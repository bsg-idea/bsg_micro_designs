

module top
(
  clk_i,
  reset_i,
  cache_pkt_i,
  v_i,
  ready_o,
  data_o,
  v_o,
  yumi_i,
  dma_pkt_o,
  dma_pkt_v_o,
  dma_pkt_yumi_i,
  dma_data_i,
  dma_data_v_i,
  dma_data_ready_o,
  dma_data_o,
  dma_data_v_o,
  dma_data_yumi_i,
  v_we_o
);

  input [68:0] cache_pkt_i;
  output [31:0] data_o;
  output [28:0] dma_pkt_o;
  input [31:0] dma_data_i;
  output [31:0] dma_data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  input dma_pkt_yumi_i;
  input dma_data_v_i;
  input dma_data_yumi_i;
  output ready_o;
  output v_o;
  output dma_pkt_v_o;
  output dma_data_ready_o;
  output dma_data_v_o;
  output v_we_o;

  bsg_cache
  wrapper
  (
    .cache_pkt_i(cache_pkt_i),
    .data_o(data_o),
    .dma_pkt_o(dma_pkt_o),
    .dma_data_i(dma_data_i),
    .dma_data_o(dma_data_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .yumi_i(yumi_i),
    .dma_pkt_yumi_i(dma_pkt_yumi_i),
    .dma_data_v_i(dma_data_v_i),
    .dma_data_yumi_i(dma_data_yumi_i),
    .ready_o(ready_o),
    .v_o(v_o),
    .dma_pkt_v_o(dma_pkt_v_o),
    .dma_data_ready_o(dma_data_ready_o),
    .dma_data_v_o(dma_data_v_o),
    .v_we_o(v_we_o)
  );


endmodule



module bsg_cache_pkt_decode_data_width_p32_addr_width_p28
(
  cache_pkt_i,
  decode_o
);

  input [68:0] cache_pkt_i;
  output [15:0] decode_o;
  wire [15:0] decode_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N42,
  N43,N44,N46,N48,N49,N50,N51,N52,N54,N56,N57,N59,N61,N62,N63,N64,N66,N67,N68,N69,
  N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,
  N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,
  N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,
  N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135;
  assign N7 = cache_pkt_i[67] | cache_pkt_i[66];
  assign N8 = N42 | N36;
  assign N9 = N7 | N8;
  assign N10 = N48 | cache_pkt_i[66];
  assign N11 = N10 | N8;
  assign N12 = cache_pkt_i[67] | N61;
  assign N13 = N12 | N8;
  assign N15 = N42 | cache_pkt_i[64];
  assign N16 = N7 | N15;
  assign N17 = N10 | N15;
  assign N18 = N12 | N15;
  assign N20 = cache_pkt_i[65] | N36;
  assign N21 = N7 | N20;
  assign N22 = N10 | N20;
  assign N23 = N12 | N20;
  assign N25 = N48 & N61;
  assign N26 = N42 & N36;
  assign N27 = N25 & N26;
  assign N28 = cache_pkt_i[65] | cache_pkt_i[64];
  assign N29 = N10 | N28;
  assign N30 = N12 | N28;
  assign N32 = cache_pkt_i[67] & cache_pkt_i[66];
  assign N35 = ~cache_pkt_i[68];
  assign N36 = ~cache_pkt_i[64];
  assign N37 = cache_pkt_i[67] | N35;
  assign N38 = cache_pkt_i[66] | N37;
  assign N39 = cache_pkt_i[65] | N38;
  assign N40 = N36 | N39;
  assign decode_o[8] = ~N40;
  assign N42 = ~cache_pkt_i[65];
  assign N43 = N42 | N38;
  assign N44 = cache_pkt_i[64] | N43;
  assign decode_o[7] = ~N44;
  assign N46 = N36 | N43;
  assign decode_o[6] = ~N46;
  assign N48 = ~cache_pkt_i[67];
  assign N49 = N48 | N35;
  assign N50 = cache_pkt_i[66] | N49;
  assign N51 = cache_pkt_i[65] | N50;
  assign N52 = cache_pkt_i[64] | N51;
  assign decode_o[5] = ~N52;
  assign N54 = N36 | N51;
  assign decode_o[4] = ~N54;
  assign N56 = N42 | N50;
  assign N57 = cache_pkt_i[64] | N56;
  assign decode_o[3] = ~N57;
  assign N59 = N36 | N56;
  assign decode_o[2] = ~N59;
  assign N61 = ~cache_pkt_i[66];
  assign N62 = N61 | N49;
  assign N63 = cache_pkt_i[65] | N62;
  assign N64 = cache_pkt_i[64] | N63;
  assign decode_o[1] = ~N64;
  assign N66 = cache_pkt_i[67] | cache_pkt_i[68];
  assign N67 = cache_pkt_i[66] | N66;
  assign N68 = cache_pkt_i[65] | N67;
  assign N69 = cache_pkt_i[64] | N68;
  assign N70 = ~N69;
  assign N71 = N36 | N68;
  assign N72 = ~N71;
  assign N73 = N42 | N67;
  assign N74 = cache_pkt_i[64] | N73;
  assign N75 = ~N74;
  assign N76 = N36 | N73;
  assign N77 = ~N76;
  assign N78 = N48 | cache_pkt_i[68];
  assign N79 = N61 | N78;
  assign N80 = cache_pkt_i[65] | N79;
  assign N81 = cache_pkt_i[64] | N80;
  assign N82 = ~N81;
  assign N83 = N36 | N80;
  assign N84 = ~N83;
  assign N85 = N61 | N66;
  assign N86 = cache_pkt_i[65] | N85;
  assign N87 = cache_pkt_i[64] | N86;
  assign N88 = ~N87;
  assign N89 = N36 | N86;
  assign N90 = ~N89;
  assign N91 = N42 | N85;
  assign N92 = cache_pkt_i[64] | N91;
  assign N93 = ~N92;
  assign N94 = N36 | N91;
  assign N95 = ~N94;
  assign N96 = cache_pkt_i[66] | N78;
  assign N97 = cache_pkt_i[65] | N96;
  assign N98 = cache_pkt_i[64] | N97;
  assign N99 = ~N98;
  assign N100 = N36 | N97;
  assign N101 = ~N100;
  assign N102 = N42 | N96;
  assign N103 = cache_pkt_i[64] | N102;
  assign N104 = ~N103;
  assign N105 = N36 | N102;
  assign N106 = ~N105;
  assign N107 = cache_pkt_i[64] | N39;
  assign decode_o[9] = ~N107;
  assign { N34, N33 } = (N0)? { 1'b1, 1'b1 } : 
                        (N1)? { 1'b1, 1'b0 } : 
                        (N2)? { 1'b0, 1'b1 } : 
                        (N3)? { 1'b0, 1'b0 } : 
                        (N4)? { 1'b0, 1'b0 } : 1'b0;
  assign N0 = N14;
  assign N1 = N19;
  assign N2 = N24;
  assign N3 = N31;
  assign N4 = N32;
  assign decode_o[15:14] = (N5)? { N34, N33 } : 
                           (N6)? { 1'b0, 1'b0 } : 1'b0;
  assign N5 = N35;
  assign N6 = cache_pkt_i[68];
  assign N14 = N111 | N112;
  assign N111 = N109 | N110;
  assign N109 = ~N9;
  assign N110 = ~N11;
  assign N112 = ~N13;
  assign N19 = N115 | N116;
  assign N115 = N113 | N114;
  assign N113 = ~N16;
  assign N114 = ~N17;
  assign N116 = ~N18;
  assign N24 = N119 | N120;
  assign N119 = N117 | N118;
  assign N117 = ~N21;
  assign N118 = ~N22;
  assign N120 = ~N23;
  assign N31 = N122 | N123;
  assign N122 = N27 | N121;
  assign N121 = ~N29;
  assign N123 = ~N30;
  assign decode_o[12] = N82 | N84;
  assign decode_o[13] = N125 | N77;
  assign N125 = N124 | N75;
  assign N124 = N70 | N72;
  assign decode_o[11] = N132 | N82;
  assign N132 = N131 | N95;
  assign N131 = N130 | N93;
  assign N130 = N129 | N90;
  assign N129 = N128 | N88;
  assign N128 = N127 | N77;
  assign N127 = N126 | N75;
  assign N126 = N70 | N72;
  assign decode_o[10] = N135 | N84;
  assign N135 = N134 | N106;
  assign N134 = N133 | N104;
  assign N133 = N99 | N101;
  assign decode_o[0] = ~decode_o[9];

endmodule



module bsg_dff_width_p1
(
  clk_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  reg [0:0] data_o;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { data_o[0:0] } <= { data_i[0:0] };
    end 
  end


endmodule



module bsg_dff_en_width_p80_harden_p0_strength_p0
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [79:0] data_i;
  output [79:0] data_o;
  input clk_i;
  input en_i;
  reg [79:0] data_o;

  always @(posedge clk_i) begin
    if(en_i) begin
      { data_o[79:0] } <= { data_i[79:0] };
    end 
  end


endmodule



module bsg_dff_en_bypass_width_p80
(
  clk_i,
  en_i,
  data_i,
  data_o
);

  input [79:0] data_i;
  output [79:0] data_o;
  input clk_i;
  input en_i;
  wire [79:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_en_width_p80_harden_p0_strength_p0
  dff
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .en_i(en_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_mem_1rw_sync_mask_write_bit_synth_width_p80_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [79:0] data_i;
  input [5:0] addr_i;
  input [79:0] w_mask_i;
  output [79:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [79:0] data_o,data_out;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,read_en,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
  llr_read_en_r,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,
  N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,
  N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,
  N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,
  N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,
  N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,
  N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,
  N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,
  N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,
  N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,
  N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,
  N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,
  N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,
  N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,
  N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,
  N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,
  N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,
  N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,
  N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,
  N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,
  N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,
  N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,
  N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,
  N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,
  N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,
  N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,
  N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,
  N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,
  N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,
  N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,
  N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,
  N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,
  N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
  N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,
  N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,
  N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,
  N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,
  N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,
  N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,
  N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,
  N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,
  N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,
  N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,
  N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,
  N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,
  N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,
  N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,
  N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,
  N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,
  N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,
  N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,
  N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,
  N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,
  N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,
  N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,
  N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,
  N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,
  N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,
  N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,
  N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,
  N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,
  N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,
  N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,
  N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,
  N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,
  N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,
  N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,
  N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,
  N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,
  N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,
  N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,
  N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,
  N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,
  N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,
  N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,
  N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,
  N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,
  N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,
  N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,
  N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,
  N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,
  N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,
  N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,
  N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,
  N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,
  N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,
  N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,
  N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,
  N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,
  N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,
  N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,
  N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,
  N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,
  N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,
  N1608,N1609,N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,
  N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,
  N1634,N1635,N1636,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,
  N1648,N1649,N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,
  N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,
  N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,
  N1688,N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,
  N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,
  N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,
  N1728,N1729,N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,
  N1741,N1742,N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,
  N1754,N1755,N1756,N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,
  N1768,N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,
  N1781,N1782,N1783,N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,
  N1794,N1795,N1796,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,
  N1808,N1809,N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,
  N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,
  N1834,N1835,N1836,N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,
  N1848,N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,
  N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,
  N1874,N1875,N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,
  N1888,N1889,N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,
  N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,
  N1914,N1915,N1916,N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,
  N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,
  N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,
  N1954,N1955,N1956,N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,
  N1968,N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,
  N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,
  N1994,N1995,N1996,N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,
  N2008,N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,
  N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,
  N2034,N2035,N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,
  N2048,N2049,N2050,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,
  N2061,N2062,N2063,N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,
  N2074,N2075,N2076,N2077,N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,
  N2088,N2089,N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,
  N2101,N2102,N2103,N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,
  N2114,N2115,N2116,N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,
  N2128,N2129,N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,
  N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,
  N2154,N2155,N2156,N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,
  N2168,N2169,N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,
  N2181,N2182,N2183,N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,
  N2194,N2195,N2196,N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,
  N2208,N2209,N2210,N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,
  N2221,N2222,N2223,N2224,N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,
  N2234,N2235,N2236,N2237,N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,
  N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,
  N2261,N2262,N2263,N2264,N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,
  N2274,N2275,N2276,N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,
  N2288,N2289,N2290,N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300,
  N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,
  N2314,N2315,N2316,N2317,N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,
  N2328,N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,
  N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,
  N2354,N2355,N2356,N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,
  N2368,N2369,N2370,N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,N2380,
  N2381,N2382,N2383,N2384,N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,
  N2394,N2395,N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2407,
  N2408,N2409,N2410,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,N2420,
  N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,
  N2434,N2435,N2436,N2437,N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,N2447,
  N2448,N2449,N2450,N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,N2460,
  N2461,N2462,N2463,N2464,N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,
  N2474,N2475,N2476,N2477,N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487,
  N2488,N2489,N2490,N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,N2500,
  N2501,N2502,N2503,N2504,N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,N2513,
  N2514,N2515,N2516,N2517,N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,N2527,
  N2528,N2529,N2530,N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,N2539,N2540,
  N2541,N2542,N2543,N2544,N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,
  N2554,N2555,N2556,N2557,N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,N2567,
  N2568,N2569,N2570,N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,N2579,N2580,
  N2581,N2582,N2583,N2584,N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,N2593,
  N2594,N2595,N2596,N2597,N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,N2607,
  N2608,N2609,N2610,N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,N2620,
  N2621,N2622,N2623,N2624,N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,N2633,
  N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,
  N2648,N2649,N2650,N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,N2659,N2660,
  N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,
  N2674,N2675,N2676,N2677,N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,N2687,
  N2688,N2689,N2690,N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,N2699,N2700,
  N2701,N2702,N2703,N2704,N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,N2713,
  N2714,N2715,N2716,N2717,N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,N2727,
  N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,N2740,
  N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,N2753,
  N2754,N2755,N2756,N2757,N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,N2767,
  N2768,N2769,N2770,N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,N2779,N2780,
  N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,N2793,
  N2794,N2795,N2796,N2797,N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806,N2807,
  N2808,N2809,N2810,N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,N2819,N2820,
  N2821,N2822,N2823,N2824,N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,
  N2834,N2835,N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,N2847,
  N2848,N2849,N2850,N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,N2859,N2860,
  N2861,N2862,N2863,N2864,N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,N2873,
  N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,N2886,N2887,
  N2888,N2889,N2890,N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,N2899,N2900,
  N2901,N2902,N2903,N2904,N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912,N2913,
  N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,
  N2928,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,N2939,N2940,
  N2941,N2942,N2943,N2944,N2945,N2946,N2947,N2948,N2949,N2950,N2951,N2952,N2953,
  N2954,N2955,N2956,N2957,N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2965,N2966,N2967,
  N2968,N2969,N2970,N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,N2979,N2980,
  N2981,N2982,N2983,N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,N2993,
  N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,N3007,
  N3008,N3009,N3010,N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,
  N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,N3033,
  N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,N3042,N3043,N3044,N3045,N3046,N3047,
  N3048,N3049,N3050,N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,
  N3061,N3062,N3063,N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,
  N3074,N3075,N3076,N3077,N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085,N3086,N3087,
  N3088,N3089,N3090,N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100,
  N3101,N3102,N3103,N3104,N3105,N3106,N3107,N3108,N3109,N3110,N3111,N3112,N3113,
  N3114,N3115,N3116,N3117,N3118,N3119,N3120,N3121,N3122,N3123,N3124,N3125,N3126,N3127,
  N3128,N3129,N3130,N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,N3139,N3140,
  N3141,N3142,N3143,N3144,N3145,N3146,N3147,N3148,N3149,N3150,N3151,N3152,N3153,
  N3154,N3155,N3156,N3157,N3158,N3159,N3160,N3161,N3162,N3163,N3164,N3165,N3166,N3167,
  N3168,N3169,N3170,N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,N3179,N3180,
  N3181,N3182,N3183,N3184,N3185,N3186,N3187,N3188,N3189,N3190,N3191,N3192,N3193,
  N3194,N3195,N3196,N3197,N3198,N3199,N3200,N3201,N3202,N3203,N3204,N3205,N3206,N3207,
  N3208,N3209,N3210,N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,N3219,N3220,
  N3221,N3222,N3223,N3224,N3225,N3226,N3227,N3228,N3229,N3230,N3231,N3232,N3233,
  N3234,N3235,N3236,N3237,N3238,N3239,N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247,
  N3248,N3249,N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,N3260,
  N3261,N3262,N3263,N3264,N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272,N3273,
  N3274,N3275,N3276,N3277,N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,
  N3288,N3289,N3290,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299,N3300,
  N3301,N3302,N3303,N3304,N3305,N3306,N3307,N3308,N3309,N3310,N3311,N3312,N3313,
  N3314,N3315,N3316,N3317,N3318,N3319,N3320,N3321,N3322,N3323,N3324,N3325,N3326,N3327,
  N3328,N3329,N3330,N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,N3339,N3340,
  N3341,N3342,N3343,N3344,N3345,N3346,N3347,N3348,N3349,N3350,N3351,N3352,N3353,
  N3354,N3355,N3356,N3357,N3358,N3359,N3360,N3361,N3362,N3363,N3364,N3365,N3366,N3367,
  N3368,N3369,N3370,N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,N3379,N3380,
  N3381,N3382,N3383,N3384,N3385,N3386,N3387,N3388,N3389,N3390,N3391,N3392,N3393,
  N3394,N3395,N3396,N3397,N3398,N3399,N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,
  N3408,N3409,N3410,N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,N3419,N3420,
  N3421,N3422,N3423,N3424,N3425,N3426,N3427,N3428,N3429,N3430,N3431,N3432,N3433,
  N3434,N3435,N3436,N3437,N3438,N3439,N3440,N3441,N3442,N3443,N3444,N3445,N3446,N3447,
  N3448,N3449,N3450,N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,N3459,N3460,
  N3461,N3462,N3463,N3464,N3465,N3466,N3467,N3468,N3469,N3470,N3471,N3472,N3473,
  N3474,N3475,N3476,N3477,N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,N3487,
  N3488,N3489,N3490,N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,N3499,N3500,
  N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,N3513,
  N3514,N3515,N3516,N3517,N3518,N3519,N3520,N3521,N3522,N3523,N3524,N3525,N3526,N3527,
  N3528,N3529,N3530,N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538,N3539,N3540,
  N3541,N3542,N3543,N3544,N3545,N3546,N3547,N3548,N3549,N3550,N3551,N3552,N3553,
  N3554,N3555,N3556,N3557,N3558,N3559,N3560,N3561,N3562,N3563,N3564,N3565,N3566,N3567,
  N3568,N3569,N3570,N3571,N3572,N3573,N3574,N3575,N3576,N3577,N3578,N3579,N3580,
  N3581,N3582,N3583,N3584,N3585,N3586,N3587,N3588,N3589,N3590,N3591,N3592,N3593,
  N3594,N3595,N3596,N3597,N3598,N3599,N3600,N3601,N3602,N3603,N3604,N3605,N3606,N3607,
  N3608,N3609,N3610,N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618,N3619,N3620,
  N3621,N3622,N3623,N3624,N3625,N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,
  N3634,N3635,N3636,N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3646,N3647,
  N3648,N3649,N3650,N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,N3659,N3660,
  N3661,N3662,N3663,N3664,N3665,N3666,N3667,N3668,N3669,N3670,N3671,N3672,N3673,
  N3674,N3675,N3676,N3677,N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685,N3686,N3687,
  N3688,N3689,N3690,N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3698,N3699,N3700,
  N3701,N3702,N3703,N3704,N3705,N3706,N3707,N3708,N3709,N3710,N3711,N3712,N3713,
  N3714,N3715,N3716,N3717,N3718,N3719,N3720,N3721,N3722,N3723,N3724,N3725,N3726,N3727,
  N3728,N3729,N3730,N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3738,N3739,N3740,
  N3741,N3742,N3743,N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3751,N3752,N3753,
  N3754,N3755,N3756,N3757,N3758,N3759,N3760,N3761,N3762,N3763,N3764,N3765,N3766,N3767,
  N3768,N3769,N3770,N3771,N3772,N3773,N3774,N3775,N3776,N3777,N3778,N3779,N3780,
  N3781,N3782,N3783,N3784,N3785,N3786,N3787,N3788,N3789,N3790,N3791,N3792,N3793,
  N3794,N3795,N3796,N3797,N3798,N3799,N3800,N3801,N3802,N3803,N3804,N3805,N3806,N3807,
  N3808,N3809,N3810,N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,N3819,N3820,
  N3821,N3822,N3823,N3824,N3825,N3826,N3827,N3828,N3829,N3830,N3831,N3832,N3833,
  N3834,N3835,N3836,N3837,N3838,N3839,N3840,N3841,N3842,N3843,N3844,N3845,N3846,N3847,
  N3848,N3849,N3850,N3851,N3852,N3853,N3854,N3855,N3856,N3857,N3858,N3859,N3860,
  N3861,N3862,N3863,N3864,N3865,N3866,N3867,N3868,N3869,N3870,N3871,N3872,N3873,
  N3874,N3875,N3876,N3877,N3878,N3879,N3880,N3881,N3882,N3883,N3884,N3885,N3886,N3887,
  N3888,N3889,N3890,N3891,N3892,N3893,N3894,N3895,N3896,N3897,N3898,N3899,N3900,
  N3901,N3902,N3903,N3904,N3905,N3906,N3907,N3908,N3909,N3910,N3911,N3912,N3913,
  N3914,N3915,N3916,N3917,N3918,N3919,N3920,N3921,N3922,N3923,N3924,N3925,N3926,N3927,
  N3928,N3929,N3930,N3931,N3932,N3933,N3934,N3935,N3936,N3937,N3938,N3939,N3940,
  N3941,N3942,N3943,N3944,N3945,N3946,N3947,N3948,N3949,N3950,N3951,N3952,N3953,
  N3954,N3955,N3956,N3957,N3958,N3959,N3960,N3961,N3962,N3963,N3964,N3965,N3966,N3967,
  N3968,N3969,N3970,N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3978,N3979,N3980,
  N3981,N3982,N3983,N3984,N3985,N3986,N3987,N3988,N3989,N3990,N3991,N3992,N3993,
  N3994,N3995,N3996,N3997,N3998,N3999,N4000,N4001,N4002,N4003,N4004,N4005,N4006,N4007,
  N4008,N4009,N4010,N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,N4019,N4020,
  N4021,N4022,N4023,N4024,N4025,N4026,N4027,N4028,N4029,N4030,N4031,N4032,N4033,
  N4034,N4035,N4036,N4037,N4038,N4039,N4040,N4041,N4042,N4043,N4044,N4045,N4046,N4047,
  N4048,N4049,N4050,N4051,N4052,N4053,N4054,N4055,N4056,N4057,N4058,N4059,N4060,
  N4061,N4062,N4063,N4064,N4065,N4066,N4067,N4068,N4069,N4070,N4071,N4072,N4073,
  N4074,N4075,N4076,N4077,N4078,N4079,N4080,N4081,N4082,N4083,N4084,N4085,N4086,N4087,
  N4088,N4089,N4090,N4091,N4092,N4093,N4094,N4095,N4096,N4097,N4098,N4099,N4100,
  N4101,N4102,N4103,N4104,N4105,N4106,N4107,N4108,N4109,N4110,N4111,N4112,N4113,
  N4114,N4115,N4116,N4117,N4118,N4119,N4120,N4121,N4122,N4123,N4124,N4125,N4126,N4127,
  N4128,N4129,N4130,N4131,N4132,N4133,N4134,N4135,N4136,N4137,N4138,N4139,N4140,
  N4141,N4142,N4143,N4144,N4145,N4146,N4147,N4148,N4149,N4150,N4151,N4152,N4153,
  N4154,N4155,N4156,N4157,N4158,N4159,N4160,N4161,N4162,N4163,N4164,N4165,N4166,N4167,
  N4168,N4169,N4170,N4171,N4172,N4173,N4174,N4175,N4176,N4177,N4178,N4179,N4180,
  N4181,N4182,N4183,N4184,N4185,N4186,N4187,N4188,N4189,N4190,N4191,N4192,N4193,
  N4194,N4195,N4196,N4197,N4198,N4199,N4200,N4201,N4202,N4203,N4204,N4205,N4206,N4207,
  N4208,N4209,N4210,N4211,N4212,N4213,N4214,N4215,N4216,N4217,N4218,N4219,N4220,
  N4221,N4222,N4223,N4224,N4225,N4226,N4227,N4228,N4229,N4230,N4231,N4232,N4233,
  N4234,N4235,N4236,N4237,N4238,N4239,N4240,N4241,N4242,N4243,N4244,N4245,N4246,N4247,
  N4248,N4249,N4250,N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,N4259,N4260,
  N4261,N4262,N4263,N4264,N4265,N4266,N4267,N4268,N4269,N4270,N4271,N4272,N4273,
  N4274,N4275,N4276,N4277,N4278,N4279,N4280,N4281,N4282,N4283,N4284,N4285,N4286,N4287,
  N4288,N4289,N4290,N4291,N4292,N4293,N4294,N4295,N4296,N4297,N4298,N4299,N4300,
  N4301,N4302,N4303,N4304,N4305,N4306,N4307,N4308,N4309,N4310,N4311,N4312,N4313,
  N4314,N4315,N4316,N4317,N4318,N4319,N4320,N4321,N4322,N4323,N4324,N4325,N4326,N4327,
  N4328,N4329,N4330,N4331,N4332,N4333,N4334,N4335,N4336,N4337,N4338,N4339,N4340,
  N4341,N4342,N4343,N4344,N4345,N4346,N4347,N4348,N4349,N4350,N4351,N4352,N4353,
  N4354,N4355,N4356,N4357,N4358,N4359,N4360,N4361,N4362,N4363,N4364,N4365,N4366,N4367,
  N4368,N4369,N4370,N4371,N4372,N4373,N4374,N4375,N4376,N4377,N4378,N4379,N4380,
  N4381,N4382,N4383,N4384,N4385,N4386,N4387,N4388,N4389,N4390,N4391,N4392,N4393,
  N4394,N4395,N4396,N4397,N4398,N4399,N4400,N4401,N4402,N4403,N4404,N4405,N4406,N4407,
  N4408,N4409,N4410,N4411,N4412,N4413,N4414,N4415,N4416,N4417,N4418,N4419,N4420,
  N4421,N4422,N4423,N4424,N4425,N4426,N4427,N4428,N4429,N4430,N4431,N4432,N4433,
  N4434,N4435,N4436,N4437,N4438,N4439,N4440,N4441,N4442,N4443,N4444,N4445,N4446,N4447,
  N4448,N4449,N4450,N4451,N4452,N4453,N4454,N4455,N4456,N4457,N4458,N4459,N4460,
  N4461,N4462,N4463,N4464,N4465,N4466,N4467,N4468,N4469,N4470,N4471,N4472,N4473,
  N4474,N4475,N4476,N4477,N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,N4486,N4487,
  N4488,N4489,N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498,N4499,N4500,
  N4501,N4502,N4503,N4504,N4505,N4506,N4507,N4508,N4509,N4510,N4511,N4512,N4513,
  N4514,N4515,N4516,N4517,N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,N4527,
  N4528,N4529,N4530,N4531,N4532,N4533,N4534,N4535,N4536,N4537,N4538,N4539,N4540,
  N4541,N4542,N4543,N4544,N4545,N4546,N4547,N4548,N4549,N4550,N4551,N4552,N4553,
  N4554,N4555,N4556,N4557,N4558,N4559,N4560,N4561,N4562,N4563,N4564,N4565,N4566,N4567,
  N4568,N4569,N4570,N4571,N4572,N4573,N4574,N4575,N4576,N4577,N4578,N4579,N4580,
  N4581,N4582,N4583,N4584,N4585,N4586,N4587,N4588,N4589,N4590,N4591,N4592,N4593,
  N4594,N4595,N4596,N4597,N4598,N4599,N4600,N4601,N4602,N4603,N4604,N4605,N4606,N4607,
  N4608,N4609,N4610,N4611,N4612,N4613,N4614,N4615,N4616,N4617,N4618,N4619,N4620,
  N4621,N4622,N4623,N4624,N4625,N4626,N4627,N4628,N4629,N4630,N4631,N4632,N4633,
  N4634,N4635,N4636,N4637,N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,N4647,
  N4648,N4649,N4650,N4651,N4652,N4653,N4654,N4655,N4656,N4657,N4658,N4659,N4660,
  N4661,N4662,N4663,N4664,N4665,N4666,N4667,N4668,N4669,N4670,N4671,N4672,N4673,
  N4674,N4675,N4676,N4677,N4678,N4679,N4680,N4681,N4682,N4683,N4684,N4685,N4686,N4687,
  N4688,N4689,N4690,N4691,N4692,N4693,N4694,N4695,N4696,N4697,N4698,N4699,N4700,
  N4701,N4702,N4703,N4704,N4705,N4706,N4707,N4708,N4709,N4710,N4711,N4712,N4713,
  N4714,N4715,N4716,N4717,N4718,N4719,N4720,N4721,N4722,N4723,N4724,N4725,N4726,N4727,
  N4728,N4729,N4730,N4731,N4732,N4733,N4734,N4735,N4736,N4737,N4738,N4739,N4740,
  N4741,N4742,N4743,N4744,N4745,N4746,N4747,N4748,N4749,N4750,N4751,N4752,N4753,
  N4754,N4755,N4756,N4757,N4758,N4759,N4760,N4761,N4762,N4763,N4764,N4765,N4766,N4767,
  N4768,N4769,N4770,N4771,N4772,N4773,N4774,N4775,N4776,N4777,N4778,N4779,N4780,
  N4781,N4782,N4783,N4784,N4785,N4786,N4787,N4788,N4789,N4790,N4791,N4792,N4793,
  N4794,N4795,N4796,N4797,N4798,N4799,N4800,N4801,N4802,N4803,N4804,N4805,N4806,N4807,
  N4808,N4809,N4810,N4811,N4812,N4813,N4814,N4815,N4816,N4817,N4818,N4819,N4820,
  N4821,N4822,N4823,N4824,N4825,N4826,N4827,N4828,N4829,N4830,N4831,N4832,N4833,
  N4834,N4835,N4836,N4837,N4838,N4839,N4840,N4841,N4842,N4843,N4844,N4845,N4846,N4847,
  N4848,N4849,N4850,N4851,N4852,N4853,N4854,N4855,N4856,N4857,N4858,N4859,N4860,
  N4861,N4862,N4863,N4864,N4865,N4866,N4867,N4868,N4869,N4870,N4871,N4872,N4873,
  N4874,N4875,N4876,N4877,N4878,N4879,N4880,N4881,N4882,N4883,N4884,N4885,N4886,N4887,
  N4888,N4889,N4890,N4891,N4892,N4893,N4894,N4895,N4896,N4897,N4898,N4899,N4900,
  N4901,N4902,N4903,N4904,N4905,N4906,N4907,N4908,N4909,N4910,N4911,N4912,N4913,
  N4914,N4915,N4916,N4917,N4918,N4919,N4920,N4921,N4922,N4923,N4924,N4925,N4926,N4927,
  N4928,N4929,N4930,N4931,N4932,N4933,N4934,N4935,N4936,N4937,N4938,N4939,N4940,
  N4941,N4942,N4943,N4944,N4945,N4946,N4947,N4948,N4949,N4950,N4951,N4952,N4953,
  N4954,N4955,N4956,N4957,N4958,N4959,N4960,N4961,N4962,N4963,N4964,N4965,N4966,N4967,
  N4968,N4969,N4970,N4971,N4972,N4973,N4974,N4975,N4976,N4977,N4978,N4979,N4980,
  N4981,N4982,N4983,N4984,N4985,N4986,N4987,N4988,N4989,N4990,N4991,N4992,N4993,
  N4994,N4995,N4996,N4997,N4998,N4999,N5000,N5001,N5002,N5003,N5004,N5005,N5006,N5007,
  N5008,N5009,N5010,N5011,N5012,N5013,N5014,N5015,N5016,N5017,N5018,N5019,N5020,
  N5021,N5022,N5023,N5024,N5025,N5026,N5027,N5028,N5029,N5030,N5031,N5032,N5033,
  N5034,N5035,N5036,N5037,N5038,N5039,N5040,N5041,N5042,N5043,N5044,N5045,N5046,N5047,
  N5048,N5049,N5050,N5051,N5052,N5053,N5054,N5055,N5056,N5057,N5058,N5059,N5060,
  N5061,N5062,N5063,N5064,N5065,N5066,N5067,N5068,N5069,N5070,N5071,N5072,N5073,
  N5074,N5075,N5076,N5077,N5078,N5079,N5080,N5081,N5082,N5083,N5084,N5085,N5086,N5087,
  N5088,N5089,N5090,N5091,N5092,N5093,N5094,N5095,N5096,N5097,N5098,N5099,N5100,
  N5101,N5102,N5103,N5104,N5105,N5106,N5107,N5108,N5109,N5110,N5111,N5112,N5113,
  N5114,N5115,N5116,N5117,N5118,N5119,N5120,N5121,N5122,N5123,N5124,N5125,N5126,N5127,
  N5128,N5129,N5130,N5131,N5132,N5133,N5134,N5135,N5136,N5137,N5138,N5139,N5140,
  N5141,N5142,N5143,N5144,N5145,N5146,N5147,N5148,N5149,N5150,N5151,N5152,N5153,
  N5154,N5155,N5156,N5157,N5158,N5159,N5160,N5161,N5162,N5163,N5164,N5165,N5166,N5167,
  N5168,N5169,N5170,N5171,N5172,N5173,N5174,N5175,N5176,N5177,N5178,N5179,N5180,
  N5181,N5182,N5183,N5184,N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,N5193,
  N5194,N5195,N5196,N5197,N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,N5207,
  N5208,N5209,N5210,N5211,N5212,N5213,N5214,N5215,N5216,N5217,N5218,N5219,N5220,
  N5221,N5222,N5223,N5224,N5225,N5226,N5227,N5228,N5229,N5230,N5231,N5232,N5233,
  N5234,N5235,N5236,N5237,N5238,N5239,N5240,N5241,N5242,N5243,N5244,N5245,N5246,N5247,
  N5248,N5249,N5250,N5251,N5252,N5253,N5254,N5255,N5256,N5257,N5258,N5259,N5260,
  N5261,N5262,N5263,N5264,N5265,N5266,N5267,N5268,N5269,N5270,N5271,N5272,N5273,
  N5274,N5275,N5276,N5277,N5278,N5279,N5280,N5281,N5282,N5283,N5284,N5285,N5286,N5287,
  N5288,N5289,N5290,N5291,N5292,N5293,N5294,N5295,N5296,N5297,N5298,N5299,N5300,
  N5301,N5302,N5303,N5304,N5305,N5306,N5307,N5308,N5309,N5310,N5311,N5312,N5313,
  N5314,N5315,N5316,N5317,N5318,N5319,N5320,N5321,N5322,N5323,N5324,N5325,N5326,N5327,
  N5328,N5329,N5330,N5331,N5332,N5333,N5334,N5335,N5336,N5337,N5338,N5339,N5340,
  N5341,N5342,N5343,N5344,N5345,N5346,N5347,N5348,N5349,N5350,N5351,N5352,N5353,
  N5354,N5355,N5356,N5357,N5358,N5359,N5360,N5361,N5362,N5363,N5364,N5365,N5366,N5367,
  N5368,N5369,N5370,N5371,N5372,N5373,N5374,N5375,N5376,N5377,N5378,N5379,N5380,
  N5381,N5382,N5383,N5384,N5385,N5386,N5387,N5388,N5389,N5390,N5391,N5392,N5393,
  N5394,N5395,N5396,N5397,N5398,N5399,N5400,N5401,N5402,N5403,N5404,N5405,N5406,N5407,
  N5408,N5409,N5410,N5411,N5412,N5413,N5414,N5415,N5416,N5417,N5418,N5419,N5420,
  N5421,N5422,N5423,N5424,N5425,N5426,N5427,N5428,N5429,N5430,N5431,N5432,N5433,
  N5434,N5435,N5436,N5437,N5438,N5439,N5440,N5441,N5442,N5443,N5444,N5445,N5446,N5447,
  N5448,N5449,N5450,N5451,N5452,N5453,N5454,N5455,N5456,N5457,N5458,N5459,N5460,
  N5461,N5462,N5463,N5464,N5465,N5466,N5467,N5468,N5469,N5470,N5471,N5472,N5473,
  N5474,N5475,N5476,N5477,N5478,N5479,N5480,N5481,N5482,N5483,N5484,N5485,N5486,N5487,
  N5488,N5489,N5490,N5491,N5492,N5493,N5494,N5495,N5496,N5497,N5498,N5499,N5500,
  N5501,N5502,N5503,N5504,N5505,N5506,N5507,N5508,N5509,N5510,N5511,N5512,N5513,
  N5514,N5515,N5516,N5517,N5518,N5519,N5520,N5521,N5522,N5523,N5524,N5525,N5526,N5527,
  N5528,N5529,N5530,N5531,N5532,N5533,N5534,N5535,N5536,N5537,N5538,N5539,N5540,
  N5541,N5542,N5543,N5544,N5545,N5546,N5547,N5548,N5549,N5550,N5551,N5552,N5553,
  N5554,N5555,N5556,N5557,N5558,N5559,N5560,N5561,N5562,N5563,N5564,N5565,N5566,N5567,
  N5568,N5569,N5570,N5571,N5572,N5573,N5574,N5575,N5576,N5577,N5578,N5579,N5580,
  N5581,N5582,N5583,N5584,N5585,N5586,N5587,N5588,N5589,N5590,N5591,N5592,N5593,
  N5594,N5595,N5596,N5597,N5598,N5599,N5600,N5601,N5602,N5603,N5604,N5605,N5606,N5607,
  N5608,N5609,N5610,N5611,N5612,N5613,N5614,N5615,N5616,N5617,N5618,N5619,N5620,
  N5621,N5622,N5623,N5624,N5625,N5626,N5627,N5628,N5629,N5630,N5631,N5632,N5633,
  N5634,N5635,N5636,N5637,N5638,N5639,N5640,N5641,N5642,N5643,N5644,N5645,N5646,N5647,
  N5648,N5649,N5650,N5651,N5652,N5653,N5654,N5655,N5656,N5657,N5658,N5659,N5660,
  N5661,N5662,N5663,N5664,N5665,N5666,N5667,N5668,N5669,N5670,N5671,N5672,N5673,
  N5674,N5675,N5676,N5677,N5678,N5679,N5680,N5681,N5682,N5683,N5684,N5685,N5686,N5687,
  N5688,N5689,N5690,N5691,N5692,N5693,N5694,N5695,N5696,N5697,N5698,N5699,N5700,
  N5701,N5702,N5703,N5704,N5705,N5706,N5707,N5708,N5709,N5710,N5711,N5712,N5713,
  N5714,N5715,N5716,N5717,N5718,N5719,N5720,N5721,N5722,N5723,N5724,N5725,N5726,N5727,
  N5728,N5729,N5730,N5731,N5732,N5733,N5734,N5735,N5736,N5737,N5738,N5739,N5740,
  N5741,N5742,N5743,N5744,N5745,N5746,N5747,N5748,N5749,N5750,N5751,N5752,N5753,
  N5754,N5755,N5756,N5757,N5758,N5759,N5760,N5761,N5762,N5763,N5764,N5765,N5766,N5767,
  N5768,N5769,N5770,N5771,N5772,N5773,N5774,N5775,N5776,N5777,N5778,N5779,N5780,
  N5781,N5782,N5783,N5784,N5785,N5786,N5787,N5788,N5789,N5790,N5791,N5792,N5793,
  N5794,N5795,N5796,N5797,N5798,N5799,N5800,N5801,N5802,N5803,N5804,N5805,N5806,N5807,
  N5808,N5809,N5810,N5811,N5812,N5813,N5814,N5815,N5816,N5817,N5818,N5819,N5820,
  N5821,N5822,N5823,N5824,N5825,N5826,N5827,N5828,N5829,N5830,N5831,N5832,N5833,
  N5834,N5835,N5836,N5837,N5838,N5839,N5840,N5841,N5842,N5843,N5844,N5845,N5846,N5847,
  N5848,N5849,N5850,N5851,N5852,N5853,N5854,N5855,N5856,N5857,N5858,N5859,N5860,
  N5861,N5862,N5863,N5864,N5865,N5866,N5867,N5868,N5869,N5870,N5871,N5872,N5873,
  N5874,N5875,N5876,N5877,N5878,N5879,N5880,N5881,N5882,N5883,N5884,N5885,N5886,N5887,
  N5888,N5889,N5890,N5891,N5892,N5893,N5894,N5895,N5896,N5897,N5898,N5899,N5900,
  N5901,N5902,N5903,N5904,N5905,N5906,N5907,N5908,N5909,N5910,N5911,N5912,N5913,
  N5914,N5915,N5916,N5917,N5918,N5919,N5920,N5921,N5922,N5923,N5924,N5925,N5926,N5927,
  N5928,N5929,N5930,N5931,N5932,N5933,N5934,N5935,N5936,N5937,N5938,N5939,N5940,
  N5941,N5942,N5943,N5944,N5945,N5946,N5947,N5948,N5949,N5950,N5951,N5952,N5953,
  N5954,N5955,N5956,N5957,N5958,N5959,N5960,N5961,N5962,N5963,N5964,N5965,N5966,N5967,
  N5968,N5969,N5970,N5971,N5972,N5973,N5974,N5975,N5976,N5977,N5978,N5979,N5980,
  N5981,N5982,N5983,N5984,N5985,N5986,N5987,N5988,N5989,N5990,N5991,N5992,N5993,
  N5994,N5995,N5996,N5997,N5998,N5999,N6000,N6001,N6002,N6003,N6004,N6005,N6006,N6007,
  N6008,N6009,N6010,N6011,N6012,N6013,N6014,N6015,N6016,N6017,N6018,N6019,N6020,
  N6021,N6022,N6023,N6024,N6025,N6026,N6027,N6028,N6029,N6030,N6031,N6032,N6033,
  N6034,N6035,N6036,N6037,N6038,N6039,N6040,N6041,N6042,N6043,N6044,N6045,N6046,N6047,
  N6048,N6049,N6050,N6051,N6052,N6053,N6054,N6055,N6056,N6057,N6058,N6059,N6060,
  N6061,N6062,N6063,N6064,N6065,N6066,N6067,N6068,N6069,N6070,N6071,N6072,N6073,
  N6074,N6075,N6076,N6077,N6078,N6079,N6080,N6081,N6082,N6083,N6084,N6085,N6086,N6087,
  N6088,N6089,N6090,N6091,N6092,N6093,N6094,N6095,N6096,N6097,N6098,N6099,N6100,
  N6101,N6102,N6103,N6104,N6105,N6106,N6107,N6108,N6109,N6110,N6111,N6112,N6113,
  N6114,N6115,N6116,N6117,N6118,N6119,N6120,N6121,N6122,N6123,N6124,N6125,N6126,N6127,
  N6128,N6129,N6130,N6131,N6132,N6133,N6134,N6135,N6136,N6137,N6138,N6139,N6140,
  N6141,N6142,N6143,N6144,N6145,N6146,N6147,N6148,N6149,N6150,N6151,N6152,N6153,
  N6154,N6155,N6156,N6157,N6158,N6159,N6160,N6161,N6162,N6163,N6164,N6165,N6166,N6167,
  N6168,N6169,N6170,N6171,N6172,N6173,N6174,N6175,N6176,N6177,N6178,N6179,N6180,
  N6181,N6182,N6183,N6184,N6185,N6186,N6187,N6188,N6189,N6190,N6191,N6192,N6193,
  N6194,N6195,N6196,N6197,N6198,N6199,N6200,N6201,N6202,N6203,N6204,N6205,N6206,N6207,
  N6208,N6209,N6210,N6211,N6212,N6213,N6214,N6215,N6216,N6217,N6218,N6219,N6220,
  N6221,N6222,N6223,N6224,N6225,N6226,N6227,N6228,N6229,N6230,N6231,N6232,N6233,
  N6234,N6235,N6236,N6237,N6238,N6239,N6240,N6241,N6242,N6243,N6244,N6245,N6246,N6247,
  N6248,N6249,N6250,N6251,N6252,N6253,N6254,N6255,N6256,N6257,N6258,N6259,N6260,
  N6261,N6262,N6263,N6264,N6265,N6266,N6267,N6268,N6269,N6270,N6271,N6272,N6273,
  N6274,N6275,N6276,N6277,N6278,N6279,N6280,N6281,N6282,N6283,N6284,N6285,N6286,N6287,
  N6288,N6289,N6290,N6291,N6292,N6293,N6294,N6295,N6296,N6297,N6298,N6299,N6300,
  N6301,N6302,N6303,N6304,N6305,N6306,N6307,N6308,N6309,N6310,N6311,N6312,N6313,
  N6314,N6315,N6316,N6317,N6318,N6319,N6320,N6321,N6322,N6323,N6324,N6325,N6326,N6327,
  N6328,N6329,N6330,N6331,N6332,N6333,N6334,N6335,N6336,N6337,N6338,N6339,N6340,
  N6341,N6342,N6343,N6344,N6345,N6346,N6347,N6348,N6349,N6350,N6351,N6352,N6353,
  N6354,N6355,N6356,N6357,N6358,N6359,N6360,N6361,N6362,N6363,N6364,N6365,N6366,N6367,
  N6368,N6369,N6370,N6371,N6372,N6373,N6374,N6375,N6376,N6377,N6378,N6379,N6380,
  N6381,N6382,N6383,N6384,N6385,N6386,N6387,N6388,N6389,N6390,N6391,N6392,N6393,
  N6394,N6395,N6396,N6397,N6398,N6399,N6400,N6401,N6402,N6403,N6404,N6405,N6406,N6407,
  N6408,N6409,N6410,N6411,N6412,N6413,N6414,N6415,N6416,N6417,N6418,N6419,N6420,
  N6421,N6422,N6423,N6424,N6425,N6426,N6427,N6428,N6429,N6430,N6431,N6432,N6433,
  N6434,N6435,N6436,N6437,N6438,N6439,N6440,N6441,N6442,N6443,N6444,N6445,N6446,N6447,
  N6448,N6449,N6450,N6451,N6452,N6453,N6454,N6455,N6456,N6457,N6458,N6459,N6460,
  N6461,N6462,N6463,N6464,N6465,N6466,N6467,N6468,N6469,N6470,N6471,N6472,N6473,
  N6474,N6475,N6476,N6477,N6478,N6479,N6480,N6481,N6482,N6483,N6484,N6485,N6486,N6487,
  N6488,N6489,N6490,N6491,N6492,N6493,N6494,N6495,N6496,N6497,N6498,N6499,N6500,
  N6501,N6502,N6503,N6504,N6505,N6506,N6507,N6508,N6509,N6510,N6511,N6512,N6513,
  N6514,N6515,N6516,N6517,N6518,N6519,N6520,N6521,N6522,N6523,N6524,N6525,N6526,N6527,
  N6528,N6529,N6530,N6531,N6532,N6533,N6534,N6535,N6536,N6537,N6538,N6539,N6540,
  N6541,N6542,N6543,N6544,N6545,N6546,N6547,N6548,N6549,N6550,N6551,N6552,N6553,
  N6554,N6555,N6556,N6557,N6558,N6559,N6560,N6561,N6562,N6563,N6564,N6565,N6566,N6567,
  N6568,N6569,N6570,N6571,N6572,N6573,N6574,N6575,N6576,N6577,N6578,N6579,N6580,
  N6581,N6582,N6583,N6584,N6585,N6586,N6587,N6588,N6589,N6590,N6591,N6592,N6593,
  N6594,N6595,N6596,N6597,N6598,N6599,N6600,N6601,N6602,N6603,N6604,N6605,N6606,N6607,
  N6608,N6609,N6610,N6611,N6612,N6613,N6614,N6615,N6616,N6617,N6618,N6619,N6620,
  N6621,N6622,N6623,N6624,N6625,N6626,N6627,N6628,N6629,N6630,N6631,N6632,N6633,
  N6634,N6635,N6636,N6637,N6638,N6639,N6640,N6641,N6642,N6643,N6644,N6645,N6646,N6647,
  N6648,N6649,N6650,N6651,N6652,N6653,N6654,N6655,N6656,N6657,N6658,N6659,N6660,
  N6661,N6662,N6663,N6664,N6665,N6666,N6667,N6668,N6669,N6670,N6671,N6672,N6673,
  N6674,N6675,N6676,N6677,N6678,N6679,N6680,N6681,N6682,N6683,N6684,N6685,N6686,N6687,
  N6688,N6689,N6690,N6691,N6692,N6693,N6694,N6695,N6696,N6697,N6698,N6699,N6700,
  N6701,N6702,N6703,N6704,N6705,N6706,N6707,N6708,N6709,N6710,N6711,N6712,N6713,
  N6714,N6715,N6716,N6717,N6718,N6719,N6720,N6721,N6722,N6723,N6724,N6725,N6726,N6727,
  N6728,N6729,N6730,N6731,N6732,N6733,N6734,N6735,N6736,N6737,N6738,N6739,N6740,
  N6741,N6742,N6743,N6744,N6745,N6746,N6747,N6748,N6749,N6750,N6751,N6752,N6753,
  N6754,N6755,N6756,N6757,N6758,N6759,N6760,N6761,N6762,N6763,N6764,N6765,N6766,N6767,
  N6768,N6769,N6770,N6771,N6772,N6773,N6774,N6775,N6776,N6777,N6778,N6779,N6780,
  N6781,N6782,N6783,N6784,N6785,N6786,N6787,N6788,N6789,N6790,N6791,N6792,N6793,
  N6794,N6795,N6796,N6797,N6798,N6799,N6800,N6801,N6802,N6803,N6804,N6805,N6806,N6807,
  N6808,N6809,N6810,N6811,N6812,N6813,N6814,N6815,N6816,N6817,N6818,N6819,N6820,
  N6821,N6822,N6823,N6824,N6825,N6826,N6827,N6828,N6829,N6830,N6831,N6832,N6833,
  N6834,N6835,N6836,N6837,N6838,N6839,N6840,N6841,N6842,N6843,N6844,N6845,N6846,N6847,
  N6848,N6849,N6850,N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6858,N6859,N6860,
  N6861,N6862,N6863,N6864,N6865,N6866,N6867,N6868,N6869,N6870,N6871,N6872,N6873,
  N6874,N6875,N6876,N6877,N6878,N6879,N6880,N6881,N6882,N6883,N6884,N6885,N6886,N6887,
  N6888,N6889,N6890,N6891,N6892,N6893,N6894,N6895,N6896,N6897,N6898,N6899,N6900,
  N6901,N6902,N6903,N6904,N6905,N6906,N6907,N6908,N6909,N6910,N6911,N6912,N6913,
  N6914,N6915,N6916,N6917,N6918,N6919,N6920,N6921,N6922,N6923,N6924,N6925,N6926,N6927,
  N6928,N6929,N6930,N6931,N6932,N6933,N6934,N6935,N6936,N6937,N6938,N6939,N6940,
  N6941,N6942,N6943,N6944,N6945,N6946,N6947,N6948,N6949,N6950,N6951,N6952,N6953,
  N6954,N6955,N6956,N6957,N6958,N6959,N6960,N6961,N6962,N6963,N6964,N6965,N6966,N6967,
  N6968,N6969,N6970,N6971,N6972,N6973,N6974,N6975,N6976,N6977,N6978,N6979,N6980,
  N6981,N6982,N6983,N6984,N6985,N6986,N6987,N6988,N6989,N6990,N6991,N6992,N6993,
  N6994,N6995,N6996,N6997,N6998,N6999,N7000,N7001,N7002,N7003,N7004,N7005,N7006,N7007,
  N7008,N7009,N7010,N7011,N7012,N7013,N7014,N7015,N7016,N7017,N7018,N7019,N7020,
  N7021,N7022,N7023,N7024,N7025,N7026,N7027,N7028,N7029,N7030,N7031,N7032,N7033,
  N7034,N7035,N7036,N7037,N7038,N7039,N7040,N7041,N7042,N7043,N7044,N7045,N7046,N7047,
  N7048,N7049,N7050,N7051,N7052,N7053,N7054,N7055,N7056,N7057,N7058,N7059,N7060,
  N7061,N7062,N7063,N7064,N7065,N7066,N7067,N7068,N7069,N7070,N7071,N7072,N7073,
  N7074,N7075,N7076,N7077,N7078,N7079,N7080,N7081,N7082,N7083,N7084,N7085,N7086,N7087,
  N7088,N7089,N7090,N7091,N7092,N7093,N7094,N7095,N7096,N7097,N7098,N7099,N7100,
  N7101,N7102,N7103,N7104,N7105,N7106,N7107,N7108,N7109,N7110,N7111,N7112,N7113,
  N7114,N7115,N7116,N7117,N7118,N7119,N7120,N7121,N7122,N7123,N7124,N7125,N7126,N7127,
  N7128,N7129,N7130,N7131,N7132,N7133,N7134,N7135,N7136,N7137,N7138,N7139,N7140,
  N7141,N7142,N7143,N7144,N7145,N7146,N7147,N7148,N7149,N7150,N7151,N7152,N7153,
  N7154,N7155,N7156,N7157,N7158,N7159,N7160,N7161,N7162,N7163,N7164,N7165,N7166,N7167,
  N7168,N7169,N7170,N7171,N7172,N7173,N7174,N7175,N7176,N7177,N7178,N7179,N7180,
  N7181,N7182,N7183,N7184,N7185,N7186,N7187,N7188,N7189,N7190,N7191,N7192,N7193,
  N7194,N7195,N7196,N7197,N7198,N7199,N7200,N7201,N7202,N7203,N7204,N7205,N7206,N7207,
  N7208,N7209,N7210,N7211,N7212,N7213,N7214,N7215,N7216,N7217,N7218,N7219,N7220,
  N7221,N7222,N7223,N7224,N7225,N7226,N7227,N7228,N7229,N7230,N7231,N7232,N7233,
  N7234,N7235,N7236,N7237,N7238,N7239,N7240,N7241,N7242,N7243,N7244,N7245,N7246,N7247,
  N7248,N7249,N7250,N7251,N7252,N7253,N7254,N7255,N7256,N7257,N7258,N7259,N7260,
  N7261,N7262,N7263,N7264,N7265,N7266,N7267,N7268,N7269,N7270,N7271,N7272,N7273,
  N7274,N7275,N7276,N7277,N7278,N7279,N7280,N7281,N7282,N7283,N7284,N7285,N7286,N7287,
  N7288,N7289,N7290,N7291,N7292,N7293,N7294,N7295,N7296,N7297,N7298,N7299,N7300,
  N7301,N7302,N7303,N7304,N7305,N7306,N7307,N7308,N7309,N7310,N7311,N7312,N7313,
  N7314,N7315,N7316,N7317,N7318,N7319,N7320,N7321,N7322,N7323,N7324,N7325,N7326,N7327,
  N7328,N7329,N7330,N7331,N7332,N7333,N7334,N7335,N7336,N7337,N7338,N7339,N7340,
  N7341,N7342,N7343,N7344,N7345,N7346,N7347,N7348,N7349,N7350,N7351,N7352,N7353,
  N7354,N7355,N7356,N7357,N7358,N7359,N7360,N7361,N7362,N7363,N7364,N7365,N7366,N7367,
  N7368,N7369,N7370,N7371,N7372,N7373,N7374,N7375,N7376,N7377,N7378,N7379,N7380,
  N7381,N7382,N7383,N7384,N7385,N7386,N7387,N7388,N7389,N7390,N7391,N7392,N7393,
  N7394,N7395,N7396,N7397,N7398,N7399,N7400,N7401,N7402,N7403,N7404,N7405,N7406,N7407,
  N7408,N7409,N7410,N7411,N7412,N7413,N7414,N7415,N7416,N7417,N7418,N7419,N7420,
  N7421,N7422,N7423,N7424,N7425,N7426,N7427,N7428,N7429,N7430,N7431,N7432,N7433,
  N7434,N7435,N7436,N7437,N7438,N7439,N7440,N7441,N7442,N7443,N7444,N7445,N7446,N7447,
  N7448,N7449,N7450,N7451,N7452,N7453,N7454,N7455,N7456,N7457,N7458,N7459,N7460,
  N7461,N7462,N7463,N7464,N7465,N7466,N7467,N7468,N7469,N7470,N7471,N7472,N7473,
  N7474,N7475,N7476,N7477,N7478,N7479,N7480,N7481,N7482,N7483,N7484,N7485,N7486,N7487,
  N7488,N7489,N7490,N7491,N7492,N7493,N7494,N7495,N7496,N7497,N7498,N7499,N7500,
  N7501,N7502,N7503,N7504,N7505,N7506,N7507,N7508,N7509,N7510,N7511,N7512,N7513,
  N7514,N7515,N7516,N7517,N7518,N7519,N7520,N7521,N7522,N7523,N7524,N7525,N7526,N7527,
  N7528,N7529,N7530,N7531,N7532,N7533,N7534,N7535,N7536,N7537,N7538,N7539,N7540,
  N7541,N7542,N7543,N7544,N7545,N7546,N7547,N7548,N7549,N7550,N7551,N7552,N7553,
  N7554,N7555,N7556,N7557,N7558,N7559,N7560,N7561,N7562,N7563,N7564,N7565,N7566,N7567,
  N7568,N7569,N7570,N7571,N7572,N7573,N7574,N7575,N7576,N7577,N7578,N7579,N7580,
  N7581,N7582,N7583,N7584,N7585,N7586,N7587,N7588,N7589,N7590,N7591,N7592,N7593,
  N7594,N7595,N7596,N7597,N7598,N7599,N7600,N7601,N7602,N7603,N7604,N7605,N7606,N7607,
  N7608,N7609,N7610,N7611,N7612,N7613,N7614,N7615,N7616,N7617,N7618,N7619,N7620,
  N7621,N7622,N7623,N7624,N7625,N7626,N7627,N7628,N7629,N7630,N7631,N7632,N7633,
  N7634,N7635,N7636,N7637,N7638,N7639,N7640,N7641,N7642,N7643,N7644,N7645,N7646,N7647,
  N7648,N7649,N7650,N7651,N7652,N7653,N7654,N7655,N7656,N7657,N7658,N7659,N7660,
  N7661,N7662,N7663,N7664,N7665,N7666,N7667,N7668,N7669,N7670,N7671,N7672,N7673,
  N7674,N7675,N7676,N7677,N7678,N7679,N7680,N7681,N7682,N7683,N7684,N7685,N7686,N7687,
  N7688,N7689,N7690,N7691,N7692,N7693,N7694,N7695,N7696,N7697,N7698,N7699,N7700,
  N7701,N7702,N7703,N7704,N7705,N7706,N7707,N7708,N7709,N7710,N7711,N7712,N7713,
  N7714,N7715,N7716,N7717,N7718,N7719,N7720,N7721,N7722,N7723,N7724,N7725,N7726,N7727,
  N7728,N7729,N7730,N7731,N7732,N7733,N7734,N7735,N7736,N7737,N7738,N7739,N7740,
  N7741,N7742,N7743,N7744,N7745,N7746,N7747,N7748,N7749,N7750,N7751,N7752,N7753,
  N7754,N7755,N7756,N7757,N7758,N7759,N7760,N7761,N7762,N7763,N7764,N7765,N7766,N7767,
  N7768,N7769,N7770,N7771,N7772,N7773,N7774,N7775,N7776,N7777,N7778,N7779,N7780,
  N7781,N7782,N7783,N7784,N7785,N7786,N7787,N7788,N7789,N7790,N7791,N7792,N7793,
  N7794,N7795,N7796,N7797,N7798,N7799,N7800,N7801,N7802,N7803,N7804,N7805,N7806,N7807,
  N7808,N7809,N7810,N7811,N7812,N7813,N7814,N7815,N7816,N7817,N7818,N7819,N7820,
  N7821,N7822,N7823,N7824,N7825,N7826,N7827,N7828,N7829,N7830,N7831,N7832,N7833,
  N7834,N7835,N7836,N7837,N7838,N7839,N7840,N7841,N7842,N7843,N7844,N7845,N7846,N7847,
  N7848,N7849,N7850,N7851,N7852,N7853,N7854,N7855,N7856,N7857,N7858,N7859,N7860,
  N7861,N7862,N7863,N7864,N7865,N7866,N7867,N7868,N7869,N7870,N7871,N7872,N7873,
  N7874,N7875,N7876,N7877,N7878,N7879,N7880,N7881,N7882,N7883,N7884,N7885,N7886,N7887,
  N7888,N7889,N7890,N7891,N7892,N7893,N7894,N7895,N7896,N7897,N7898,N7899,N7900,
  N7901,N7902,N7903,N7904,N7905,N7906,N7907,N7908,N7909,N7910,N7911,N7912,N7913,
  N7914,N7915,N7916,N7917,N7918,N7919,N7920,N7921,N7922,N7923,N7924,N7925,N7926,N7927,
  N7928,N7929,N7930,N7931,N7932,N7933,N7934,N7935,N7936,N7937,N7938,N7939,N7940,
  N7941,N7942,N7943,N7944,N7945,N7946,N7947,N7948,N7949,N7950,N7951,N7952,N7953,
  N7954,N7955,N7956,N7957,N7958,N7959,N7960,N7961,N7962,N7963,N7964,N7965,N7966,N7967,
  N7968,N7969,N7970,N7971,N7972,N7973,N7974,N7975,N7976,N7977,N7978,N7979,N7980,
  N7981,N7982,N7983,N7984,N7985,N7986,N7987,N7988,N7989,N7990,N7991,N7992,N7993,
  N7994,N7995,N7996,N7997,N7998,N7999,N8000,N8001,N8002,N8003,N8004,N8005,N8006,N8007,
  N8008,N8009,N8010,N8011,N8012,N8013,N8014,N8015,N8016,N8017,N8018,N8019,N8020,
  N8021,N8022,N8023,N8024,N8025,N8026,N8027,N8028,N8029,N8030,N8031,N8032,N8033,
  N8034,N8035,N8036,N8037,N8038,N8039,N8040,N8041,N8042,N8043,N8044,N8045,N8046,N8047,
  N8048,N8049,N8050,N8051,N8052,N8053,N8054,N8055,N8056,N8057,N8058,N8059,N8060,
  N8061,N8062,N8063,N8064,N8065,N8066,N8067,N8068,N8069,N8070,N8071,N8072,N8073,
  N8074,N8075,N8076,N8077,N8078,N8079,N8080,N8081,N8082,N8083,N8084,N8085,N8086,N8087,
  N8088,N8089,N8090,N8091,N8092,N8093,N8094,N8095,N8096,N8097,N8098,N8099,N8100,
  N8101,N8102,N8103,N8104,N8105,N8106,N8107,N8108,N8109,N8110,N8111,N8112,N8113,
  N8114,N8115,N8116,N8117,N8118,N8119,N8120,N8121,N8122,N8123,N8124,N8125,N8126,N8127,
  N8128,N8129,N8130,N8131,N8132,N8133,N8134,N8135,N8136,N8137,N8138,N8139,N8140,
  N8141,N8142,N8143,N8144,N8145,N8146,N8147,N8148,N8149,N8150,N8151,N8152,N8153,
  N8154,N8155,N8156,N8157,N8158,N8159,N8160,N8161,N8162,N8163,N8164,N8165,N8166,N8167,
  N8168,N8169,N8170,N8171,N8172,N8173,N8174,N8175,N8176,N8177,N8178,N8179,N8180,
  N8181,N8182,N8183,N8184,N8185,N8186,N8187,N8188,N8189,N8190,N8191,N8192,N8193,
  N8194,N8195,N8196,N8197,N8198,N8199,N8200,N8201,N8202,N8203,N8204,N8205,N8206,N8207,
  N8208,N8209,N8210,N8211,N8212,N8213,N8214,N8215,N8216,N8217,N8218,N8219,N8220,
  N8221,N8222,N8223,N8224,N8225,N8226,N8227,N8228,N8229,N8230,N8231,N8232,N8233,
  N8234,N8235,N8236,N8237,N8238,N8239,N8240,N8241,N8242,N8243,N8244,N8245,N8246,N8247,
  N8248,N8249,N8250,N8251,N8252,N8253,N8254,N8255,N8256,N8257,N8258,N8259,N8260,
  N8261,N8262,N8263,N8264,N8265,N8266,N8267,N8268,N8269,N8270,N8271,N8272,N8273,
  N8274,N8275,N8276,N8277,N8278,N8279,N8280,N8281,N8282,N8283,N8284,N8285,N8286,N8287,
  N8288,N8289,N8290,N8291,N8292,N8293,N8294,N8295,N8296,N8297,N8298,N8299,N8300,
  N8301,N8302,N8303,N8304,N8305,N8306,N8307,N8308,N8309,N8310,N8311,N8312,N8313,
  N8314,N8315,N8316,N8317,N8318,N8319,N8320,N8321,N8322,N8323,N8324,N8325,N8326,N8327,
  N8328,N8329,N8330,N8331,N8332,N8333,N8334,N8335,N8336,N8337,N8338,N8339,N8340,
  N8341,N8342,N8343,N8344,N8345,N8346,N8347,N8348,N8349,N8350,N8351,N8352,N8353,
  N8354,N8355,N8356,N8357,N8358,N8359,N8360,N8361,N8362,N8363,N8364,N8365,N8366,N8367,
  N8368,N8369,N8370,N8371,N8372,N8373,N8374,N8375,N8376,N8377,N8378,N8379,N8380,
  N8381,N8382,N8383,N8384,N8385,N8386,N8387,N8388,N8389,N8390,N8391,N8392,N8393,
  N8394,N8395,N8396,N8397,N8398,N8399,N8400,N8401,N8402,N8403,N8404,N8405,N8406,N8407,
  N8408,N8409,N8410,N8411,N8412,N8413,N8414,N8415,N8416,N8417,N8418,N8419,N8420,
  N8421,N8422,N8423,N8424,N8425,N8426,N8427,N8428,N8429,N8430,N8431,N8432,N8433,
  N8434,N8435,N8436,N8437,N8438,N8439,N8440,N8441,N8442,N8443,N8444,N8445,N8446,N8447,
  N8448,N8449,N8450,N8451,N8452,N8453,N8454,N8455,N8456,N8457,N8458,N8459,N8460,
  N8461,N8462,N8463,N8464,N8465,N8466,N8467,N8468,N8469,N8470,N8471,N8472,N8473,
  N8474,N8475,N8476,N8477,N8478,N8479,N8480,N8481,N8482,N8483,N8484,N8485,N8486,N8487,
  N8488,N8489,N8490,N8491,N8492,N8493,N8494,N8495,N8496,N8497,N8498,N8499,N8500,
  N8501,N8502,N8503,N8504,N8505,N8506,N8507,N8508,N8509,N8510,N8511,N8512,N8513,
  N8514,N8515,N8516,N8517,N8518,N8519,N8520,N8521,N8522,N8523,N8524,N8525,N8526,N8527,
  N8528,N8529,N8530,N8531,N8532,N8533,N8534,N8535,N8536,N8537,N8538,N8539,N8540,
  N8541,N8542,N8543,N8544,N8545,N8546,N8547,N8548,N8549,N8550,N8551,N8552,N8553,
  N8554,N8555,N8556,N8557,N8558,N8559,N8560,N8561,N8562,N8563,N8564,N8565,N8566,N8567,
  N8568,N8569,N8570,N8571,N8572,N8573,N8574,N8575,N8576,N8577,N8578,N8579,N8580,
  N8581,N8582,N8583,N8584,N8585,N8586,N8587,N8588,N8589,N8590,N8591,N8592,N8593,
  N8594,N8595,N8596,N8597,N8598,N8599,N8600,N8601,N8602,N8603,N8604,N8605,N8606,N8607,
  N8608,N8609,N8610,N8611,N8612,N8613,N8614,N8615,N8616,N8617,N8618,N8619,N8620,
  N8621,N8622,N8623,N8624,N8625,N8626,N8627,N8628,N8629,N8630,N8631,N8632,N8633,
  N8634,N8635,N8636,N8637,N8638,N8639,N8640,N8641,N8642,N8643,N8644,N8645,N8646,N8647,
  N8648,N8649,N8650,N8651,N8652,N8653,N8654,N8655,N8656,N8657,N8658,N8659,N8660,
  N8661,N8662,N8663,N8664,N8665,N8666,N8667,N8668,N8669,N8670,N8671,N8672,N8673,
  N8674,N8675,N8676,N8677,N8678,N8679,N8680,N8681,N8682,N8683,N8684,N8685,N8686,N8687,
  N8688,N8689,N8690,N8691,N8692,N8693,N8694,N8695,N8696,N8697,N8698,N8699,N8700,
  N8701,N8702,N8703,N8704,N8705,N8706,N8707,N8708,N8709,N8710,N8711,N8712,N8713,
  N8714,N8715,N8716,N8717,N8718,N8719,N8720,N8721,N8722,N8723,N8724,N8725,N8726,N8727,
  N8728,N8729,N8730,N8731,N8732,N8733,N8734,N8735,N8736,N8737,N8738,N8739,N8740,
  N8741,N8742,N8743,N8744,N8745,N8746,N8747,N8748,N8749,N8750,N8751,N8752,N8753,
  N8754,N8755,N8756,N8757,N8758,N8759,N8760,N8761,N8762,N8763,N8764,N8765,N8766,N8767,
  N8768,N8769,N8770,N8771,N8772,N8773,N8774,N8775,N8776,N8777,N8778,N8779,N8780,
  N8781,N8782,N8783,N8784,N8785,N8786,N8787,N8788,N8789,N8790,N8791,N8792,N8793,
  N8794,N8795,N8796,N8797,N8798,N8799,N8800,N8801,N8802,N8803,N8804,N8805,N8806,N8807,
  N8808,N8809,N8810,N8811,N8812,N8813,N8814,N8815,N8816,N8817,N8818,N8819,N8820,
  N8821,N8822,N8823,N8824,N8825,N8826,N8827,N8828,N8829,N8830,N8831,N8832,N8833,
  N8834,N8835,N8836,N8837,N8838,N8839,N8840,N8841,N8842,N8843,N8844,N8845,N8846,N8847,
  N8848,N8849,N8850,N8851,N8852,N8853,N8854,N8855,N8856,N8857,N8858,N8859,N8860,
  N8861,N8862,N8863,N8864,N8865,N8866,N8867,N8868,N8869,N8870,N8871,N8872,N8873,
  N8874,N8875,N8876,N8877,N8878,N8879,N8880,N8881,N8882,N8883,N8884,N8885,N8886,N8887,
  N8888,N8889,N8890,N8891,N8892,N8893,N8894,N8895,N8896,N8897,N8898,N8899,N8900,
  N8901,N8902,N8903,N8904,N8905,N8906,N8907,N8908,N8909,N8910,N8911,N8912,N8913,
  N8914,N8915,N8916,N8917,N8918,N8919,N8920,N8921,N8922,N8923,N8924,N8925,N8926,N8927,
  N8928,N8929,N8930,N8931,N8932,N8933,N8934,N8935,N8936,N8937,N8938,N8939,N8940,
  N8941,N8942,N8943,N8944,N8945,N8946,N8947,N8948,N8949,N8950,N8951,N8952,N8953,
  N8954,N8955,N8956,N8957,N8958,N8959,N8960,N8961,N8962,N8963,N8964,N8965,N8966,N8967,
  N8968,N8969,N8970,N8971,N8972,N8973,N8974,N8975,N8976,N8977,N8978,N8979,N8980,
  N8981,N8982,N8983,N8984,N8985,N8986,N8987,N8988,N8989,N8990,N8991,N8992,N8993,
  N8994,N8995,N8996,N8997,N8998,N8999,N9000,N9001,N9002,N9003,N9004,N9005,N9006,N9007,
  N9008,N9009,N9010,N9011,N9012,N9013,N9014,N9015,N9016,N9017,N9018,N9019,N9020,
  N9021,N9022,N9023,N9024,N9025,N9026,N9027,N9028,N9029,N9030,N9031,N9032,N9033,
  N9034,N9035,N9036,N9037,N9038,N9039,N9040,N9041,N9042,N9043,N9044,N9045,N9046,N9047,
  N9048,N9049,N9050,N9051,N9052,N9053,N9054,N9055,N9056,N9057,N9058,N9059,N9060,
  N9061,N9062,N9063,N9064,N9065,N9066,N9067,N9068,N9069,N9070,N9071,N9072,N9073,
  N9074,N9075,N9076,N9077,N9078,N9079,N9080,N9081,N9082,N9083,N9084,N9085,N9086,N9087,
  N9088,N9089,N9090,N9091,N9092,N9093,N9094,N9095,N9096,N9097,N9098,N9099,N9100,
  N9101,N9102,N9103,N9104,N9105,N9106,N9107,N9108,N9109,N9110,N9111,N9112,N9113,
  N9114,N9115,N9116,N9117,N9118,N9119,N9120,N9121,N9122,N9123,N9124,N9125,N9126,N9127,
  N9128,N9129,N9130,N9131,N9132,N9133,N9134,N9135,N9136,N9137,N9138,N9139,N9140,
  N9141,N9142,N9143,N9144,N9145,N9146,N9147,N9148,N9149,N9150,N9151,N9152,N9153,
  N9154,N9155,N9156,N9157,N9158,N9159,N9160,N9161,N9162,N9163,N9164,N9165,N9166,N9167,
  N9168,N9169,N9170,N9171,N9172,N9173,N9174,N9175,N9176,N9177,N9178,N9179,N9180,
  N9181,N9182,N9183,N9184,N9185,N9186,N9187,N9188,N9189,N9190,N9191,N9192,N9193,
  N9194,N9195,N9196,N9197,N9198,N9199,N9200,N9201,N9202,N9203,N9204,N9205,N9206,N9207,
  N9208,N9209,N9210,N9211,N9212,N9213,N9214,N9215,N9216,N9217,N9218,N9219,N9220,
  N9221,N9222,N9223,N9224,N9225,N9226,N9227,N9228,N9229,N9230,N9231,N9232,N9233,
  N9234,N9235,N9236,N9237,N9238,N9239,N9240,N9241,N9242,N9243,N9244,N9245,N9246,N9247,
  N9248,N9249,N9250,N9251,N9252,N9253,N9254,N9255,N9256,N9257,N9258,N9259,N9260,
  N9261,N9262,N9263,N9264,N9265,N9266,N9267,N9268,N9269,N9270,N9271,N9272,N9273,
  N9274,N9275,N9276,N9277,N9278,N9279,N9280,N9281,N9282,N9283,N9284,N9285,N9286,N9287,
  N9288,N9289,N9290,N9291,N9292,N9293,N9294,N9295,N9296,N9297,N9298,N9299,N9300,
  N9301,N9302,N9303,N9304,N9305,N9306,N9307,N9308,N9309,N9310,N9311,N9312,N9313,
  N9314,N9315,N9316,N9317,N9318,N9319,N9320,N9321,N9322,N9323,N9324,N9325,N9326,N9327,
  N9328,N9329,N9330,N9331,N9332,N9333,N9334,N9335,N9336,N9337,N9338,N9339,N9340,
  N9341,N9342,N9343,N9344,N9345,N9346,N9347,N9348,N9349,N9350,N9351,N9352,N9353,
  N9354,N9355,N9356,N9357,N9358,N9359,N9360,N9361,N9362,N9363,N9364,N9365,N9366,N9367,
  N9368,N9369,N9370,N9371,N9372,N9373,N9374,N9375,N9376,N9377,N9378,N9379,N9380,
  N9381,N9382,N9383,N9384,N9385,N9386,N9387,N9388,N9389,N9390,N9391,N9392,N9393,
  N9394,N9395,N9396,N9397,N9398,N9399,N9400,N9401,N9402,N9403,N9404,N9405,N9406,N9407,
  N9408,N9409,N9410,N9411,N9412,N9413,N9414,N9415,N9416,N9417,N9418,N9419,N9420,
  N9421,N9422,N9423,N9424,N9425,N9426,N9427,N9428,N9429,N9430,N9431,N9432,N9433,
  N9434,N9435,N9436,N9437,N9438,N9439,N9440,N9441,N9442,N9443,N9444,N9445,N9446,N9447,
  N9448,N9449,N9450,N9451,N9452,N9453,N9454,N9455,N9456,N9457,N9458,N9459,N9460,
  N9461,N9462,N9463,N9464,N9465,N9466,N9467,N9468,N9469,N9470,N9471,N9472,N9473,
  N9474,N9475,N9476,N9477,N9478,N9479,N9480,N9481,N9482,N9483,N9484,N9485,N9486,N9487,
  N9488,N9489,N9490,N9491,N9492,N9493,N9494,N9495,N9496,N9497,N9498,N9499,N9500,
  N9501,N9502,N9503,N9504,N9505,N9506,N9507,N9508,N9509,N9510,N9511,N9512,N9513,
  N9514,N9515,N9516,N9517,N9518,N9519,N9520,N9521,N9522,N9523,N9524,N9525,N9526,N9527,
  N9528,N9529,N9530,N9531,N9532,N9533,N9534,N9535,N9536,N9537,N9538,N9539,N9540,
  N9541,N9542,N9543,N9544,N9545,N9546,N9547,N9548,N9549,N9550,N9551,N9552,N9553,
  N9554,N9555,N9556,N9557,N9558,N9559,N9560,N9561,N9562,N9563,N9564,N9565,N9566,N9567,
  N9568,N9569,N9570,N9571,N9572,N9573,N9574,N9575,N9576,N9577,N9578,N9579,N9580,
  N9581,N9582,N9583,N9584,N9585,N9586,N9587,N9588,N9589,N9590,N9591,N9592,N9593,
  N9594,N9595,N9596,N9597,N9598,N9599,N9600,N9601,N9602,N9603,N9604,N9605,N9606,N9607,
  N9608,N9609,N9610,N9611,N9612,N9613,N9614,N9615,N9616,N9617,N9618,N9619,N9620,
  N9621,N9622,N9623,N9624,N9625,N9626,N9627,N9628,N9629,N9630,N9631,N9632,N9633,
  N9634,N9635,N9636,N9637,N9638,N9639,N9640,N9641,N9642,N9643,N9644,N9645,N9646,N9647,
  N9648,N9649,N9650,N9651,N9652,N9653,N9654,N9655,N9656,N9657,N9658,N9659,N9660,
  N9661,N9662,N9663,N9664,N9665,N9666,N9667,N9668,N9669,N9670,N9671,N9672,N9673,
  N9674,N9675,N9676,N9677,N9678,N9679,N9680,N9681,N9682,N9683,N9684,N9685,N9686,N9687,
  N9688,N9689,N9690,N9691,N9692,N9693,N9694,N9695,N9696,N9697,N9698,N9699,N9700,
  N9701,N9702,N9703,N9704,N9705,N9706,N9707,N9708,N9709,N9710,N9711,N9712,N9713,
  N9714,N9715,N9716,N9717,N9718,N9719,N9720,N9721,N9722,N9723,N9724,N9725,N9726,N9727,
  N9728,N9729,N9730,N9731,N9732,N9733,N9734,N9735,N9736,N9737,N9738,N9739,N9740,
  N9741,N9742,N9743,N9744,N9745,N9746,N9747,N9748,N9749,N9750,N9751,N9752,N9753,
  N9754,N9755,N9756,N9757,N9758,N9759,N9760,N9761,N9762,N9763,N9764,N9765,N9766,N9767,
  N9768,N9769,N9770,N9771,N9772,N9773,N9774,N9775,N9776,N9777,N9778,N9779,N9780,
  N9781,N9782,N9783,N9784,N9785,N9786,N9787,N9788,N9789,N9790,N9791,N9792,N9793,
  N9794,N9795,N9796,N9797,N9798,N9799,N9800,N9801,N9802,N9803,N9804,N9805,N9806,N9807,
  N9808,N9809,N9810,N9811,N9812,N9813,N9814,N9815,N9816,N9817,N9818,N9819,N9820,
  N9821,N9822,N9823,N9824,N9825,N9826,N9827,N9828,N9829,N9830,N9831,N9832,N9833,
  N9834,N9835,N9836,N9837,N9838,N9839,N9840,N9841,N9842,N9843,N9844,N9845,N9846,N9847,
  N9848,N9849,N9850,N9851,N9852,N9853,N9854,N9855,N9856,N9857,N9858,N9859,N9860,
  N9861,N9862,N9863,N9864,N9865,N9866,N9867,N9868,N9869,N9870,N9871,N9872,N9873,
  N9874,N9875,N9876,N9877,N9878,N9879,N9880,N9881,N9882,N9883,N9884,N9885,N9886,N9887,
  N9888,N9889,N9890,N9891,N9892,N9893,N9894,N9895,N9896,N9897,N9898,N9899,N9900,
  N9901,N9902,N9903,N9904,N9905,N9906,N9907,N9908,N9909,N9910,N9911,N9912,N9913,
  N9914,N9915,N9916,N9917,N9918,N9919,N9920,N9921,N9922,N9923,N9924,N9925,N9926,N9927,
  N9928,N9929,N9930,N9931,N9932,N9933,N9934,N9935,N9936,N9937,N9938,N9939,N9940,
  N9941,N9942,N9943,N9944,N9945,N9946,N9947,N9948,N9949,N9950,N9951,N9952,N9953,
  N9954,N9955,N9956,N9957,N9958,N9959,N9960,N9961,N9962,N9963,N9964,N9965,N9966,N9967,
  N9968,N9969,N9970,N9971,N9972,N9973,N9974,N9975,N9976,N9977,N9978,N9979,N9980,
  N9981,N9982,N9983,N9984,N9985,N9986,N9987,N9988,N9989,N9990,N9991,N9992,N9993,
  N9994,N9995,N9996,N9997,N9998,N9999,N10000,N10001,N10002,N10003,N10004,N10005,
  N10006,N10007,N10008,N10009,N10010,N10011,N10012,N10013,N10014,N10015,N10016,N10017,
  N10018,N10019,N10020,N10021,N10022,N10023,N10024,N10025,N10026,N10027,N10028,
  N10029,N10030,N10031,N10032,N10033,N10034,N10035,N10036,N10037,N10038,N10039,N10040,
  N10041,N10042,N10043,N10044,N10045,N10046,N10047,N10048,N10049,N10050,N10051,
  N10052,N10053,N10054,N10055,N10056,N10057,N10058,N10059,N10060,N10061,N10062,N10063,
  N10064,N10065,N10066,N10067,N10068,N10069,N10070,N10071,N10072,N10073,N10074,
  N10075,N10076,N10077,N10078,N10079,N10080,N10081,N10082,N10083,N10084,N10085,
  N10086,N10087,N10088,N10089,N10090,N10091,N10092,N10093,N10094,N10095,N10096,N10097,
  N10098,N10099,N10100,N10101,N10102,N10103,N10104,N10105,N10106,N10107,N10108,
  N10109,N10110,N10111,N10112,N10113,N10114,N10115,N10116,N10117,N10118,N10119,N10120,
  N10121,N10122,N10123,N10124,N10125,N10126,N10127,N10128,N10129,N10130,N10131,
  N10132,N10133,N10134,N10135,N10136,N10137,N10138,N10139,N10140,N10141,N10142,N10143,
  N10144,N10145,N10146,N10147,N10148,N10149,N10150,N10151,N10152,N10153,N10154,
  N10155,N10156,N10157,N10158,N10159,N10160,N10161,N10162,N10163,N10164,N10165,
  N10166,N10167,N10168,N10169,N10170,N10171,N10172,N10173,N10174,N10175,N10176,N10177,
  N10178,N10179,N10180,N10181,N10182,N10183,N10184,N10185,N10186,N10187,N10188,
  N10189,N10190,N10191,N10192,N10193,N10194,N10195,N10196,N10197,N10198,N10199,N10200,
  N10201,N10202,N10203,N10204,N10205,N10206,N10207,N10208,N10209,N10210,N10211,
  N10212,N10213,N10214,N10215,N10216,N10217,N10218,N10219,N10220,N10221,N10222,N10223,
  N10224,N10225,N10226,N10227,N10228,N10229,N10230,N10231,N10232,N10233,N10234,
  N10235,N10236,N10237,N10238,N10239,N10240,N10241,N10242,N10243,N10244,N10245,
  N10246,N10247,N10248,N10249,N10250,N10251,N10252,N10253,N10254,N10255,N10256,N10257,
  N10258,N10259,N10260,N10261,N10262,N10263,N10264,N10265,N10266,N10267,N10268,
  N10269,N10270,N10271,N10272,N10273,N10274,N10275,N10276,N10277,N10278,N10279,N10280,
  N10281,N10282,N10283,N10284,N10285,N10286,N10287,N10288,N10289,N10290,N10291,
  N10292,N10293,N10294,N10295,N10296,N10297,N10298,N10299,N10300,N10301,N10302,N10303,
  N10304,N10305,N10306,N10307,N10308,N10309,N10310,N10311,N10312,N10313,N10314,
  N10315,N10316,N10317,N10318,N10319,N10320,N10321,N10322,N10323,N10324,N10325,
  N10326,N10327,N10328,N10329,N10330,N10331,N10332,N10333,N10334,N10335,N10336,N10337,
  N10338,N10339,N10340,N10341,N10342,N10343,N10344,N10345,N10346,N10347,N10348,
  N10349,N10350,N10351,N10352,N10353,N10354,N10355,N10356,N10357,N10358,N10359,N10360,
  N10361,N10362,N10363,N10364,N10365,N10366,N10367,N10368,N10369,N10370,N10371,
  N10372,N10373,N10374,N10375,N10376,N10377,N10378,N10379,N10380,N10381,N10382,N10383,
  N10384,N10385,N10386,N10387,N10388,N10389,N10390,N10391,N10392,N10393,N10394,
  N10395,N10396,N10397,N10398,N10399,N10400,N10401,N10402,N10403,N10404,N10405,
  N10406,N10407,N10408,N10409,N10410,N10411,N10412,N10413,N10414,N10415,N10416,N10417,
  N10418,N10419,N10420,N10421,N10422,N10423,N10424,N10425,N10426,N10427,N10428,
  N10429,N10430,N10431,N10432,N10433,N10434,N10435,N10436,N10437,N10438,N10439,N10440,
  N10441,N10442,N10443,N10444,N10445,N10446,N10447,N10448,N10449,N10450,N10451,
  N10452,N10453,N10454,N10455,N10456,N10457,N10458,N10459,N10460,N10461,N10462,N10463,
  N10464,N10465,N10466,N10467,N10468,N10469,N10470,N10471,N10472,N10473,N10474,
  N10475,N10476,N10477,N10478,N10479,N10480,N10481,N10482,N10483,N10484,N10485,
  N10486,N10487,N10488,N10489,N10490,N10491,N10492,N10493,N10494,N10495,N10496,N10497,
  N10498,N10499,N10500,N10501,N10502,N10503,N10504,N10505,N10506,N10507,N10508,
  N10509,N10510,N10511,N10512,N10513,N10514,N10515,N10516,N10517,N10518,N10519,N10520,
  N10521,N10522,N10523,N10524,N10525,N10526,N10527,N10528,N10529,N10530,N10531,
  N10532,N10533,N10534,N10535,N10536,N10537,N10538,N10539,N10540,N10541,N10542,N10543,
  N10544,N10545,N10546,N10547,N10548,N10549,N10550,N10551,N10552,N10553,N10554,
  N10555,N10556,N10557,N10558,N10559,N10560,N10561,N10562,N10563,N10564,N10565,
  N10566,N10567,N10568,N10569,N10570,N10571,N10572,N10573,N10574,N10575,N10576,N10577,
  N10578,N10579,N10580,N10581,N10582,N10583,N10584,N10585,N10586,N10587,N10588,
  N10589,N10590,N10591,N10592,N10593,N10594,N10595,N10596,N10597,N10598,N10599,N10600,
  N10601,N10602,N10603,N10604,N10605,N10606,N10607,N10608,N10609,N10610,N10611,
  N10612,N10613,N10614,N10615,N10616,N10617,N10618,N10619,N10620,N10621,N10622,N10623,
  N10624,N10625,N10626,N10627,N10628,N10629,N10630,N10631,N10632,N10633,N10634,
  N10635,N10636,N10637,N10638,N10639,N10640,N10641,N10642,N10643,N10644,N10645,
  N10646,N10647,N10648,N10649,N10650,N10651,N10652,N10653,N10654,N10655,N10656,N10657,
  N10658,N10659,N10660,N10661,N10662,N10663,N10664,N10665,N10666,N10667,N10668,
  N10669,N10670,N10671,N10672,N10673,N10674,N10675,N10676,N10677,N10678,N10679,N10680,
  N10681,N10682,N10683,N10684,N10685,N10686,N10687,N10688,N10689,N10690,N10691,
  N10692,N10693,N10694,N10695,N10696,N10697,N10698,N10699,N10700,N10701,N10702,N10703,
  N10704,N10705,N10706,N10707,N10708,N10709,N10710,N10711,N10712,N10713,N10714,
  N10715,N10716,N10717,N10718,N10719,N10720,N10721,N10722,N10723,N10724,N10725,
  N10726,N10727,N10728,N10729,N10730,N10731,N10732,N10733,N10734,N10735,N10736,N10737,
  N10738,N10739,N10740,N10741,N10742,N10743,N10744,N10745,N10746,N10747,N10748,
  N10749,N10750,N10751,N10752,N10753,N10754,N10755,N10756,N10757,N10758,N10759,N10760,
  N10761,N10762,N10763,N10764,N10765,N10766,N10767,N10768,N10769,N10770,N10771,
  N10772,N10773,N10774,N10775,N10776,N10777,N10778,N10779,N10780,N10781,N10782,N10783,
  N10784,N10785,N10786,N10787,N10788,N10789,N10790,N10791,N10792,N10793,N10794,
  N10795,N10796,N10797,N10798,N10799,N10800,N10801,N10802,N10803,N10804,N10805,
  N10806,N10807,N10808,N10809,N10810,N10811,N10812,N10813,N10814,N10815,N10816,N10817,
  N10818,N10819,N10820,N10821,N10822,N10823,N10824,N10825,N10826,N10827,N10828,
  N10829,N10830,N10831,N10832,N10833,N10834,N10835,N10836,N10837,N10838,N10839,N10840,
  N10841,N10842,N10843,N10844,N10845,N10846,N10847,N10848,N10849,N10850,N10851,
  N10852,N10853,N10854,N10855,N10856,N10857,N10858,N10859,N10860,N10861,N10862,N10863,
  N10864,N10865,N10866,N10867,N10868,N10869,N10870,N10871,N10872,N10873,N10874,
  N10875,N10876,N10877,N10878,N10879,N10880,N10881,N10882,N10883,N10884,N10885,
  N10886,N10887,N10888,N10889,N10890,N10891,N10892,N10893,N10894,N10895,N10896,N10897,
  N10898,N10899,N10900,N10901,N10902,N10903,N10904,N10905,N10906,N10907,N10908,
  N10909,N10910,N10911,N10912,N10913,N10914,N10915,N10916,N10917,N10918,N10919,N10920,
  N10921,N10922,N10923,N10924,N10925,N10926,N10927,N10928,N10929,N10930,N10931,
  N10932,N10933,N10934,N10935,N10936,N10937,N10938,N10939,N10940,N10941,N10942,N10943,
  N10944,N10945,N10946,N10947,N10948,N10949,N10950,N10951,N10952,N10953,N10954,
  N10955,N10956,N10957,N10958,N10959,N10960,N10961,N10962,N10963,N10964,N10965,
  N10966,N10967,N10968,N10969,N10970,N10971,N10972,N10973,N10974,N10975,N10976,N10977,
  N10978,N10979,N10980,N10981,N10982,N10983,N10984,N10985,N10986,N10987,N10988,
  N10989,N10990,N10991,N10992,N10993,N10994,N10995,N10996,N10997,N10998,N10999,N11000,
  N11001,N11002,N11003,N11004,N11005,N11006,N11007,N11008,N11009,N11010,N11011,
  N11012,N11013,N11014,N11015,N11016,N11017,N11018,N11019,N11020,N11021,N11022,N11023,
  N11024,N11025,N11026,N11027,N11028,N11029,N11030,N11031,N11032,N11033,N11034,
  N11035,N11036,N11037,N11038,N11039,N11040,N11041,N11042,N11043,N11044,N11045,
  N11046,N11047,N11048,N11049,N11050,N11051,N11052,N11053,N11054,N11055,N11056,N11057,
  N11058,N11059,N11060,N11061,N11062,N11063,N11064,N11065,N11066,N11067,N11068,
  N11069,N11070,N11071,N11072,N11073,N11074,N11075,N11076,N11077,N11078,N11079,N11080,
  N11081,N11082,N11083,N11084,N11085,N11086,N11087,N11088,N11089,N11090,N11091,
  N11092,N11093,N11094,N11095,N11096,N11097,N11098,N11099,N11100,N11101,N11102,N11103,
  N11104,N11105,N11106,N11107,N11108,N11109,N11110,N11111,N11112,N11113,N11114,
  N11115,N11116,N11117,N11118,N11119,N11120,N11121,N11122,N11123,N11124,N11125,
  N11126,N11127,N11128,N11129,N11130,N11131,N11132,N11133,N11134,N11135,N11136,N11137,
  N11138,N11139,N11140,N11141,N11142,N11143,N11144,N11145,N11146,N11147,N11148,
  N11149,N11150,N11151,N11152,N11153,N11154,N11155,N11156,N11157,N11158,N11159,N11160,
  N11161,N11162,N11163,N11164,N11165,N11166,N11167,N11168,N11169,N11170,N11171,
  N11172,N11173,N11174,N11175,N11176,N11177,N11178,N11179,N11180,N11181,N11182,N11183,
  N11184,N11185,N11186,N11187,N11188,N11189,N11190,N11191,N11192,N11193,N11194,
  N11195,N11196,N11197,N11198,N11199,N11200,N11201,N11202,N11203,N11204,N11205,
  N11206,N11207,N11208,N11209,N11210,N11211,N11212,N11213,N11214,N11215,N11216,N11217,
  N11218,N11219,N11220,N11221,N11222,N11223,N11224,N11225,N11226,N11227,N11228,
  N11229,N11230,N11231,N11232,N11233,N11234,N11235,N11236,N11237,N11238,N11239,N11240,
  N11241,N11242,N11243,N11244,N11245,N11246,N11247,N11248,N11249,N11250,N11251,
  N11252,N11253,N11254,N11255,N11256,N11257,N11258,N11259,N11260,N11261,N11262,N11263,
  N11264,N11265,N11266,N11267,N11268,N11269,N11270,N11271,N11272,N11273,N11274,
  N11275,N11276,N11277,N11278,N11279,N11280,N11281,N11282,N11283,N11284,N11285,
  N11286,N11287,N11288,N11289,N11290,N11291,N11292,N11293,N11294,N11295,N11296,N11297,
  N11298,N11299,N11300,N11301,N11302,N11303,N11304,N11305,N11306,N11307,N11308,
  N11309,N11310,N11311,N11312,N11313,N11314,N11315,N11316,N11317,N11318,N11319,N11320,
  N11321,N11322,N11323,N11324,N11325,N11326,N11327,N11328,N11329,N11330,N11331,
  N11332,N11333,N11334,N11335,N11336,N11337,N11338,N11339,N11340,N11341,N11342,N11343,
  N11344,N11345,N11346,N11347,N11348,N11349,N11350,N11351,N11352,N11353,N11354,
  N11355,N11356,N11357,N11358,N11359,N11360,N11361,N11362,N11363,N11364,N11365,
  N11366,N11367,N11368,N11369,N11370,N11371,N11372,N11373,N11374,N11375,N11376,N11377,
  N11378,N11379,N11380,N11381,N11382,N11383,N11384,N11385,N11386,N11387,N11388,
  N11389,N11390,N11391,N11392,N11393,N11394,N11395,N11396,N11397,N11398,N11399,N11400,
  N11401,N11402,N11403,N11404,N11405,N11406,N11407,N11408,N11409,N11410,N11411,
  N11412,N11413,N11414,N11415,N11416,N11417,N11418,N11419,N11420,N11421,N11422,N11423,
  N11424,N11425,N11426,N11427,N11428,N11429,N11430,N11431,N11432,N11433,N11434,
  N11435,N11436,N11437,N11438,N11439,N11440,N11441,N11442,N11443,N11444,N11445,
  N11446,N11447,N11448,N11449,N11450,N11451,N11452,N11453,N11454,N11455,N11456,N11457,
  N11458,N11459,N11460,N11461,N11462,N11463,N11464,N11465,N11466,N11467,N11468,
  N11469,N11470,N11471,N11472,N11473,N11474,N11475,N11476,N11477,N11478,N11479,N11480,
  N11481,N11482,N11483,N11484,N11485,N11486,N11487,N11488,N11489,N11490,N11491,
  N11492,N11493,N11494,N11495,N11496,N11497,N11498,N11499,N11500,N11501,N11502,N11503,
  N11504,N11505,N11506,N11507,N11508,N11509,N11510,N11511,N11512,N11513,N11514,
  N11515,N11516,N11517,N11518,N11519,N11520,N11521,N11522,N11523,N11524,N11525,
  N11526,N11527,N11528,N11529,N11530,N11531,N11532,N11533,N11534,N11535,N11536,N11537,
  N11538,N11539,N11540,N11541,N11542,N11543,N11544,N11545,N11546,N11547,N11548,
  N11549,N11550,N11551,N11552,N11553,N11554,N11555,N11556,N11557,N11558,N11559,N11560,
  N11561,N11562,N11563,N11564,N11565,N11566,N11567,N11568,N11569,N11570,N11571,
  N11572,N11573,N11574,N11575,N11576,N11577,N11578,N11579,N11580,N11581,N11582,N11583,
  N11584,N11585,N11586,N11587,N11588,N11589,N11590,N11591,N11592,N11593,N11594,
  N11595,N11596,N11597,N11598,N11599,N11600,N11601,N11602,N11603,N11604,N11605,
  N11606,N11607,N11608,N11609,N11610,N11611,N11612,N11613,N11614,N11615,N11616,N11617,
  N11618,N11619,N11620,N11621,N11622,N11623,N11624,N11625,N11626,N11627,N11628,
  N11629,N11630,N11631,N11632,N11633,N11634,N11635,N11636,N11637,N11638,N11639,N11640,
  N11641,N11642,N11643,N11644,N11645,N11646,N11647,N11648,N11649,N11650,N11651,
  N11652,N11653,N11654,N11655,N11656,N11657,N11658,N11659;
  reg [5:0] addr_r;
  reg [5119:0] mem;
  assign data_out[79] = (N163)? mem[79] : 
                        (N165)? mem[159] : 
                        (N167)? mem[239] : 
                        (N169)? mem[319] : 
                        (N171)? mem[399] : 
                        (N173)? mem[479] : 
                        (N175)? mem[559] : 
                        (N177)? mem[639] : 
                        (N179)? mem[719] : 
                        (N181)? mem[799] : 
                        (N183)? mem[879] : 
                        (N185)? mem[959] : 
                        (N187)? mem[1039] : 
                        (N189)? mem[1119] : 
                        (N191)? mem[1199] : 
                        (N193)? mem[1279] : 
                        (N195)? mem[1359] : 
                        (N197)? mem[1439] : 
                        (N199)? mem[1519] : 
                        (N201)? mem[1599] : 
                        (N203)? mem[1679] : 
                        (N205)? mem[1759] : 
                        (N207)? mem[1839] : 
                        (N209)? mem[1919] : 
                        (N211)? mem[1999] : 
                        (N213)? mem[2079] : 
                        (N215)? mem[2159] : 
                        (N217)? mem[2239] : 
                        (N219)? mem[2319] : 
                        (N221)? mem[2399] : 
                        (N223)? mem[2479] : 
                        (N225)? mem[2559] : 
                        (N164)? mem[2639] : 
                        (N166)? mem[2719] : 
                        (N168)? mem[2799] : 
                        (N170)? mem[2879] : 
                        (N172)? mem[2959] : 
                        (N174)? mem[3039] : 
                        (N176)? mem[3119] : 
                        (N178)? mem[3199] : 
                        (N180)? mem[3279] : 
                        (N182)? mem[3359] : 
                        (N184)? mem[3439] : 
                        (N186)? mem[3519] : 
                        (N188)? mem[3599] : 
                        (N190)? mem[3679] : 
                        (N192)? mem[3759] : 
                        (N194)? mem[3839] : 
                        (N196)? mem[3919] : 
                        (N198)? mem[3999] : 
                        (N200)? mem[4079] : 
                        (N202)? mem[4159] : 
                        (N204)? mem[4239] : 
                        (N206)? mem[4319] : 
                        (N208)? mem[4399] : 
                        (N210)? mem[4479] : 
                        (N212)? mem[4559] : 
                        (N214)? mem[4639] : 
                        (N216)? mem[4719] : 
                        (N218)? mem[4799] : 
                        (N220)? mem[4879] : 
                        (N222)? mem[4959] : 
                        (N224)? mem[5039] : 
                        (N226)? mem[5119] : 1'b0;
  assign data_out[78] = (N163)? mem[78] : 
                        (N165)? mem[158] : 
                        (N167)? mem[238] : 
                        (N169)? mem[318] : 
                        (N171)? mem[398] : 
                        (N173)? mem[478] : 
                        (N175)? mem[558] : 
                        (N177)? mem[638] : 
                        (N179)? mem[718] : 
                        (N181)? mem[798] : 
                        (N183)? mem[878] : 
                        (N185)? mem[958] : 
                        (N187)? mem[1038] : 
                        (N189)? mem[1118] : 
                        (N191)? mem[1198] : 
                        (N193)? mem[1278] : 
                        (N195)? mem[1358] : 
                        (N197)? mem[1438] : 
                        (N199)? mem[1518] : 
                        (N201)? mem[1598] : 
                        (N203)? mem[1678] : 
                        (N205)? mem[1758] : 
                        (N207)? mem[1838] : 
                        (N209)? mem[1918] : 
                        (N211)? mem[1998] : 
                        (N213)? mem[2078] : 
                        (N215)? mem[2158] : 
                        (N217)? mem[2238] : 
                        (N219)? mem[2318] : 
                        (N221)? mem[2398] : 
                        (N223)? mem[2478] : 
                        (N225)? mem[2558] : 
                        (N164)? mem[2638] : 
                        (N166)? mem[2718] : 
                        (N168)? mem[2798] : 
                        (N170)? mem[2878] : 
                        (N172)? mem[2958] : 
                        (N174)? mem[3038] : 
                        (N176)? mem[3118] : 
                        (N178)? mem[3198] : 
                        (N180)? mem[3278] : 
                        (N182)? mem[3358] : 
                        (N184)? mem[3438] : 
                        (N186)? mem[3518] : 
                        (N188)? mem[3598] : 
                        (N190)? mem[3678] : 
                        (N192)? mem[3758] : 
                        (N194)? mem[3838] : 
                        (N196)? mem[3918] : 
                        (N198)? mem[3998] : 
                        (N200)? mem[4078] : 
                        (N202)? mem[4158] : 
                        (N204)? mem[4238] : 
                        (N206)? mem[4318] : 
                        (N208)? mem[4398] : 
                        (N210)? mem[4478] : 
                        (N212)? mem[4558] : 
                        (N214)? mem[4638] : 
                        (N216)? mem[4718] : 
                        (N218)? mem[4798] : 
                        (N220)? mem[4878] : 
                        (N222)? mem[4958] : 
                        (N224)? mem[5038] : 
                        (N226)? mem[5118] : 1'b0;
  assign data_out[77] = (N163)? mem[77] : 
                        (N165)? mem[157] : 
                        (N167)? mem[237] : 
                        (N169)? mem[317] : 
                        (N171)? mem[397] : 
                        (N173)? mem[477] : 
                        (N175)? mem[557] : 
                        (N177)? mem[637] : 
                        (N179)? mem[717] : 
                        (N181)? mem[797] : 
                        (N183)? mem[877] : 
                        (N185)? mem[957] : 
                        (N187)? mem[1037] : 
                        (N189)? mem[1117] : 
                        (N191)? mem[1197] : 
                        (N193)? mem[1277] : 
                        (N195)? mem[1357] : 
                        (N197)? mem[1437] : 
                        (N199)? mem[1517] : 
                        (N201)? mem[1597] : 
                        (N203)? mem[1677] : 
                        (N205)? mem[1757] : 
                        (N207)? mem[1837] : 
                        (N209)? mem[1917] : 
                        (N211)? mem[1997] : 
                        (N213)? mem[2077] : 
                        (N215)? mem[2157] : 
                        (N217)? mem[2237] : 
                        (N219)? mem[2317] : 
                        (N221)? mem[2397] : 
                        (N223)? mem[2477] : 
                        (N225)? mem[2557] : 
                        (N164)? mem[2637] : 
                        (N166)? mem[2717] : 
                        (N168)? mem[2797] : 
                        (N170)? mem[2877] : 
                        (N172)? mem[2957] : 
                        (N174)? mem[3037] : 
                        (N176)? mem[3117] : 
                        (N178)? mem[3197] : 
                        (N180)? mem[3277] : 
                        (N182)? mem[3357] : 
                        (N184)? mem[3437] : 
                        (N186)? mem[3517] : 
                        (N188)? mem[3597] : 
                        (N190)? mem[3677] : 
                        (N192)? mem[3757] : 
                        (N194)? mem[3837] : 
                        (N196)? mem[3917] : 
                        (N198)? mem[3997] : 
                        (N200)? mem[4077] : 
                        (N202)? mem[4157] : 
                        (N204)? mem[4237] : 
                        (N206)? mem[4317] : 
                        (N208)? mem[4397] : 
                        (N210)? mem[4477] : 
                        (N212)? mem[4557] : 
                        (N214)? mem[4637] : 
                        (N216)? mem[4717] : 
                        (N218)? mem[4797] : 
                        (N220)? mem[4877] : 
                        (N222)? mem[4957] : 
                        (N224)? mem[5037] : 
                        (N226)? mem[5117] : 1'b0;
  assign data_out[76] = (N163)? mem[76] : 
                        (N165)? mem[156] : 
                        (N167)? mem[236] : 
                        (N169)? mem[316] : 
                        (N171)? mem[396] : 
                        (N173)? mem[476] : 
                        (N175)? mem[556] : 
                        (N177)? mem[636] : 
                        (N179)? mem[716] : 
                        (N181)? mem[796] : 
                        (N183)? mem[876] : 
                        (N185)? mem[956] : 
                        (N187)? mem[1036] : 
                        (N189)? mem[1116] : 
                        (N191)? mem[1196] : 
                        (N193)? mem[1276] : 
                        (N195)? mem[1356] : 
                        (N197)? mem[1436] : 
                        (N199)? mem[1516] : 
                        (N201)? mem[1596] : 
                        (N203)? mem[1676] : 
                        (N205)? mem[1756] : 
                        (N207)? mem[1836] : 
                        (N209)? mem[1916] : 
                        (N211)? mem[1996] : 
                        (N213)? mem[2076] : 
                        (N215)? mem[2156] : 
                        (N217)? mem[2236] : 
                        (N219)? mem[2316] : 
                        (N221)? mem[2396] : 
                        (N223)? mem[2476] : 
                        (N225)? mem[2556] : 
                        (N164)? mem[2636] : 
                        (N166)? mem[2716] : 
                        (N168)? mem[2796] : 
                        (N170)? mem[2876] : 
                        (N172)? mem[2956] : 
                        (N174)? mem[3036] : 
                        (N176)? mem[3116] : 
                        (N178)? mem[3196] : 
                        (N180)? mem[3276] : 
                        (N182)? mem[3356] : 
                        (N184)? mem[3436] : 
                        (N186)? mem[3516] : 
                        (N188)? mem[3596] : 
                        (N190)? mem[3676] : 
                        (N192)? mem[3756] : 
                        (N194)? mem[3836] : 
                        (N196)? mem[3916] : 
                        (N198)? mem[3996] : 
                        (N200)? mem[4076] : 
                        (N202)? mem[4156] : 
                        (N204)? mem[4236] : 
                        (N206)? mem[4316] : 
                        (N208)? mem[4396] : 
                        (N210)? mem[4476] : 
                        (N212)? mem[4556] : 
                        (N214)? mem[4636] : 
                        (N216)? mem[4716] : 
                        (N218)? mem[4796] : 
                        (N220)? mem[4876] : 
                        (N222)? mem[4956] : 
                        (N224)? mem[5036] : 
                        (N226)? mem[5116] : 1'b0;
  assign data_out[75] = (N163)? mem[75] : 
                        (N165)? mem[155] : 
                        (N167)? mem[235] : 
                        (N169)? mem[315] : 
                        (N171)? mem[395] : 
                        (N173)? mem[475] : 
                        (N175)? mem[555] : 
                        (N177)? mem[635] : 
                        (N179)? mem[715] : 
                        (N181)? mem[795] : 
                        (N183)? mem[875] : 
                        (N185)? mem[955] : 
                        (N187)? mem[1035] : 
                        (N189)? mem[1115] : 
                        (N191)? mem[1195] : 
                        (N193)? mem[1275] : 
                        (N195)? mem[1355] : 
                        (N197)? mem[1435] : 
                        (N199)? mem[1515] : 
                        (N201)? mem[1595] : 
                        (N203)? mem[1675] : 
                        (N205)? mem[1755] : 
                        (N207)? mem[1835] : 
                        (N209)? mem[1915] : 
                        (N211)? mem[1995] : 
                        (N213)? mem[2075] : 
                        (N215)? mem[2155] : 
                        (N217)? mem[2235] : 
                        (N219)? mem[2315] : 
                        (N221)? mem[2395] : 
                        (N223)? mem[2475] : 
                        (N225)? mem[2555] : 
                        (N164)? mem[2635] : 
                        (N166)? mem[2715] : 
                        (N168)? mem[2795] : 
                        (N170)? mem[2875] : 
                        (N172)? mem[2955] : 
                        (N174)? mem[3035] : 
                        (N176)? mem[3115] : 
                        (N178)? mem[3195] : 
                        (N180)? mem[3275] : 
                        (N182)? mem[3355] : 
                        (N184)? mem[3435] : 
                        (N186)? mem[3515] : 
                        (N188)? mem[3595] : 
                        (N190)? mem[3675] : 
                        (N192)? mem[3755] : 
                        (N194)? mem[3835] : 
                        (N196)? mem[3915] : 
                        (N198)? mem[3995] : 
                        (N200)? mem[4075] : 
                        (N202)? mem[4155] : 
                        (N204)? mem[4235] : 
                        (N206)? mem[4315] : 
                        (N208)? mem[4395] : 
                        (N210)? mem[4475] : 
                        (N212)? mem[4555] : 
                        (N214)? mem[4635] : 
                        (N216)? mem[4715] : 
                        (N218)? mem[4795] : 
                        (N220)? mem[4875] : 
                        (N222)? mem[4955] : 
                        (N224)? mem[5035] : 
                        (N226)? mem[5115] : 1'b0;
  assign data_out[74] = (N163)? mem[74] : 
                        (N165)? mem[154] : 
                        (N167)? mem[234] : 
                        (N169)? mem[314] : 
                        (N171)? mem[394] : 
                        (N173)? mem[474] : 
                        (N175)? mem[554] : 
                        (N177)? mem[634] : 
                        (N179)? mem[714] : 
                        (N181)? mem[794] : 
                        (N183)? mem[874] : 
                        (N185)? mem[954] : 
                        (N187)? mem[1034] : 
                        (N189)? mem[1114] : 
                        (N191)? mem[1194] : 
                        (N193)? mem[1274] : 
                        (N195)? mem[1354] : 
                        (N197)? mem[1434] : 
                        (N199)? mem[1514] : 
                        (N201)? mem[1594] : 
                        (N203)? mem[1674] : 
                        (N205)? mem[1754] : 
                        (N207)? mem[1834] : 
                        (N209)? mem[1914] : 
                        (N211)? mem[1994] : 
                        (N213)? mem[2074] : 
                        (N215)? mem[2154] : 
                        (N217)? mem[2234] : 
                        (N219)? mem[2314] : 
                        (N221)? mem[2394] : 
                        (N223)? mem[2474] : 
                        (N225)? mem[2554] : 
                        (N164)? mem[2634] : 
                        (N166)? mem[2714] : 
                        (N168)? mem[2794] : 
                        (N170)? mem[2874] : 
                        (N172)? mem[2954] : 
                        (N174)? mem[3034] : 
                        (N176)? mem[3114] : 
                        (N178)? mem[3194] : 
                        (N180)? mem[3274] : 
                        (N182)? mem[3354] : 
                        (N184)? mem[3434] : 
                        (N186)? mem[3514] : 
                        (N188)? mem[3594] : 
                        (N190)? mem[3674] : 
                        (N192)? mem[3754] : 
                        (N194)? mem[3834] : 
                        (N196)? mem[3914] : 
                        (N198)? mem[3994] : 
                        (N200)? mem[4074] : 
                        (N202)? mem[4154] : 
                        (N204)? mem[4234] : 
                        (N206)? mem[4314] : 
                        (N208)? mem[4394] : 
                        (N210)? mem[4474] : 
                        (N212)? mem[4554] : 
                        (N214)? mem[4634] : 
                        (N216)? mem[4714] : 
                        (N218)? mem[4794] : 
                        (N220)? mem[4874] : 
                        (N222)? mem[4954] : 
                        (N224)? mem[5034] : 
                        (N226)? mem[5114] : 1'b0;
  assign data_out[73] = (N163)? mem[73] : 
                        (N165)? mem[153] : 
                        (N167)? mem[233] : 
                        (N169)? mem[313] : 
                        (N171)? mem[393] : 
                        (N173)? mem[473] : 
                        (N175)? mem[553] : 
                        (N177)? mem[633] : 
                        (N179)? mem[713] : 
                        (N181)? mem[793] : 
                        (N183)? mem[873] : 
                        (N185)? mem[953] : 
                        (N187)? mem[1033] : 
                        (N189)? mem[1113] : 
                        (N191)? mem[1193] : 
                        (N193)? mem[1273] : 
                        (N195)? mem[1353] : 
                        (N197)? mem[1433] : 
                        (N199)? mem[1513] : 
                        (N201)? mem[1593] : 
                        (N203)? mem[1673] : 
                        (N205)? mem[1753] : 
                        (N207)? mem[1833] : 
                        (N209)? mem[1913] : 
                        (N211)? mem[1993] : 
                        (N213)? mem[2073] : 
                        (N215)? mem[2153] : 
                        (N217)? mem[2233] : 
                        (N219)? mem[2313] : 
                        (N221)? mem[2393] : 
                        (N223)? mem[2473] : 
                        (N225)? mem[2553] : 
                        (N164)? mem[2633] : 
                        (N166)? mem[2713] : 
                        (N168)? mem[2793] : 
                        (N170)? mem[2873] : 
                        (N172)? mem[2953] : 
                        (N174)? mem[3033] : 
                        (N176)? mem[3113] : 
                        (N178)? mem[3193] : 
                        (N180)? mem[3273] : 
                        (N182)? mem[3353] : 
                        (N184)? mem[3433] : 
                        (N186)? mem[3513] : 
                        (N188)? mem[3593] : 
                        (N190)? mem[3673] : 
                        (N192)? mem[3753] : 
                        (N194)? mem[3833] : 
                        (N196)? mem[3913] : 
                        (N198)? mem[3993] : 
                        (N200)? mem[4073] : 
                        (N202)? mem[4153] : 
                        (N204)? mem[4233] : 
                        (N206)? mem[4313] : 
                        (N208)? mem[4393] : 
                        (N210)? mem[4473] : 
                        (N212)? mem[4553] : 
                        (N214)? mem[4633] : 
                        (N216)? mem[4713] : 
                        (N218)? mem[4793] : 
                        (N220)? mem[4873] : 
                        (N222)? mem[4953] : 
                        (N224)? mem[5033] : 
                        (N226)? mem[5113] : 1'b0;
  assign data_out[72] = (N163)? mem[72] : 
                        (N165)? mem[152] : 
                        (N167)? mem[232] : 
                        (N169)? mem[312] : 
                        (N171)? mem[392] : 
                        (N173)? mem[472] : 
                        (N175)? mem[552] : 
                        (N177)? mem[632] : 
                        (N179)? mem[712] : 
                        (N181)? mem[792] : 
                        (N183)? mem[872] : 
                        (N185)? mem[952] : 
                        (N187)? mem[1032] : 
                        (N189)? mem[1112] : 
                        (N191)? mem[1192] : 
                        (N193)? mem[1272] : 
                        (N195)? mem[1352] : 
                        (N197)? mem[1432] : 
                        (N199)? mem[1512] : 
                        (N201)? mem[1592] : 
                        (N203)? mem[1672] : 
                        (N205)? mem[1752] : 
                        (N207)? mem[1832] : 
                        (N209)? mem[1912] : 
                        (N211)? mem[1992] : 
                        (N213)? mem[2072] : 
                        (N215)? mem[2152] : 
                        (N217)? mem[2232] : 
                        (N219)? mem[2312] : 
                        (N221)? mem[2392] : 
                        (N223)? mem[2472] : 
                        (N225)? mem[2552] : 
                        (N164)? mem[2632] : 
                        (N166)? mem[2712] : 
                        (N168)? mem[2792] : 
                        (N170)? mem[2872] : 
                        (N172)? mem[2952] : 
                        (N174)? mem[3032] : 
                        (N176)? mem[3112] : 
                        (N178)? mem[3192] : 
                        (N180)? mem[3272] : 
                        (N182)? mem[3352] : 
                        (N184)? mem[3432] : 
                        (N186)? mem[3512] : 
                        (N188)? mem[3592] : 
                        (N190)? mem[3672] : 
                        (N192)? mem[3752] : 
                        (N194)? mem[3832] : 
                        (N196)? mem[3912] : 
                        (N198)? mem[3992] : 
                        (N200)? mem[4072] : 
                        (N202)? mem[4152] : 
                        (N204)? mem[4232] : 
                        (N206)? mem[4312] : 
                        (N208)? mem[4392] : 
                        (N210)? mem[4472] : 
                        (N212)? mem[4552] : 
                        (N214)? mem[4632] : 
                        (N216)? mem[4712] : 
                        (N218)? mem[4792] : 
                        (N220)? mem[4872] : 
                        (N222)? mem[4952] : 
                        (N224)? mem[5032] : 
                        (N226)? mem[5112] : 1'b0;
  assign data_out[71] = (N163)? mem[71] : 
                        (N165)? mem[151] : 
                        (N167)? mem[231] : 
                        (N169)? mem[311] : 
                        (N171)? mem[391] : 
                        (N173)? mem[471] : 
                        (N175)? mem[551] : 
                        (N177)? mem[631] : 
                        (N179)? mem[711] : 
                        (N181)? mem[791] : 
                        (N183)? mem[871] : 
                        (N185)? mem[951] : 
                        (N187)? mem[1031] : 
                        (N189)? mem[1111] : 
                        (N191)? mem[1191] : 
                        (N193)? mem[1271] : 
                        (N195)? mem[1351] : 
                        (N197)? mem[1431] : 
                        (N199)? mem[1511] : 
                        (N201)? mem[1591] : 
                        (N203)? mem[1671] : 
                        (N205)? mem[1751] : 
                        (N207)? mem[1831] : 
                        (N209)? mem[1911] : 
                        (N211)? mem[1991] : 
                        (N213)? mem[2071] : 
                        (N215)? mem[2151] : 
                        (N217)? mem[2231] : 
                        (N219)? mem[2311] : 
                        (N221)? mem[2391] : 
                        (N223)? mem[2471] : 
                        (N225)? mem[2551] : 
                        (N164)? mem[2631] : 
                        (N166)? mem[2711] : 
                        (N168)? mem[2791] : 
                        (N170)? mem[2871] : 
                        (N172)? mem[2951] : 
                        (N174)? mem[3031] : 
                        (N176)? mem[3111] : 
                        (N178)? mem[3191] : 
                        (N180)? mem[3271] : 
                        (N182)? mem[3351] : 
                        (N184)? mem[3431] : 
                        (N186)? mem[3511] : 
                        (N188)? mem[3591] : 
                        (N190)? mem[3671] : 
                        (N192)? mem[3751] : 
                        (N194)? mem[3831] : 
                        (N196)? mem[3911] : 
                        (N198)? mem[3991] : 
                        (N200)? mem[4071] : 
                        (N202)? mem[4151] : 
                        (N204)? mem[4231] : 
                        (N206)? mem[4311] : 
                        (N208)? mem[4391] : 
                        (N210)? mem[4471] : 
                        (N212)? mem[4551] : 
                        (N214)? mem[4631] : 
                        (N216)? mem[4711] : 
                        (N218)? mem[4791] : 
                        (N220)? mem[4871] : 
                        (N222)? mem[4951] : 
                        (N224)? mem[5031] : 
                        (N226)? mem[5111] : 1'b0;
  assign data_out[70] = (N163)? mem[70] : 
                        (N165)? mem[150] : 
                        (N167)? mem[230] : 
                        (N169)? mem[310] : 
                        (N171)? mem[390] : 
                        (N173)? mem[470] : 
                        (N175)? mem[550] : 
                        (N177)? mem[630] : 
                        (N179)? mem[710] : 
                        (N181)? mem[790] : 
                        (N183)? mem[870] : 
                        (N185)? mem[950] : 
                        (N187)? mem[1030] : 
                        (N189)? mem[1110] : 
                        (N191)? mem[1190] : 
                        (N193)? mem[1270] : 
                        (N195)? mem[1350] : 
                        (N197)? mem[1430] : 
                        (N199)? mem[1510] : 
                        (N201)? mem[1590] : 
                        (N203)? mem[1670] : 
                        (N205)? mem[1750] : 
                        (N207)? mem[1830] : 
                        (N209)? mem[1910] : 
                        (N211)? mem[1990] : 
                        (N213)? mem[2070] : 
                        (N215)? mem[2150] : 
                        (N217)? mem[2230] : 
                        (N219)? mem[2310] : 
                        (N221)? mem[2390] : 
                        (N223)? mem[2470] : 
                        (N225)? mem[2550] : 
                        (N164)? mem[2630] : 
                        (N166)? mem[2710] : 
                        (N168)? mem[2790] : 
                        (N170)? mem[2870] : 
                        (N172)? mem[2950] : 
                        (N174)? mem[3030] : 
                        (N176)? mem[3110] : 
                        (N178)? mem[3190] : 
                        (N180)? mem[3270] : 
                        (N182)? mem[3350] : 
                        (N184)? mem[3430] : 
                        (N186)? mem[3510] : 
                        (N188)? mem[3590] : 
                        (N190)? mem[3670] : 
                        (N192)? mem[3750] : 
                        (N194)? mem[3830] : 
                        (N196)? mem[3910] : 
                        (N198)? mem[3990] : 
                        (N200)? mem[4070] : 
                        (N202)? mem[4150] : 
                        (N204)? mem[4230] : 
                        (N206)? mem[4310] : 
                        (N208)? mem[4390] : 
                        (N210)? mem[4470] : 
                        (N212)? mem[4550] : 
                        (N214)? mem[4630] : 
                        (N216)? mem[4710] : 
                        (N218)? mem[4790] : 
                        (N220)? mem[4870] : 
                        (N222)? mem[4950] : 
                        (N224)? mem[5030] : 
                        (N226)? mem[5110] : 1'b0;
  assign data_out[69] = (N163)? mem[69] : 
                        (N165)? mem[149] : 
                        (N167)? mem[229] : 
                        (N169)? mem[309] : 
                        (N171)? mem[389] : 
                        (N173)? mem[469] : 
                        (N175)? mem[549] : 
                        (N177)? mem[629] : 
                        (N179)? mem[709] : 
                        (N181)? mem[789] : 
                        (N183)? mem[869] : 
                        (N185)? mem[949] : 
                        (N187)? mem[1029] : 
                        (N189)? mem[1109] : 
                        (N191)? mem[1189] : 
                        (N193)? mem[1269] : 
                        (N195)? mem[1349] : 
                        (N197)? mem[1429] : 
                        (N199)? mem[1509] : 
                        (N201)? mem[1589] : 
                        (N203)? mem[1669] : 
                        (N205)? mem[1749] : 
                        (N207)? mem[1829] : 
                        (N209)? mem[1909] : 
                        (N211)? mem[1989] : 
                        (N213)? mem[2069] : 
                        (N215)? mem[2149] : 
                        (N217)? mem[2229] : 
                        (N219)? mem[2309] : 
                        (N221)? mem[2389] : 
                        (N223)? mem[2469] : 
                        (N225)? mem[2549] : 
                        (N164)? mem[2629] : 
                        (N166)? mem[2709] : 
                        (N168)? mem[2789] : 
                        (N170)? mem[2869] : 
                        (N172)? mem[2949] : 
                        (N174)? mem[3029] : 
                        (N176)? mem[3109] : 
                        (N178)? mem[3189] : 
                        (N180)? mem[3269] : 
                        (N182)? mem[3349] : 
                        (N184)? mem[3429] : 
                        (N186)? mem[3509] : 
                        (N188)? mem[3589] : 
                        (N190)? mem[3669] : 
                        (N192)? mem[3749] : 
                        (N194)? mem[3829] : 
                        (N196)? mem[3909] : 
                        (N198)? mem[3989] : 
                        (N200)? mem[4069] : 
                        (N202)? mem[4149] : 
                        (N204)? mem[4229] : 
                        (N206)? mem[4309] : 
                        (N208)? mem[4389] : 
                        (N210)? mem[4469] : 
                        (N212)? mem[4549] : 
                        (N214)? mem[4629] : 
                        (N216)? mem[4709] : 
                        (N218)? mem[4789] : 
                        (N220)? mem[4869] : 
                        (N222)? mem[4949] : 
                        (N224)? mem[5029] : 
                        (N226)? mem[5109] : 1'b0;
  assign data_out[68] = (N163)? mem[68] : 
                        (N165)? mem[148] : 
                        (N167)? mem[228] : 
                        (N169)? mem[308] : 
                        (N171)? mem[388] : 
                        (N173)? mem[468] : 
                        (N175)? mem[548] : 
                        (N177)? mem[628] : 
                        (N179)? mem[708] : 
                        (N181)? mem[788] : 
                        (N183)? mem[868] : 
                        (N185)? mem[948] : 
                        (N187)? mem[1028] : 
                        (N189)? mem[1108] : 
                        (N191)? mem[1188] : 
                        (N193)? mem[1268] : 
                        (N195)? mem[1348] : 
                        (N197)? mem[1428] : 
                        (N199)? mem[1508] : 
                        (N201)? mem[1588] : 
                        (N203)? mem[1668] : 
                        (N205)? mem[1748] : 
                        (N207)? mem[1828] : 
                        (N209)? mem[1908] : 
                        (N211)? mem[1988] : 
                        (N213)? mem[2068] : 
                        (N215)? mem[2148] : 
                        (N217)? mem[2228] : 
                        (N219)? mem[2308] : 
                        (N221)? mem[2388] : 
                        (N223)? mem[2468] : 
                        (N225)? mem[2548] : 
                        (N164)? mem[2628] : 
                        (N166)? mem[2708] : 
                        (N168)? mem[2788] : 
                        (N170)? mem[2868] : 
                        (N172)? mem[2948] : 
                        (N174)? mem[3028] : 
                        (N176)? mem[3108] : 
                        (N178)? mem[3188] : 
                        (N180)? mem[3268] : 
                        (N182)? mem[3348] : 
                        (N184)? mem[3428] : 
                        (N186)? mem[3508] : 
                        (N188)? mem[3588] : 
                        (N190)? mem[3668] : 
                        (N192)? mem[3748] : 
                        (N194)? mem[3828] : 
                        (N196)? mem[3908] : 
                        (N198)? mem[3988] : 
                        (N200)? mem[4068] : 
                        (N202)? mem[4148] : 
                        (N204)? mem[4228] : 
                        (N206)? mem[4308] : 
                        (N208)? mem[4388] : 
                        (N210)? mem[4468] : 
                        (N212)? mem[4548] : 
                        (N214)? mem[4628] : 
                        (N216)? mem[4708] : 
                        (N218)? mem[4788] : 
                        (N220)? mem[4868] : 
                        (N222)? mem[4948] : 
                        (N224)? mem[5028] : 
                        (N226)? mem[5108] : 1'b0;
  assign data_out[67] = (N163)? mem[67] : 
                        (N165)? mem[147] : 
                        (N167)? mem[227] : 
                        (N169)? mem[307] : 
                        (N171)? mem[387] : 
                        (N173)? mem[467] : 
                        (N175)? mem[547] : 
                        (N177)? mem[627] : 
                        (N179)? mem[707] : 
                        (N181)? mem[787] : 
                        (N183)? mem[867] : 
                        (N185)? mem[947] : 
                        (N187)? mem[1027] : 
                        (N189)? mem[1107] : 
                        (N191)? mem[1187] : 
                        (N193)? mem[1267] : 
                        (N195)? mem[1347] : 
                        (N197)? mem[1427] : 
                        (N199)? mem[1507] : 
                        (N201)? mem[1587] : 
                        (N203)? mem[1667] : 
                        (N205)? mem[1747] : 
                        (N207)? mem[1827] : 
                        (N209)? mem[1907] : 
                        (N211)? mem[1987] : 
                        (N213)? mem[2067] : 
                        (N215)? mem[2147] : 
                        (N217)? mem[2227] : 
                        (N219)? mem[2307] : 
                        (N221)? mem[2387] : 
                        (N223)? mem[2467] : 
                        (N225)? mem[2547] : 
                        (N164)? mem[2627] : 
                        (N166)? mem[2707] : 
                        (N168)? mem[2787] : 
                        (N170)? mem[2867] : 
                        (N172)? mem[2947] : 
                        (N174)? mem[3027] : 
                        (N176)? mem[3107] : 
                        (N178)? mem[3187] : 
                        (N180)? mem[3267] : 
                        (N182)? mem[3347] : 
                        (N184)? mem[3427] : 
                        (N186)? mem[3507] : 
                        (N188)? mem[3587] : 
                        (N190)? mem[3667] : 
                        (N192)? mem[3747] : 
                        (N194)? mem[3827] : 
                        (N196)? mem[3907] : 
                        (N198)? mem[3987] : 
                        (N200)? mem[4067] : 
                        (N202)? mem[4147] : 
                        (N204)? mem[4227] : 
                        (N206)? mem[4307] : 
                        (N208)? mem[4387] : 
                        (N210)? mem[4467] : 
                        (N212)? mem[4547] : 
                        (N214)? mem[4627] : 
                        (N216)? mem[4707] : 
                        (N218)? mem[4787] : 
                        (N220)? mem[4867] : 
                        (N222)? mem[4947] : 
                        (N224)? mem[5027] : 
                        (N226)? mem[5107] : 1'b0;
  assign data_out[66] = (N163)? mem[66] : 
                        (N165)? mem[146] : 
                        (N167)? mem[226] : 
                        (N169)? mem[306] : 
                        (N171)? mem[386] : 
                        (N173)? mem[466] : 
                        (N175)? mem[546] : 
                        (N177)? mem[626] : 
                        (N179)? mem[706] : 
                        (N181)? mem[786] : 
                        (N183)? mem[866] : 
                        (N185)? mem[946] : 
                        (N187)? mem[1026] : 
                        (N189)? mem[1106] : 
                        (N191)? mem[1186] : 
                        (N193)? mem[1266] : 
                        (N195)? mem[1346] : 
                        (N197)? mem[1426] : 
                        (N199)? mem[1506] : 
                        (N201)? mem[1586] : 
                        (N203)? mem[1666] : 
                        (N205)? mem[1746] : 
                        (N207)? mem[1826] : 
                        (N209)? mem[1906] : 
                        (N211)? mem[1986] : 
                        (N213)? mem[2066] : 
                        (N215)? mem[2146] : 
                        (N217)? mem[2226] : 
                        (N219)? mem[2306] : 
                        (N221)? mem[2386] : 
                        (N223)? mem[2466] : 
                        (N225)? mem[2546] : 
                        (N164)? mem[2626] : 
                        (N166)? mem[2706] : 
                        (N168)? mem[2786] : 
                        (N170)? mem[2866] : 
                        (N172)? mem[2946] : 
                        (N174)? mem[3026] : 
                        (N176)? mem[3106] : 
                        (N178)? mem[3186] : 
                        (N180)? mem[3266] : 
                        (N182)? mem[3346] : 
                        (N184)? mem[3426] : 
                        (N186)? mem[3506] : 
                        (N188)? mem[3586] : 
                        (N190)? mem[3666] : 
                        (N192)? mem[3746] : 
                        (N194)? mem[3826] : 
                        (N196)? mem[3906] : 
                        (N198)? mem[3986] : 
                        (N200)? mem[4066] : 
                        (N202)? mem[4146] : 
                        (N204)? mem[4226] : 
                        (N206)? mem[4306] : 
                        (N208)? mem[4386] : 
                        (N210)? mem[4466] : 
                        (N212)? mem[4546] : 
                        (N214)? mem[4626] : 
                        (N216)? mem[4706] : 
                        (N218)? mem[4786] : 
                        (N220)? mem[4866] : 
                        (N222)? mem[4946] : 
                        (N224)? mem[5026] : 
                        (N226)? mem[5106] : 1'b0;
  assign data_out[65] = (N163)? mem[65] : 
                        (N165)? mem[145] : 
                        (N167)? mem[225] : 
                        (N169)? mem[305] : 
                        (N171)? mem[385] : 
                        (N173)? mem[465] : 
                        (N175)? mem[545] : 
                        (N177)? mem[625] : 
                        (N179)? mem[705] : 
                        (N181)? mem[785] : 
                        (N183)? mem[865] : 
                        (N185)? mem[945] : 
                        (N187)? mem[1025] : 
                        (N189)? mem[1105] : 
                        (N191)? mem[1185] : 
                        (N193)? mem[1265] : 
                        (N195)? mem[1345] : 
                        (N197)? mem[1425] : 
                        (N199)? mem[1505] : 
                        (N201)? mem[1585] : 
                        (N203)? mem[1665] : 
                        (N205)? mem[1745] : 
                        (N207)? mem[1825] : 
                        (N209)? mem[1905] : 
                        (N211)? mem[1985] : 
                        (N213)? mem[2065] : 
                        (N215)? mem[2145] : 
                        (N217)? mem[2225] : 
                        (N219)? mem[2305] : 
                        (N221)? mem[2385] : 
                        (N223)? mem[2465] : 
                        (N225)? mem[2545] : 
                        (N164)? mem[2625] : 
                        (N166)? mem[2705] : 
                        (N168)? mem[2785] : 
                        (N170)? mem[2865] : 
                        (N172)? mem[2945] : 
                        (N174)? mem[3025] : 
                        (N176)? mem[3105] : 
                        (N178)? mem[3185] : 
                        (N180)? mem[3265] : 
                        (N182)? mem[3345] : 
                        (N184)? mem[3425] : 
                        (N186)? mem[3505] : 
                        (N188)? mem[3585] : 
                        (N190)? mem[3665] : 
                        (N192)? mem[3745] : 
                        (N194)? mem[3825] : 
                        (N196)? mem[3905] : 
                        (N198)? mem[3985] : 
                        (N200)? mem[4065] : 
                        (N202)? mem[4145] : 
                        (N204)? mem[4225] : 
                        (N206)? mem[4305] : 
                        (N208)? mem[4385] : 
                        (N210)? mem[4465] : 
                        (N212)? mem[4545] : 
                        (N214)? mem[4625] : 
                        (N216)? mem[4705] : 
                        (N218)? mem[4785] : 
                        (N220)? mem[4865] : 
                        (N222)? mem[4945] : 
                        (N224)? mem[5025] : 
                        (N226)? mem[5105] : 1'b0;
  assign data_out[64] = (N163)? mem[64] : 
                        (N165)? mem[144] : 
                        (N167)? mem[224] : 
                        (N169)? mem[304] : 
                        (N171)? mem[384] : 
                        (N173)? mem[464] : 
                        (N175)? mem[544] : 
                        (N177)? mem[624] : 
                        (N179)? mem[704] : 
                        (N181)? mem[784] : 
                        (N183)? mem[864] : 
                        (N185)? mem[944] : 
                        (N187)? mem[1024] : 
                        (N189)? mem[1104] : 
                        (N191)? mem[1184] : 
                        (N193)? mem[1264] : 
                        (N195)? mem[1344] : 
                        (N197)? mem[1424] : 
                        (N199)? mem[1504] : 
                        (N201)? mem[1584] : 
                        (N203)? mem[1664] : 
                        (N205)? mem[1744] : 
                        (N207)? mem[1824] : 
                        (N209)? mem[1904] : 
                        (N211)? mem[1984] : 
                        (N213)? mem[2064] : 
                        (N215)? mem[2144] : 
                        (N217)? mem[2224] : 
                        (N219)? mem[2304] : 
                        (N221)? mem[2384] : 
                        (N223)? mem[2464] : 
                        (N225)? mem[2544] : 
                        (N164)? mem[2624] : 
                        (N166)? mem[2704] : 
                        (N168)? mem[2784] : 
                        (N170)? mem[2864] : 
                        (N172)? mem[2944] : 
                        (N174)? mem[3024] : 
                        (N176)? mem[3104] : 
                        (N178)? mem[3184] : 
                        (N180)? mem[3264] : 
                        (N182)? mem[3344] : 
                        (N184)? mem[3424] : 
                        (N186)? mem[3504] : 
                        (N188)? mem[3584] : 
                        (N190)? mem[3664] : 
                        (N192)? mem[3744] : 
                        (N194)? mem[3824] : 
                        (N196)? mem[3904] : 
                        (N198)? mem[3984] : 
                        (N200)? mem[4064] : 
                        (N202)? mem[4144] : 
                        (N204)? mem[4224] : 
                        (N206)? mem[4304] : 
                        (N208)? mem[4384] : 
                        (N210)? mem[4464] : 
                        (N212)? mem[4544] : 
                        (N214)? mem[4624] : 
                        (N216)? mem[4704] : 
                        (N218)? mem[4784] : 
                        (N220)? mem[4864] : 
                        (N222)? mem[4944] : 
                        (N224)? mem[5024] : 
                        (N226)? mem[5104] : 1'b0;
  assign data_out[63] = (N163)? mem[63] : 
                        (N165)? mem[143] : 
                        (N167)? mem[223] : 
                        (N169)? mem[303] : 
                        (N171)? mem[383] : 
                        (N173)? mem[463] : 
                        (N175)? mem[543] : 
                        (N177)? mem[623] : 
                        (N179)? mem[703] : 
                        (N181)? mem[783] : 
                        (N183)? mem[863] : 
                        (N185)? mem[943] : 
                        (N187)? mem[1023] : 
                        (N189)? mem[1103] : 
                        (N191)? mem[1183] : 
                        (N193)? mem[1263] : 
                        (N195)? mem[1343] : 
                        (N197)? mem[1423] : 
                        (N199)? mem[1503] : 
                        (N201)? mem[1583] : 
                        (N203)? mem[1663] : 
                        (N205)? mem[1743] : 
                        (N207)? mem[1823] : 
                        (N209)? mem[1903] : 
                        (N211)? mem[1983] : 
                        (N213)? mem[2063] : 
                        (N215)? mem[2143] : 
                        (N217)? mem[2223] : 
                        (N219)? mem[2303] : 
                        (N221)? mem[2383] : 
                        (N223)? mem[2463] : 
                        (N225)? mem[2543] : 
                        (N164)? mem[2623] : 
                        (N166)? mem[2703] : 
                        (N168)? mem[2783] : 
                        (N170)? mem[2863] : 
                        (N172)? mem[2943] : 
                        (N174)? mem[3023] : 
                        (N176)? mem[3103] : 
                        (N178)? mem[3183] : 
                        (N180)? mem[3263] : 
                        (N182)? mem[3343] : 
                        (N184)? mem[3423] : 
                        (N186)? mem[3503] : 
                        (N188)? mem[3583] : 
                        (N190)? mem[3663] : 
                        (N192)? mem[3743] : 
                        (N194)? mem[3823] : 
                        (N196)? mem[3903] : 
                        (N198)? mem[3983] : 
                        (N200)? mem[4063] : 
                        (N202)? mem[4143] : 
                        (N204)? mem[4223] : 
                        (N206)? mem[4303] : 
                        (N208)? mem[4383] : 
                        (N210)? mem[4463] : 
                        (N212)? mem[4543] : 
                        (N214)? mem[4623] : 
                        (N216)? mem[4703] : 
                        (N218)? mem[4783] : 
                        (N220)? mem[4863] : 
                        (N222)? mem[4943] : 
                        (N224)? mem[5023] : 
                        (N226)? mem[5103] : 1'b0;
  assign data_out[62] = (N163)? mem[62] : 
                        (N165)? mem[142] : 
                        (N167)? mem[222] : 
                        (N169)? mem[302] : 
                        (N171)? mem[382] : 
                        (N173)? mem[462] : 
                        (N175)? mem[542] : 
                        (N177)? mem[622] : 
                        (N179)? mem[702] : 
                        (N181)? mem[782] : 
                        (N183)? mem[862] : 
                        (N185)? mem[942] : 
                        (N187)? mem[1022] : 
                        (N189)? mem[1102] : 
                        (N191)? mem[1182] : 
                        (N193)? mem[1262] : 
                        (N195)? mem[1342] : 
                        (N197)? mem[1422] : 
                        (N199)? mem[1502] : 
                        (N201)? mem[1582] : 
                        (N203)? mem[1662] : 
                        (N205)? mem[1742] : 
                        (N207)? mem[1822] : 
                        (N209)? mem[1902] : 
                        (N211)? mem[1982] : 
                        (N213)? mem[2062] : 
                        (N215)? mem[2142] : 
                        (N217)? mem[2222] : 
                        (N219)? mem[2302] : 
                        (N221)? mem[2382] : 
                        (N223)? mem[2462] : 
                        (N225)? mem[2542] : 
                        (N164)? mem[2622] : 
                        (N166)? mem[2702] : 
                        (N168)? mem[2782] : 
                        (N170)? mem[2862] : 
                        (N172)? mem[2942] : 
                        (N174)? mem[3022] : 
                        (N176)? mem[3102] : 
                        (N178)? mem[3182] : 
                        (N180)? mem[3262] : 
                        (N182)? mem[3342] : 
                        (N184)? mem[3422] : 
                        (N186)? mem[3502] : 
                        (N188)? mem[3582] : 
                        (N190)? mem[3662] : 
                        (N192)? mem[3742] : 
                        (N194)? mem[3822] : 
                        (N196)? mem[3902] : 
                        (N198)? mem[3982] : 
                        (N200)? mem[4062] : 
                        (N202)? mem[4142] : 
                        (N204)? mem[4222] : 
                        (N206)? mem[4302] : 
                        (N208)? mem[4382] : 
                        (N210)? mem[4462] : 
                        (N212)? mem[4542] : 
                        (N214)? mem[4622] : 
                        (N216)? mem[4702] : 
                        (N218)? mem[4782] : 
                        (N220)? mem[4862] : 
                        (N222)? mem[4942] : 
                        (N224)? mem[5022] : 
                        (N226)? mem[5102] : 1'b0;
  assign data_out[61] = (N163)? mem[61] : 
                        (N165)? mem[141] : 
                        (N167)? mem[221] : 
                        (N169)? mem[301] : 
                        (N171)? mem[381] : 
                        (N173)? mem[461] : 
                        (N175)? mem[541] : 
                        (N177)? mem[621] : 
                        (N179)? mem[701] : 
                        (N181)? mem[781] : 
                        (N183)? mem[861] : 
                        (N185)? mem[941] : 
                        (N187)? mem[1021] : 
                        (N189)? mem[1101] : 
                        (N191)? mem[1181] : 
                        (N193)? mem[1261] : 
                        (N195)? mem[1341] : 
                        (N197)? mem[1421] : 
                        (N199)? mem[1501] : 
                        (N201)? mem[1581] : 
                        (N203)? mem[1661] : 
                        (N205)? mem[1741] : 
                        (N207)? mem[1821] : 
                        (N209)? mem[1901] : 
                        (N211)? mem[1981] : 
                        (N213)? mem[2061] : 
                        (N215)? mem[2141] : 
                        (N217)? mem[2221] : 
                        (N219)? mem[2301] : 
                        (N221)? mem[2381] : 
                        (N223)? mem[2461] : 
                        (N225)? mem[2541] : 
                        (N164)? mem[2621] : 
                        (N166)? mem[2701] : 
                        (N168)? mem[2781] : 
                        (N170)? mem[2861] : 
                        (N172)? mem[2941] : 
                        (N174)? mem[3021] : 
                        (N176)? mem[3101] : 
                        (N178)? mem[3181] : 
                        (N180)? mem[3261] : 
                        (N182)? mem[3341] : 
                        (N184)? mem[3421] : 
                        (N186)? mem[3501] : 
                        (N188)? mem[3581] : 
                        (N190)? mem[3661] : 
                        (N192)? mem[3741] : 
                        (N194)? mem[3821] : 
                        (N196)? mem[3901] : 
                        (N198)? mem[3981] : 
                        (N200)? mem[4061] : 
                        (N202)? mem[4141] : 
                        (N204)? mem[4221] : 
                        (N206)? mem[4301] : 
                        (N208)? mem[4381] : 
                        (N210)? mem[4461] : 
                        (N212)? mem[4541] : 
                        (N214)? mem[4621] : 
                        (N216)? mem[4701] : 
                        (N218)? mem[4781] : 
                        (N220)? mem[4861] : 
                        (N222)? mem[4941] : 
                        (N224)? mem[5021] : 
                        (N226)? mem[5101] : 1'b0;
  assign data_out[60] = (N163)? mem[60] : 
                        (N165)? mem[140] : 
                        (N167)? mem[220] : 
                        (N169)? mem[300] : 
                        (N171)? mem[380] : 
                        (N173)? mem[460] : 
                        (N175)? mem[540] : 
                        (N177)? mem[620] : 
                        (N179)? mem[700] : 
                        (N181)? mem[780] : 
                        (N183)? mem[860] : 
                        (N185)? mem[940] : 
                        (N187)? mem[1020] : 
                        (N189)? mem[1100] : 
                        (N191)? mem[1180] : 
                        (N193)? mem[1260] : 
                        (N195)? mem[1340] : 
                        (N197)? mem[1420] : 
                        (N199)? mem[1500] : 
                        (N201)? mem[1580] : 
                        (N203)? mem[1660] : 
                        (N205)? mem[1740] : 
                        (N207)? mem[1820] : 
                        (N209)? mem[1900] : 
                        (N211)? mem[1980] : 
                        (N213)? mem[2060] : 
                        (N215)? mem[2140] : 
                        (N217)? mem[2220] : 
                        (N219)? mem[2300] : 
                        (N221)? mem[2380] : 
                        (N223)? mem[2460] : 
                        (N225)? mem[2540] : 
                        (N164)? mem[2620] : 
                        (N166)? mem[2700] : 
                        (N168)? mem[2780] : 
                        (N170)? mem[2860] : 
                        (N172)? mem[2940] : 
                        (N174)? mem[3020] : 
                        (N176)? mem[3100] : 
                        (N178)? mem[3180] : 
                        (N180)? mem[3260] : 
                        (N182)? mem[3340] : 
                        (N184)? mem[3420] : 
                        (N186)? mem[3500] : 
                        (N188)? mem[3580] : 
                        (N190)? mem[3660] : 
                        (N192)? mem[3740] : 
                        (N194)? mem[3820] : 
                        (N196)? mem[3900] : 
                        (N198)? mem[3980] : 
                        (N200)? mem[4060] : 
                        (N202)? mem[4140] : 
                        (N204)? mem[4220] : 
                        (N206)? mem[4300] : 
                        (N208)? mem[4380] : 
                        (N210)? mem[4460] : 
                        (N212)? mem[4540] : 
                        (N214)? mem[4620] : 
                        (N216)? mem[4700] : 
                        (N218)? mem[4780] : 
                        (N220)? mem[4860] : 
                        (N222)? mem[4940] : 
                        (N224)? mem[5020] : 
                        (N226)? mem[5100] : 1'b0;
  assign data_out[59] = (N163)? mem[59] : 
                        (N165)? mem[139] : 
                        (N167)? mem[219] : 
                        (N169)? mem[299] : 
                        (N171)? mem[379] : 
                        (N173)? mem[459] : 
                        (N175)? mem[539] : 
                        (N177)? mem[619] : 
                        (N179)? mem[699] : 
                        (N181)? mem[779] : 
                        (N183)? mem[859] : 
                        (N185)? mem[939] : 
                        (N187)? mem[1019] : 
                        (N189)? mem[1099] : 
                        (N191)? mem[1179] : 
                        (N193)? mem[1259] : 
                        (N195)? mem[1339] : 
                        (N197)? mem[1419] : 
                        (N199)? mem[1499] : 
                        (N201)? mem[1579] : 
                        (N203)? mem[1659] : 
                        (N205)? mem[1739] : 
                        (N207)? mem[1819] : 
                        (N209)? mem[1899] : 
                        (N211)? mem[1979] : 
                        (N213)? mem[2059] : 
                        (N215)? mem[2139] : 
                        (N217)? mem[2219] : 
                        (N219)? mem[2299] : 
                        (N221)? mem[2379] : 
                        (N223)? mem[2459] : 
                        (N225)? mem[2539] : 
                        (N164)? mem[2619] : 
                        (N166)? mem[2699] : 
                        (N168)? mem[2779] : 
                        (N170)? mem[2859] : 
                        (N172)? mem[2939] : 
                        (N174)? mem[3019] : 
                        (N176)? mem[3099] : 
                        (N178)? mem[3179] : 
                        (N180)? mem[3259] : 
                        (N182)? mem[3339] : 
                        (N184)? mem[3419] : 
                        (N186)? mem[3499] : 
                        (N188)? mem[3579] : 
                        (N190)? mem[3659] : 
                        (N192)? mem[3739] : 
                        (N194)? mem[3819] : 
                        (N196)? mem[3899] : 
                        (N198)? mem[3979] : 
                        (N200)? mem[4059] : 
                        (N202)? mem[4139] : 
                        (N204)? mem[4219] : 
                        (N206)? mem[4299] : 
                        (N208)? mem[4379] : 
                        (N210)? mem[4459] : 
                        (N212)? mem[4539] : 
                        (N214)? mem[4619] : 
                        (N216)? mem[4699] : 
                        (N218)? mem[4779] : 
                        (N220)? mem[4859] : 
                        (N222)? mem[4939] : 
                        (N224)? mem[5019] : 
                        (N226)? mem[5099] : 1'b0;
  assign data_out[58] = (N163)? mem[58] : 
                        (N165)? mem[138] : 
                        (N167)? mem[218] : 
                        (N169)? mem[298] : 
                        (N171)? mem[378] : 
                        (N173)? mem[458] : 
                        (N175)? mem[538] : 
                        (N177)? mem[618] : 
                        (N179)? mem[698] : 
                        (N181)? mem[778] : 
                        (N183)? mem[858] : 
                        (N185)? mem[938] : 
                        (N187)? mem[1018] : 
                        (N189)? mem[1098] : 
                        (N191)? mem[1178] : 
                        (N193)? mem[1258] : 
                        (N195)? mem[1338] : 
                        (N197)? mem[1418] : 
                        (N199)? mem[1498] : 
                        (N201)? mem[1578] : 
                        (N203)? mem[1658] : 
                        (N205)? mem[1738] : 
                        (N207)? mem[1818] : 
                        (N209)? mem[1898] : 
                        (N211)? mem[1978] : 
                        (N213)? mem[2058] : 
                        (N215)? mem[2138] : 
                        (N217)? mem[2218] : 
                        (N219)? mem[2298] : 
                        (N221)? mem[2378] : 
                        (N223)? mem[2458] : 
                        (N225)? mem[2538] : 
                        (N164)? mem[2618] : 
                        (N166)? mem[2698] : 
                        (N168)? mem[2778] : 
                        (N170)? mem[2858] : 
                        (N172)? mem[2938] : 
                        (N174)? mem[3018] : 
                        (N176)? mem[3098] : 
                        (N178)? mem[3178] : 
                        (N180)? mem[3258] : 
                        (N182)? mem[3338] : 
                        (N184)? mem[3418] : 
                        (N186)? mem[3498] : 
                        (N188)? mem[3578] : 
                        (N190)? mem[3658] : 
                        (N192)? mem[3738] : 
                        (N194)? mem[3818] : 
                        (N196)? mem[3898] : 
                        (N198)? mem[3978] : 
                        (N200)? mem[4058] : 
                        (N202)? mem[4138] : 
                        (N204)? mem[4218] : 
                        (N206)? mem[4298] : 
                        (N208)? mem[4378] : 
                        (N210)? mem[4458] : 
                        (N212)? mem[4538] : 
                        (N214)? mem[4618] : 
                        (N216)? mem[4698] : 
                        (N218)? mem[4778] : 
                        (N220)? mem[4858] : 
                        (N222)? mem[4938] : 
                        (N224)? mem[5018] : 
                        (N226)? mem[5098] : 1'b0;
  assign data_out[57] = (N163)? mem[57] : 
                        (N165)? mem[137] : 
                        (N167)? mem[217] : 
                        (N169)? mem[297] : 
                        (N171)? mem[377] : 
                        (N173)? mem[457] : 
                        (N175)? mem[537] : 
                        (N177)? mem[617] : 
                        (N179)? mem[697] : 
                        (N181)? mem[777] : 
                        (N183)? mem[857] : 
                        (N185)? mem[937] : 
                        (N187)? mem[1017] : 
                        (N189)? mem[1097] : 
                        (N191)? mem[1177] : 
                        (N193)? mem[1257] : 
                        (N195)? mem[1337] : 
                        (N197)? mem[1417] : 
                        (N199)? mem[1497] : 
                        (N201)? mem[1577] : 
                        (N203)? mem[1657] : 
                        (N205)? mem[1737] : 
                        (N207)? mem[1817] : 
                        (N209)? mem[1897] : 
                        (N211)? mem[1977] : 
                        (N213)? mem[2057] : 
                        (N215)? mem[2137] : 
                        (N217)? mem[2217] : 
                        (N219)? mem[2297] : 
                        (N221)? mem[2377] : 
                        (N223)? mem[2457] : 
                        (N225)? mem[2537] : 
                        (N164)? mem[2617] : 
                        (N166)? mem[2697] : 
                        (N168)? mem[2777] : 
                        (N170)? mem[2857] : 
                        (N172)? mem[2937] : 
                        (N174)? mem[3017] : 
                        (N176)? mem[3097] : 
                        (N178)? mem[3177] : 
                        (N180)? mem[3257] : 
                        (N182)? mem[3337] : 
                        (N184)? mem[3417] : 
                        (N186)? mem[3497] : 
                        (N188)? mem[3577] : 
                        (N190)? mem[3657] : 
                        (N192)? mem[3737] : 
                        (N194)? mem[3817] : 
                        (N196)? mem[3897] : 
                        (N198)? mem[3977] : 
                        (N200)? mem[4057] : 
                        (N202)? mem[4137] : 
                        (N204)? mem[4217] : 
                        (N206)? mem[4297] : 
                        (N208)? mem[4377] : 
                        (N210)? mem[4457] : 
                        (N212)? mem[4537] : 
                        (N214)? mem[4617] : 
                        (N216)? mem[4697] : 
                        (N218)? mem[4777] : 
                        (N220)? mem[4857] : 
                        (N222)? mem[4937] : 
                        (N224)? mem[5017] : 
                        (N226)? mem[5097] : 1'b0;
  assign data_out[56] = (N163)? mem[56] : 
                        (N165)? mem[136] : 
                        (N167)? mem[216] : 
                        (N169)? mem[296] : 
                        (N171)? mem[376] : 
                        (N173)? mem[456] : 
                        (N175)? mem[536] : 
                        (N177)? mem[616] : 
                        (N179)? mem[696] : 
                        (N181)? mem[776] : 
                        (N183)? mem[856] : 
                        (N185)? mem[936] : 
                        (N187)? mem[1016] : 
                        (N189)? mem[1096] : 
                        (N191)? mem[1176] : 
                        (N193)? mem[1256] : 
                        (N195)? mem[1336] : 
                        (N197)? mem[1416] : 
                        (N199)? mem[1496] : 
                        (N201)? mem[1576] : 
                        (N203)? mem[1656] : 
                        (N205)? mem[1736] : 
                        (N207)? mem[1816] : 
                        (N209)? mem[1896] : 
                        (N211)? mem[1976] : 
                        (N213)? mem[2056] : 
                        (N215)? mem[2136] : 
                        (N217)? mem[2216] : 
                        (N219)? mem[2296] : 
                        (N221)? mem[2376] : 
                        (N223)? mem[2456] : 
                        (N225)? mem[2536] : 
                        (N164)? mem[2616] : 
                        (N166)? mem[2696] : 
                        (N168)? mem[2776] : 
                        (N170)? mem[2856] : 
                        (N172)? mem[2936] : 
                        (N174)? mem[3016] : 
                        (N176)? mem[3096] : 
                        (N178)? mem[3176] : 
                        (N180)? mem[3256] : 
                        (N182)? mem[3336] : 
                        (N184)? mem[3416] : 
                        (N186)? mem[3496] : 
                        (N188)? mem[3576] : 
                        (N190)? mem[3656] : 
                        (N192)? mem[3736] : 
                        (N194)? mem[3816] : 
                        (N196)? mem[3896] : 
                        (N198)? mem[3976] : 
                        (N200)? mem[4056] : 
                        (N202)? mem[4136] : 
                        (N204)? mem[4216] : 
                        (N206)? mem[4296] : 
                        (N208)? mem[4376] : 
                        (N210)? mem[4456] : 
                        (N212)? mem[4536] : 
                        (N214)? mem[4616] : 
                        (N216)? mem[4696] : 
                        (N218)? mem[4776] : 
                        (N220)? mem[4856] : 
                        (N222)? mem[4936] : 
                        (N224)? mem[5016] : 
                        (N226)? mem[5096] : 1'b0;
  assign data_out[55] = (N163)? mem[55] : 
                        (N165)? mem[135] : 
                        (N167)? mem[215] : 
                        (N169)? mem[295] : 
                        (N171)? mem[375] : 
                        (N173)? mem[455] : 
                        (N175)? mem[535] : 
                        (N177)? mem[615] : 
                        (N179)? mem[695] : 
                        (N181)? mem[775] : 
                        (N183)? mem[855] : 
                        (N185)? mem[935] : 
                        (N187)? mem[1015] : 
                        (N189)? mem[1095] : 
                        (N191)? mem[1175] : 
                        (N193)? mem[1255] : 
                        (N195)? mem[1335] : 
                        (N197)? mem[1415] : 
                        (N199)? mem[1495] : 
                        (N201)? mem[1575] : 
                        (N203)? mem[1655] : 
                        (N205)? mem[1735] : 
                        (N207)? mem[1815] : 
                        (N209)? mem[1895] : 
                        (N211)? mem[1975] : 
                        (N213)? mem[2055] : 
                        (N215)? mem[2135] : 
                        (N217)? mem[2215] : 
                        (N219)? mem[2295] : 
                        (N221)? mem[2375] : 
                        (N223)? mem[2455] : 
                        (N225)? mem[2535] : 
                        (N164)? mem[2615] : 
                        (N166)? mem[2695] : 
                        (N168)? mem[2775] : 
                        (N170)? mem[2855] : 
                        (N172)? mem[2935] : 
                        (N174)? mem[3015] : 
                        (N176)? mem[3095] : 
                        (N178)? mem[3175] : 
                        (N180)? mem[3255] : 
                        (N182)? mem[3335] : 
                        (N184)? mem[3415] : 
                        (N186)? mem[3495] : 
                        (N188)? mem[3575] : 
                        (N190)? mem[3655] : 
                        (N192)? mem[3735] : 
                        (N194)? mem[3815] : 
                        (N196)? mem[3895] : 
                        (N198)? mem[3975] : 
                        (N200)? mem[4055] : 
                        (N202)? mem[4135] : 
                        (N204)? mem[4215] : 
                        (N206)? mem[4295] : 
                        (N208)? mem[4375] : 
                        (N210)? mem[4455] : 
                        (N212)? mem[4535] : 
                        (N214)? mem[4615] : 
                        (N216)? mem[4695] : 
                        (N218)? mem[4775] : 
                        (N220)? mem[4855] : 
                        (N222)? mem[4935] : 
                        (N224)? mem[5015] : 
                        (N226)? mem[5095] : 1'b0;
  assign data_out[54] = (N163)? mem[54] : 
                        (N165)? mem[134] : 
                        (N167)? mem[214] : 
                        (N169)? mem[294] : 
                        (N171)? mem[374] : 
                        (N173)? mem[454] : 
                        (N175)? mem[534] : 
                        (N177)? mem[614] : 
                        (N179)? mem[694] : 
                        (N181)? mem[774] : 
                        (N183)? mem[854] : 
                        (N185)? mem[934] : 
                        (N187)? mem[1014] : 
                        (N189)? mem[1094] : 
                        (N191)? mem[1174] : 
                        (N193)? mem[1254] : 
                        (N195)? mem[1334] : 
                        (N197)? mem[1414] : 
                        (N199)? mem[1494] : 
                        (N201)? mem[1574] : 
                        (N203)? mem[1654] : 
                        (N205)? mem[1734] : 
                        (N207)? mem[1814] : 
                        (N209)? mem[1894] : 
                        (N211)? mem[1974] : 
                        (N213)? mem[2054] : 
                        (N215)? mem[2134] : 
                        (N217)? mem[2214] : 
                        (N219)? mem[2294] : 
                        (N221)? mem[2374] : 
                        (N223)? mem[2454] : 
                        (N225)? mem[2534] : 
                        (N164)? mem[2614] : 
                        (N166)? mem[2694] : 
                        (N168)? mem[2774] : 
                        (N170)? mem[2854] : 
                        (N172)? mem[2934] : 
                        (N174)? mem[3014] : 
                        (N176)? mem[3094] : 
                        (N178)? mem[3174] : 
                        (N180)? mem[3254] : 
                        (N182)? mem[3334] : 
                        (N184)? mem[3414] : 
                        (N186)? mem[3494] : 
                        (N188)? mem[3574] : 
                        (N190)? mem[3654] : 
                        (N192)? mem[3734] : 
                        (N194)? mem[3814] : 
                        (N196)? mem[3894] : 
                        (N198)? mem[3974] : 
                        (N200)? mem[4054] : 
                        (N202)? mem[4134] : 
                        (N204)? mem[4214] : 
                        (N206)? mem[4294] : 
                        (N208)? mem[4374] : 
                        (N210)? mem[4454] : 
                        (N212)? mem[4534] : 
                        (N214)? mem[4614] : 
                        (N216)? mem[4694] : 
                        (N218)? mem[4774] : 
                        (N220)? mem[4854] : 
                        (N222)? mem[4934] : 
                        (N224)? mem[5014] : 
                        (N226)? mem[5094] : 1'b0;
  assign data_out[53] = (N163)? mem[53] : 
                        (N165)? mem[133] : 
                        (N167)? mem[213] : 
                        (N169)? mem[293] : 
                        (N171)? mem[373] : 
                        (N173)? mem[453] : 
                        (N175)? mem[533] : 
                        (N177)? mem[613] : 
                        (N179)? mem[693] : 
                        (N181)? mem[773] : 
                        (N183)? mem[853] : 
                        (N185)? mem[933] : 
                        (N187)? mem[1013] : 
                        (N189)? mem[1093] : 
                        (N191)? mem[1173] : 
                        (N193)? mem[1253] : 
                        (N195)? mem[1333] : 
                        (N197)? mem[1413] : 
                        (N199)? mem[1493] : 
                        (N201)? mem[1573] : 
                        (N203)? mem[1653] : 
                        (N205)? mem[1733] : 
                        (N207)? mem[1813] : 
                        (N209)? mem[1893] : 
                        (N211)? mem[1973] : 
                        (N213)? mem[2053] : 
                        (N215)? mem[2133] : 
                        (N217)? mem[2213] : 
                        (N219)? mem[2293] : 
                        (N221)? mem[2373] : 
                        (N223)? mem[2453] : 
                        (N225)? mem[2533] : 
                        (N164)? mem[2613] : 
                        (N166)? mem[2693] : 
                        (N168)? mem[2773] : 
                        (N170)? mem[2853] : 
                        (N172)? mem[2933] : 
                        (N174)? mem[3013] : 
                        (N176)? mem[3093] : 
                        (N178)? mem[3173] : 
                        (N180)? mem[3253] : 
                        (N182)? mem[3333] : 
                        (N184)? mem[3413] : 
                        (N186)? mem[3493] : 
                        (N188)? mem[3573] : 
                        (N190)? mem[3653] : 
                        (N192)? mem[3733] : 
                        (N194)? mem[3813] : 
                        (N196)? mem[3893] : 
                        (N198)? mem[3973] : 
                        (N200)? mem[4053] : 
                        (N202)? mem[4133] : 
                        (N204)? mem[4213] : 
                        (N206)? mem[4293] : 
                        (N208)? mem[4373] : 
                        (N210)? mem[4453] : 
                        (N212)? mem[4533] : 
                        (N214)? mem[4613] : 
                        (N216)? mem[4693] : 
                        (N218)? mem[4773] : 
                        (N220)? mem[4853] : 
                        (N222)? mem[4933] : 
                        (N224)? mem[5013] : 
                        (N226)? mem[5093] : 1'b0;
  assign data_out[52] = (N163)? mem[52] : 
                        (N165)? mem[132] : 
                        (N167)? mem[212] : 
                        (N169)? mem[292] : 
                        (N171)? mem[372] : 
                        (N173)? mem[452] : 
                        (N175)? mem[532] : 
                        (N177)? mem[612] : 
                        (N179)? mem[692] : 
                        (N181)? mem[772] : 
                        (N183)? mem[852] : 
                        (N185)? mem[932] : 
                        (N187)? mem[1012] : 
                        (N189)? mem[1092] : 
                        (N191)? mem[1172] : 
                        (N193)? mem[1252] : 
                        (N195)? mem[1332] : 
                        (N197)? mem[1412] : 
                        (N199)? mem[1492] : 
                        (N201)? mem[1572] : 
                        (N203)? mem[1652] : 
                        (N205)? mem[1732] : 
                        (N207)? mem[1812] : 
                        (N209)? mem[1892] : 
                        (N211)? mem[1972] : 
                        (N213)? mem[2052] : 
                        (N215)? mem[2132] : 
                        (N217)? mem[2212] : 
                        (N219)? mem[2292] : 
                        (N221)? mem[2372] : 
                        (N223)? mem[2452] : 
                        (N225)? mem[2532] : 
                        (N164)? mem[2612] : 
                        (N166)? mem[2692] : 
                        (N168)? mem[2772] : 
                        (N170)? mem[2852] : 
                        (N172)? mem[2932] : 
                        (N174)? mem[3012] : 
                        (N176)? mem[3092] : 
                        (N178)? mem[3172] : 
                        (N180)? mem[3252] : 
                        (N182)? mem[3332] : 
                        (N184)? mem[3412] : 
                        (N186)? mem[3492] : 
                        (N188)? mem[3572] : 
                        (N190)? mem[3652] : 
                        (N192)? mem[3732] : 
                        (N194)? mem[3812] : 
                        (N196)? mem[3892] : 
                        (N198)? mem[3972] : 
                        (N200)? mem[4052] : 
                        (N202)? mem[4132] : 
                        (N204)? mem[4212] : 
                        (N206)? mem[4292] : 
                        (N208)? mem[4372] : 
                        (N210)? mem[4452] : 
                        (N212)? mem[4532] : 
                        (N214)? mem[4612] : 
                        (N216)? mem[4692] : 
                        (N218)? mem[4772] : 
                        (N220)? mem[4852] : 
                        (N222)? mem[4932] : 
                        (N224)? mem[5012] : 
                        (N226)? mem[5092] : 1'b0;
  assign data_out[51] = (N163)? mem[51] : 
                        (N165)? mem[131] : 
                        (N167)? mem[211] : 
                        (N169)? mem[291] : 
                        (N171)? mem[371] : 
                        (N173)? mem[451] : 
                        (N175)? mem[531] : 
                        (N177)? mem[611] : 
                        (N179)? mem[691] : 
                        (N181)? mem[771] : 
                        (N183)? mem[851] : 
                        (N185)? mem[931] : 
                        (N187)? mem[1011] : 
                        (N189)? mem[1091] : 
                        (N191)? mem[1171] : 
                        (N193)? mem[1251] : 
                        (N195)? mem[1331] : 
                        (N197)? mem[1411] : 
                        (N199)? mem[1491] : 
                        (N201)? mem[1571] : 
                        (N203)? mem[1651] : 
                        (N205)? mem[1731] : 
                        (N207)? mem[1811] : 
                        (N209)? mem[1891] : 
                        (N211)? mem[1971] : 
                        (N213)? mem[2051] : 
                        (N215)? mem[2131] : 
                        (N217)? mem[2211] : 
                        (N219)? mem[2291] : 
                        (N221)? mem[2371] : 
                        (N223)? mem[2451] : 
                        (N225)? mem[2531] : 
                        (N164)? mem[2611] : 
                        (N166)? mem[2691] : 
                        (N168)? mem[2771] : 
                        (N170)? mem[2851] : 
                        (N172)? mem[2931] : 
                        (N174)? mem[3011] : 
                        (N176)? mem[3091] : 
                        (N178)? mem[3171] : 
                        (N180)? mem[3251] : 
                        (N182)? mem[3331] : 
                        (N184)? mem[3411] : 
                        (N186)? mem[3491] : 
                        (N188)? mem[3571] : 
                        (N190)? mem[3651] : 
                        (N192)? mem[3731] : 
                        (N194)? mem[3811] : 
                        (N196)? mem[3891] : 
                        (N198)? mem[3971] : 
                        (N200)? mem[4051] : 
                        (N202)? mem[4131] : 
                        (N204)? mem[4211] : 
                        (N206)? mem[4291] : 
                        (N208)? mem[4371] : 
                        (N210)? mem[4451] : 
                        (N212)? mem[4531] : 
                        (N214)? mem[4611] : 
                        (N216)? mem[4691] : 
                        (N218)? mem[4771] : 
                        (N220)? mem[4851] : 
                        (N222)? mem[4931] : 
                        (N224)? mem[5011] : 
                        (N226)? mem[5091] : 1'b0;
  assign data_out[50] = (N163)? mem[50] : 
                        (N165)? mem[130] : 
                        (N167)? mem[210] : 
                        (N169)? mem[290] : 
                        (N171)? mem[370] : 
                        (N173)? mem[450] : 
                        (N175)? mem[530] : 
                        (N177)? mem[610] : 
                        (N179)? mem[690] : 
                        (N181)? mem[770] : 
                        (N183)? mem[850] : 
                        (N185)? mem[930] : 
                        (N187)? mem[1010] : 
                        (N189)? mem[1090] : 
                        (N191)? mem[1170] : 
                        (N193)? mem[1250] : 
                        (N195)? mem[1330] : 
                        (N197)? mem[1410] : 
                        (N199)? mem[1490] : 
                        (N201)? mem[1570] : 
                        (N203)? mem[1650] : 
                        (N205)? mem[1730] : 
                        (N207)? mem[1810] : 
                        (N209)? mem[1890] : 
                        (N211)? mem[1970] : 
                        (N213)? mem[2050] : 
                        (N215)? mem[2130] : 
                        (N217)? mem[2210] : 
                        (N219)? mem[2290] : 
                        (N221)? mem[2370] : 
                        (N223)? mem[2450] : 
                        (N225)? mem[2530] : 
                        (N164)? mem[2610] : 
                        (N166)? mem[2690] : 
                        (N168)? mem[2770] : 
                        (N170)? mem[2850] : 
                        (N172)? mem[2930] : 
                        (N174)? mem[3010] : 
                        (N176)? mem[3090] : 
                        (N178)? mem[3170] : 
                        (N180)? mem[3250] : 
                        (N182)? mem[3330] : 
                        (N184)? mem[3410] : 
                        (N186)? mem[3490] : 
                        (N188)? mem[3570] : 
                        (N190)? mem[3650] : 
                        (N192)? mem[3730] : 
                        (N194)? mem[3810] : 
                        (N196)? mem[3890] : 
                        (N198)? mem[3970] : 
                        (N200)? mem[4050] : 
                        (N202)? mem[4130] : 
                        (N204)? mem[4210] : 
                        (N206)? mem[4290] : 
                        (N208)? mem[4370] : 
                        (N210)? mem[4450] : 
                        (N212)? mem[4530] : 
                        (N214)? mem[4610] : 
                        (N216)? mem[4690] : 
                        (N218)? mem[4770] : 
                        (N220)? mem[4850] : 
                        (N222)? mem[4930] : 
                        (N224)? mem[5010] : 
                        (N226)? mem[5090] : 1'b0;
  assign data_out[49] = (N163)? mem[49] : 
                        (N165)? mem[129] : 
                        (N167)? mem[209] : 
                        (N169)? mem[289] : 
                        (N171)? mem[369] : 
                        (N173)? mem[449] : 
                        (N175)? mem[529] : 
                        (N177)? mem[609] : 
                        (N179)? mem[689] : 
                        (N181)? mem[769] : 
                        (N183)? mem[849] : 
                        (N185)? mem[929] : 
                        (N187)? mem[1009] : 
                        (N189)? mem[1089] : 
                        (N191)? mem[1169] : 
                        (N193)? mem[1249] : 
                        (N195)? mem[1329] : 
                        (N197)? mem[1409] : 
                        (N199)? mem[1489] : 
                        (N201)? mem[1569] : 
                        (N203)? mem[1649] : 
                        (N205)? mem[1729] : 
                        (N207)? mem[1809] : 
                        (N209)? mem[1889] : 
                        (N211)? mem[1969] : 
                        (N213)? mem[2049] : 
                        (N215)? mem[2129] : 
                        (N217)? mem[2209] : 
                        (N219)? mem[2289] : 
                        (N221)? mem[2369] : 
                        (N223)? mem[2449] : 
                        (N225)? mem[2529] : 
                        (N164)? mem[2609] : 
                        (N166)? mem[2689] : 
                        (N168)? mem[2769] : 
                        (N170)? mem[2849] : 
                        (N172)? mem[2929] : 
                        (N174)? mem[3009] : 
                        (N176)? mem[3089] : 
                        (N178)? mem[3169] : 
                        (N180)? mem[3249] : 
                        (N182)? mem[3329] : 
                        (N184)? mem[3409] : 
                        (N186)? mem[3489] : 
                        (N188)? mem[3569] : 
                        (N190)? mem[3649] : 
                        (N192)? mem[3729] : 
                        (N194)? mem[3809] : 
                        (N196)? mem[3889] : 
                        (N198)? mem[3969] : 
                        (N200)? mem[4049] : 
                        (N202)? mem[4129] : 
                        (N204)? mem[4209] : 
                        (N206)? mem[4289] : 
                        (N208)? mem[4369] : 
                        (N210)? mem[4449] : 
                        (N212)? mem[4529] : 
                        (N214)? mem[4609] : 
                        (N216)? mem[4689] : 
                        (N218)? mem[4769] : 
                        (N220)? mem[4849] : 
                        (N222)? mem[4929] : 
                        (N224)? mem[5009] : 
                        (N226)? mem[5089] : 1'b0;
  assign data_out[48] = (N163)? mem[48] : 
                        (N165)? mem[128] : 
                        (N167)? mem[208] : 
                        (N169)? mem[288] : 
                        (N171)? mem[368] : 
                        (N173)? mem[448] : 
                        (N175)? mem[528] : 
                        (N177)? mem[608] : 
                        (N179)? mem[688] : 
                        (N181)? mem[768] : 
                        (N183)? mem[848] : 
                        (N185)? mem[928] : 
                        (N187)? mem[1008] : 
                        (N189)? mem[1088] : 
                        (N191)? mem[1168] : 
                        (N193)? mem[1248] : 
                        (N195)? mem[1328] : 
                        (N197)? mem[1408] : 
                        (N199)? mem[1488] : 
                        (N201)? mem[1568] : 
                        (N203)? mem[1648] : 
                        (N205)? mem[1728] : 
                        (N207)? mem[1808] : 
                        (N209)? mem[1888] : 
                        (N211)? mem[1968] : 
                        (N213)? mem[2048] : 
                        (N215)? mem[2128] : 
                        (N217)? mem[2208] : 
                        (N219)? mem[2288] : 
                        (N221)? mem[2368] : 
                        (N223)? mem[2448] : 
                        (N225)? mem[2528] : 
                        (N164)? mem[2608] : 
                        (N166)? mem[2688] : 
                        (N168)? mem[2768] : 
                        (N170)? mem[2848] : 
                        (N172)? mem[2928] : 
                        (N174)? mem[3008] : 
                        (N176)? mem[3088] : 
                        (N178)? mem[3168] : 
                        (N180)? mem[3248] : 
                        (N182)? mem[3328] : 
                        (N184)? mem[3408] : 
                        (N186)? mem[3488] : 
                        (N188)? mem[3568] : 
                        (N190)? mem[3648] : 
                        (N192)? mem[3728] : 
                        (N194)? mem[3808] : 
                        (N196)? mem[3888] : 
                        (N198)? mem[3968] : 
                        (N200)? mem[4048] : 
                        (N202)? mem[4128] : 
                        (N204)? mem[4208] : 
                        (N206)? mem[4288] : 
                        (N208)? mem[4368] : 
                        (N210)? mem[4448] : 
                        (N212)? mem[4528] : 
                        (N214)? mem[4608] : 
                        (N216)? mem[4688] : 
                        (N218)? mem[4768] : 
                        (N220)? mem[4848] : 
                        (N222)? mem[4928] : 
                        (N224)? mem[5008] : 
                        (N226)? mem[5088] : 1'b0;
  assign data_out[47] = (N163)? mem[47] : 
                        (N165)? mem[127] : 
                        (N167)? mem[207] : 
                        (N169)? mem[287] : 
                        (N171)? mem[367] : 
                        (N173)? mem[447] : 
                        (N175)? mem[527] : 
                        (N177)? mem[607] : 
                        (N179)? mem[687] : 
                        (N181)? mem[767] : 
                        (N183)? mem[847] : 
                        (N185)? mem[927] : 
                        (N187)? mem[1007] : 
                        (N189)? mem[1087] : 
                        (N191)? mem[1167] : 
                        (N193)? mem[1247] : 
                        (N195)? mem[1327] : 
                        (N197)? mem[1407] : 
                        (N199)? mem[1487] : 
                        (N201)? mem[1567] : 
                        (N203)? mem[1647] : 
                        (N205)? mem[1727] : 
                        (N207)? mem[1807] : 
                        (N209)? mem[1887] : 
                        (N211)? mem[1967] : 
                        (N213)? mem[2047] : 
                        (N215)? mem[2127] : 
                        (N217)? mem[2207] : 
                        (N219)? mem[2287] : 
                        (N221)? mem[2367] : 
                        (N223)? mem[2447] : 
                        (N225)? mem[2527] : 
                        (N164)? mem[2607] : 
                        (N166)? mem[2687] : 
                        (N168)? mem[2767] : 
                        (N170)? mem[2847] : 
                        (N172)? mem[2927] : 
                        (N174)? mem[3007] : 
                        (N176)? mem[3087] : 
                        (N178)? mem[3167] : 
                        (N180)? mem[3247] : 
                        (N182)? mem[3327] : 
                        (N184)? mem[3407] : 
                        (N186)? mem[3487] : 
                        (N188)? mem[3567] : 
                        (N190)? mem[3647] : 
                        (N192)? mem[3727] : 
                        (N194)? mem[3807] : 
                        (N196)? mem[3887] : 
                        (N198)? mem[3967] : 
                        (N200)? mem[4047] : 
                        (N202)? mem[4127] : 
                        (N204)? mem[4207] : 
                        (N206)? mem[4287] : 
                        (N208)? mem[4367] : 
                        (N210)? mem[4447] : 
                        (N212)? mem[4527] : 
                        (N214)? mem[4607] : 
                        (N216)? mem[4687] : 
                        (N218)? mem[4767] : 
                        (N220)? mem[4847] : 
                        (N222)? mem[4927] : 
                        (N224)? mem[5007] : 
                        (N226)? mem[5087] : 1'b0;
  assign data_out[46] = (N163)? mem[46] : 
                        (N165)? mem[126] : 
                        (N167)? mem[206] : 
                        (N169)? mem[286] : 
                        (N171)? mem[366] : 
                        (N173)? mem[446] : 
                        (N175)? mem[526] : 
                        (N177)? mem[606] : 
                        (N179)? mem[686] : 
                        (N181)? mem[766] : 
                        (N183)? mem[846] : 
                        (N185)? mem[926] : 
                        (N187)? mem[1006] : 
                        (N189)? mem[1086] : 
                        (N191)? mem[1166] : 
                        (N193)? mem[1246] : 
                        (N195)? mem[1326] : 
                        (N197)? mem[1406] : 
                        (N199)? mem[1486] : 
                        (N201)? mem[1566] : 
                        (N203)? mem[1646] : 
                        (N205)? mem[1726] : 
                        (N207)? mem[1806] : 
                        (N209)? mem[1886] : 
                        (N211)? mem[1966] : 
                        (N213)? mem[2046] : 
                        (N215)? mem[2126] : 
                        (N217)? mem[2206] : 
                        (N219)? mem[2286] : 
                        (N221)? mem[2366] : 
                        (N223)? mem[2446] : 
                        (N225)? mem[2526] : 
                        (N164)? mem[2606] : 
                        (N166)? mem[2686] : 
                        (N168)? mem[2766] : 
                        (N170)? mem[2846] : 
                        (N172)? mem[2926] : 
                        (N174)? mem[3006] : 
                        (N176)? mem[3086] : 
                        (N178)? mem[3166] : 
                        (N180)? mem[3246] : 
                        (N182)? mem[3326] : 
                        (N184)? mem[3406] : 
                        (N186)? mem[3486] : 
                        (N188)? mem[3566] : 
                        (N190)? mem[3646] : 
                        (N192)? mem[3726] : 
                        (N194)? mem[3806] : 
                        (N196)? mem[3886] : 
                        (N198)? mem[3966] : 
                        (N200)? mem[4046] : 
                        (N202)? mem[4126] : 
                        (N204)? mem[4206] : 
                        (N206)? mem[4286] : 
                        (N208)? mem[4366] : 
                        (N210)? mem[4446] : 
                        (N212)? mem[4526] : 
                        (N214)? mem[4606] : 
                        (N216)? mem[4686] : 
                        (N218)? mem[4766] : 
                        (N220)? mem[4846] : 
                        (N222)? mem[4926] : 
                        (N224)? mem[5006] : 
                        (N226)? mem[5086] : 1'b0;
  assign data_out[45] = (N163)? mem[45] : 
                        (N165)? mem[125] : 
                        (N167)? mem[205] : 
                        (N169)? mem[285] : 
                        (N171)? mem[365] : 
                        (N173)? mem[445] : 
                        (N175)? mem[525] : 
                        (N177)? mem[605] : 
                        (N179)? mem[685] : 
                        (N181)? mem[765] : 
                        (N183)? mem[845] : 
                        (N185)? mem[925] : 
                        (N187)? mem[1005] : 
                        (N189)? mem[1085] : 
                        (N191)? mem[1165] : 
                        (N193)? mem[1245] : 
                        (N195)? mem[1325] : 
                        (N197)? mem[1405] : 
                        (N199)? mem[1485] : 
                        (N201)? mem[1565] : 
                        (N203)? mem[1645] : 
                        (N205)? mem[1725] : 
                        (N207)? mem[1805] : 
                        (N209)? mem[1885] : 
                        (N211)? mem[1965] : 
                        (N213)? mem[2045] : 
                        (N215)? mem[2125] : 
                        (N217)? mem[2205] : 
                        (N219)? mem[2285] : 
                        (N221)? mem[2365] : 
                        (N223)? mem[2445] : 
                        (N225)? mem[2525] : 
                        (N164)? mem[2605] : 
                        (N166)? mem[2685] : 
                        (N168)? mem[2765] : 
                        (N170)? mem[2845] : 
                        (N172)? mem[2925] : 
                        (N174)? mem[3005] : 
                        (N176)? mem[3085] : 
                        (N178)? mem[3165] : 
                        (N180)? mem[3245] : 
                        (N182)? mem[3325] : 
                        (N184)? mem[3405] : 
                        (N186)? mem[3485] : 
                        (N188)? mem[3565] : 
                        (N190)? mem[3645] : 
                        (N192)? mem[3725] : 
                        (N194)? mem[3805] : 
                        (N196)? mem[3885] : 
                        (N198)? mem[3965] : 
                        (N200)? mem[4045] : 
                        (N202)? mem[4125] : 
                        (N204)? mem[4205] : 
                        (N206)? mem[4285] : 
                        (N208)? mem[4365] : 
                        (N210)? mem[4445] : 
                        (N212)? mem[4525] : 
                        (N214)? mem[4605] : 
                        (N216)? mem[4685] : 
                        (N218)? mem[4765] : 
                        (N220)? mem[4845] : 
                        (N222)? mem[4925] : 
                        (N224)? mem[5005] : 
                        (N226)? mem[5085] : 1'b0;
  assign data_out[44] = (N163)? mem[44] : 
                        (N165)? mem[124] : 
                        (N167)? mem[204] : 
                        (N169)? mem[284] : 
                        (N171)? mem[364] : 
                        (N173)? mem[444] : 
                        (N175)? mem[524] : 
                        (N177)? mem[604] : 
                        (N179)? mem[684] : 
                        (N181)? mem[764] : 
                        (N183)? mem[844] : 
                        (N185)? mem[924] : 
                        (N187)? mem[1004] : 
                        (N189)? mem[1084] : 
                        (N191)? mem[1164] : 
                        (N193)? mem[1244] : 
                        (N195)? mem[1324] : 
                        (N197)? mem[1404] : 
                        (N199)? mem[1484] : 
                        (N201)? mem[1564] : 
                        (N203)? mem[1644] : 
                        (N205)? mem[1724] : 
                        (N207)? mem[1804] : 
                        (N209)? mem[1884] : 
                        (N211)? mem[1964] : 
                        (N213)? mem[2044] : 
                        (N215)? mem[2124] : 
                        (N217)? mem[2204] : 
                        (N219)? mem[2284] : 
                        (N221)? mem[2364] : 
                        (N223)? mem[2444] : 
                        (N225)? mem[2524] : 
                        (N164)? mem[2604] : 
                        (N166)? mem[2684] : 
                        (N168)? mem[2764] : 
                        (N170)? mem[2844] : 
                        (N172)? mem[2924] : 
                        (N174)? mem[3004] : 
                        (N176)? mem[3084] : 
                        (N178)? mem[3164] : 
                        (N180)? mem[3244] : 
                        (N182)? mem[3324] : 
                        (N184)? mem[3404] : 
                        (N186)? mem[3484] : 
                        (N188)? mem[3564] : 
                        (N190)? mem[3644] : 
                        (N192)? mem[3724] : 
                        (N194)? mem[3804] : 
                        (N196)? mem[3884] : 
                        (N198)? mem[3964] : 
                        (N200)? mem[4044] : 
                        (N202)? mem[4124] : 
                        (N204)? mem[4204] : 
                        (N206)? mem[4284] : 
                        (N208)? mem[4364] : 
                        (N210)? mem[4444] : 
                        (N212)? mem[4524] : 
                        (N214)? mem[4604] : 
                        (N216)? mem[4684] : 
                        (N218)? mem[4764] : 
                        (N220)? mem[4844] : 
                        (N222)? mem[4924] : 
                        (N224)? mem[5004] : 
                        (N226)? mem[5084] : 1'b0;
  assign data_out[43] = (N163)? mem[43] : 
                        (N165)? mem[123] : 
                        (N167)? mem[203] : 
                        (N169)? mem[283] : 
                        (N171)? mem[363] : 
                        (N173)? mem[443] : 
                        (N175)? mem[523] : 
                        (N177)? mem[603] : 
                        (N179)? mem[683] : 
                        (N181)? mem[763] : 
                        (N183)? mem[843] : 
                        (N185)? mem[923] : 
                        (N187)? mem[1003] : 
                        (N189)? mem[1083] : 
                        (N191)? mem[1163] : 
                        (N193)? mem[1243] : 
                        (N195)? mem[1323] : 
                        (N197)? mem[1403] : 
                        (N199)? mem[1483] : 
                        (N201)? mem[1563] : 
                        (N203)? mem[1643] : 
                        (N205)? mem[1723] : 
                        (N207)? mem[1803] : 
                        (N209)? mem[1883] : 
                        (N211)? mem[1963] : 
                        (N213)? mem[2043] : 
                        (N215)? mem[2123] : 
                        (N217)? mem[2203] : 
                        (N219)? mem[2283] : 
                        (N221)? mem[2363] : 
                        (N223)? mem[2443] : 
                        (N225)? mem[2523] : 
                        (N164)? mem[2603] : 
                        (N166)? mem[2683] : 
                        (N168)? mem[2763] : 
                        (N170)? mem[2843] : 
                        (N172)? mem[2923] : 
                        (N174)? mem[3003] : 
                        (N176)? mem[3083] : 
                        (N178)? mem[3163] : 
                        (N180)? mem[3243] : 
                        (N182)? mem[3323] : 
                        (N184)? mem[3403] : 
                        (N186)? mem[3483] : 
                        (N188)? mem[3563] : 
                        (N190)? mem[3643] : 
                        (N192)? mem[3723] : 
                        (N194)? mem[3803] : 
                        (N196)? mem[3883] : 
                        (N198)? mem[3963] : 
                        (N200)? mem[4043] : 
                        (N202)? mem[4123] : 
                        (N204)? mem[4203] : 
                        (N206)? mem[4283] : 
                        (N208)? mem[4363] : 
                        (N210)? mem[4443] : 
                        (N212)? mem[4523] : 
                        (N214)? mem[4603] : 
                        (N216)? mem[4683] : 
                        (N218)? mem[4763] : 
                        (N220)? mem[4843] : 
                        (N222)? mem[4923] : 
                        (N224)? mem[5003] : 
                        (N226)? mem[5083] : 1'b0;
  assign data_out[42] = (N163)? mem[42] : 
                        (N165)? mem[122] : 
                        (N167)? mem[202] : 
                        (N169)? mem[282] : 
                        (N171)? mem[362] : 
                        (N173)? mem[442] : 
                        (N175)? mem[522] : 
                        (N177)? mem[602] : 
                        (N179)? mem[682] : 
                        (N181)? mem[762] : 
                        (N183)? mem[842] : 
                        (N185)? mem[922] : 
                        (N187)? mem[1002] : 
                        (N189)? mem[1082] : 
                        (N191)? mem[1162] : 
                        (N193)? mem[1242] : 
                        (N195)? mem[1322] : 
                        (N197)? mem[1402] : 
                        (N199)? mem[1482] : 
                        (N201)? mem[1562] : 
                        (N203)? mem[1642] : 
                        (N205)? mem[1722] : 
                        (N207)? mem[1802] : 
                        (N209)? mem[1882] : 
                        (N211)? mem[1962] : 
                        (N213)? mem[2042] : 
                        (N215)? mem[2122] : 
                        (N217)? mem[2202] : 
                        (N219)? mem[2282] : 
                        (N221)? mem[2362] : 
                        (N223)? mem[2442] : 
                        (N225)? mem[2522] : 
                        (N164)? mem[2602] : 
                        (N166)? mem[2682] : 
                        (N168)? mem[2762] : 
                        (N170)? mem[2842] : 
                        (N172)? mem[2922] : 
                        (N174)? mem[3002] : 
                        (N176)? mem[3082] : 
                        (N178)? mem[3162] : 
                        (N180)? mem[3242] : 
                        (N182)? mem[3322] : 
                        (N184)? mem[3402] : 
                        (N186)? mem[3482] : 
                        (N188)? mem[3562] : 
                        (N190)? mem[3642] : 
                        (N192)? mem[3722] : 
                        (N194)? mem[3802] : 
                        (N196)? mem[3882] : 
                        (N198)? mem[3962] : 
                        (N200)? mem[4042] : 
                        (N202)? mem[4122] : 
                        (N204)? mem[4202] : 
                        (N206)? mem[4282] : 
                        (N208)? mem[4362] : 
                        (N210)? mem[4442] : 
                        (N212)? mem[4522] : 
                        (N214)? mem[4602] : 
                        (N216)? mem[4682] : 
                        (N218)? mem[4762] : 
                        (N220)? mem[4842] : 
                        (N222)? mem[4922] : 
                        (N224)? mem[5002] : 
                        (N226)? mem[5082] : 1'b0;
  assign data_out[41] = (N163)? mem[41] : 
                        (N165)? mem[121] : 
                        (N167)? mem[201] : 
                        (N169)? mem[281] : 
                        (N171)? mem[361] : 
                        (N173)? mem[441] : 
                        (N175)? mem[521] : 
                        (N177)? mem[601] : 
                        (N179)? mem[681] : 
                        (N181)? mem[761] : 
                        (N183)? mem[841] : 
                        (N185)? mem[921] : 
                        (N187)? mem[1001] : 
                        (N189)? mem[1081] : 
                        (N191)? mem[1161] : 
                        (N193)? mem[1241] : 
                        (N195)? mem[1321] : 
                        (N197)? mem[1401] : 
                        (N199)? mem[1481] : 
                        (N201)? mem[1561] : 
                        (N203)? mem[1641] : 
                        (N205)? mem[1721] : 
                        (N207)? mem[1801] : 
                        (N209)? mem[1881] : 
                        (N211)? mem[1961] : 
                        (N213)? mem[2041] : 
                        (N215)? mem[2121] : 
                        (N217)? mem[2201] : 
                        (N219)? mem[2281] : 
                        (N221)? mem[2361] : 
                        (N223)? mem[2441] : 
                        (N225)? mem[2521] : 
                        (N164)? mem[2601] : 
                        (N166)? mem[2681] : 
                        (N168)? mem[2761] : 
                        (N170)? mem[2841] : 
                        (N172)? mem[2921] : 
                        (N174)? mem[3001] : 
                        (N176)? mem[3081] : 
                        (N178)? mem[3161] : 
                        (N180)? mem[3241] : 
                        (N182)? mem[3321] : 
                        (N184)? mem[3401] : 
                        (N186)? mem[3481] : 
                        (N188)? mem[3561] : 
                        (N190)? mem[3641] : 
                        (N192)? mem[3721] : 
                        (N194)? mem[3801] : 
                        (N196)? mem[3881] : 
                        (N198)? mem[3961] : 
                        (N200)? mem[4041] : 
                        (N202)? mem[4121] : 
                        (N204)? mem[4201] : 
                        (N206)? mem[4281] : 
                        (N208)? mem[4361] : 
                        (N210)? mem[4441] : 
                        (N212)? mem[4521] : 
                        (N214)? mem[4601] : 
                        (N216)? mem[4681] : 
                        (N218)? mem[4761] : 
                        (N220)? mem[4841] : 
                        (N222)? mem[4921] : 
                        (N224)? mem[5001] : 
                        (N226)? mem[5081] : 1'b0;
  assign data_out[40] = (N163)? mem[40] : 
                        (N165)? mem[120] : 
                        (N167)? mem[200] : 
                        (N169)? mem[280] : 
                        (N171)? mem[360] : 
                        (N173)? mem[440] : 
                        (N175)? mem[520] : 
                        (N177)? mem[600] : 
                        (N179)? mem[680] : 
                        (N181)? mem[760] : 
                        (N183)? mem[840] : 
                        (N185)? mem[920] : 
                        (N187)? mem[1000] : 
                        (N189)? mem[1080] : 
                        (N191)? mem[1160] : 
                        (N193)? mem[1240] : 
                        (N195)? mem[1320] : 
                        (N197)? mem[1400] : 
                        (N199)? mem[1480] : 
                        (N201)? mem[1560] : 
                        (N203)? mem[1640] : 
                        (N205)? mem[1720] : 
                        (N207)? mem[1800] : 
                        (N209)? mem[1880] : 
                        (N211)? mem[1960] : 
                        (N213)? mem[2040] : 
                        (N215)? mem[2120] : 
                        (N217)? mem[2200] : 
                        (N219)? mem[2280] : 
                        (N221)? mem[2360] : 
                        (N223)? mem[2440] : 
                        (N225)? mem[2520] : 
                        (N164)? mem[2600] : 
                        (N166)? mem[2680] : 
                        (N168)? mem[2760] : 
                        (N170)? mem[2840] : 
                        (N172)? mem[2920] : 
                        (N174)? mem[3000] : 
                        (N176)? mem[3080] : 
                        (N178)? mem[3160] : 
                        (N180)? mem[3240] : 
                        (N182)? mem[3320] : 
                        (N184)? mem[3400] : 
                        (N186)? mem[3480] : 
                        (N188)? mem[3560] : 
                        (N190)? mem[3640] : 
                        (N192)? mem[3720] : 
                        (N194)? mem[3800] : 
                        (N196)? mem[3880] : 
                        (N198)? mem[3960] : 
                        (N200)? mem[4040] : 
                        (N202)? mem[4120] : 
                        (N204)? mem[4200] : 
                        (N206)? mem[4280] : 
                        (N208)? mem[4360] : 
                        (N210)? mem[4440] : 
                        (N212)? mem[4520] : 
                        (N214)? mem[4600] : 
                        (N216)? mem[4680] : 
                        (N218)? mem[4760] : 
                        (N220)? mem[4840] : 
                        (N222)? mem[4920] : 
                        (N224)? mem[5000] : 
                        (N226)? mem[5080] : 1'b0;
  assign data_out[39] = (N163)? mem[39] : 
                        (N165)? mem[119] : 
                        (N167)? mem[199] : 
                        (N169)? mem[279] : 
                        (N171)? mem[359] : 
                        (N173)? mem[439] : 
                        (N175)? mem[519] : 
                        (N177)? mem[599] : 
                        (N179)? mem[679] : 
                        (N181)? mem[759] : 
                        (N183)? mem[839] : 
                        (N185)? mem[919] : 
                        (N187)? mem[999] : 
                        (N189)? mem[1079] : 
                        (N191)? mem[1159] : 
                        (N193)? mem[1239] : 
                        (N195)? mem[1319] : 
                        (N197)? mem[1399] : 
                        (N199)? mem[1479] : 
                        (N201)? mem[1559] : 
                        (N203)? mem[1639] : 
                        (N205)? mem[1719] : 
                        (N207)? mem[1799] : 
                        (N209)? mem[1879] : 
                        (N211)? mem[1959] : 
                        (N213)? mem[2039] : 
                        (N215)? mem[2119] : 
                        (N217)? mem[2199] : 
                        (N219)? mem[2279] : 
                        (N221)? mem[2359] : 
                        (N223)? mem[2439] : 
                        (N225)? mem[2519] : 
                        (N164)? mem[2599] : 
                        (N166)? mem[2679] : 
                        (N168)? mem[2759] : 
                        (N170)? mem[2839] : 
                        (N172)? mem[2919] : 
                        (N174)? mem[2999] : 
                        (N176)? mem[3079] : 
                        (N178)? mem[3159] : 
                        (N180)? mem[3239] : 
                        (N182)? mem[3319] : 
                        (N184)? mem[3399] : 
                        (N186)? mem[3479] : 
                        (N188)? mem[3559] : 
                        (N190)? mem[3639] : 
                        (N192)? mem[3719] : 
                        (N194)? mem[3799] : 
                        (N196)? mem[3879] : 
                        (N198)? mem[3959] : 
                        (N200)? mem[4039] : 
                        (N202)? mem[4119] : 
                        (N204)? mem[4199] : 
                        (N206)? mem[4279] : 
                        (N208)? mem[4359] : 
                        (N210)? mem[4439] : 
                        (N212)? mem[4519] : 
                        (N214)? mem[4599] : 
                        (N216)? mem[4679] : 
                        (N218)? mem[4759] : 
                        (N220)? mem[4839] : 
                        (N222)? mem[4919] : 
                        (N224)? mem[4999] : 
                        (N226)? mem[5079] : 1'b0;
  assign data_out[38] = (N163)? mem[38] : 
                        (N165)? mem[118] : 
                        (N167)? mem[198] : 
                        (N169)? mem[278] : 
                        (N171)? mem[358] : 
                        (N173)? mem[438] : 
                        (N175)? mem[518] : 
                        (N177)? mem[598] : 
                        (N179)? mem[678] : 
                        (N181)? mem[758] : 
                        (N183)? mem[838] : 
                        (N185)? mem[918] : 
                        (N187)? mem[998] : 
                        (N189)? mem[1078] : 
                        (N191)? mem[1158] : 
                        (N193)? mem[1238] : 
                        (N195)? mem[1318] : 
                        (N197)? mem[1398] : 
                        (N199)? mem[1478] : 
                        (N201)? mem[1558] : 
                        (N203)? mem[1638] : 
                        (N205)? mem[1718] : 
                        (N207)? mem[1798] : 
                        (N209)? mem[1878] : 
                        (N211)? mem[1958] : 
                        (N213)? mem[2038] : 
                        (N215)? mem[2118] : 
                        (N217)? mem[2198] : 
                        (N219)? mem[2278] : 
                        (N221)? mem[2358] : 
                        (N223)? mem[2438] : 
                        (N225)? mem[2518] : 
                        (N164)? mem[2598] : 
                        (N166)? mem[2678] : 
                        (N168)? mem[2758] : 
                        (N170)? mem[2838] : 
                        (N172)? mem[2918] : 
                        (N174)? mem[2998] : 
                        (N176)? mem[3078] : 
                        (N178)? mem[3158] : 
                        (N180)? mem[3238] : 
                        (N182)? mem[3318] : 
                        (N184)? mem[3398] : 
                        (N186)? mem[3478] : 
                        (N188)? mem[3558] : 
                        (N190)? mem[3638] : 
                        (N192)? mem[3718] : 
                        (N194)? mem[3798] : 
                        (N196)? mem[3878] : 
                        (N198)? mem[3958] : 
                        (N200)? mem[4038] : 
                        (N202)? mem[4118] : 
                        (N204)? mem[4198] : 
                        (N206)? mem[4278] : 
                        (N208)? mem[4358] : 
                        (N210)? mem[4438] : 
                        (N212)? mem[4518] : 
                        (N214)? mem[4598] : 
                        (N216)? mem[4678] : 
                        (N218)? mem[4758] : 
                        (N220)? mem[4838] : 
                        (N222)? mem[4918] : 
                        (N224)? mem[4998] : 
                        (N226)? mem[5078] : 1'b0;
  assign data_out[37] = (N163)? mem[37] : 
                        (N165)? mem[117] : 
                        (N167)? mem[197] : 
                        (N169)? mem[277] : 
                        (N171)? mem[357] : 
                        (N173)? mem[437] : 
                        (N175)? mem[517] : 
                        (N177)? mem[597] : 
                        (N179)? mem[677] : 
                        (N181)? mem[757] : 
                        (N183)? mem[837] : 
                        (N185)? mem[917] : 
                        (N187)? mem[997] : 
                        (N189)? mem[1077] : 
                        (N191)? mem[1157] : 
                        (N193)? mem[1237] : 
                        (N195)? mem[1317] : 
                        (N197)? mem[1397] : 
                        (N199)? mem[1477] : 
                        (N201)? mem[1557] : 
                        (N203)? mem[1637] : 
                        (N205)? mem[1717] : 
                        (N207)? mem[1797] : 
                        (N209)? mem[1877] : 
                        (N211)? mem[1957] : 
                        (N213)? mem[2037] : 
                        (N215)? mem[2117] : 
                        (N217)? mem[2197] : 
                        (N219)? mem[2277] : 
                        (N221)? mem[2357] : 
                        (N223)? mem[2437] : 
                        (N225)? mem[2517] : 
                        (N164)? mem[2597] : 
                        (N166)? mem[2677] : 
                        (N168)? mem[2757] : 
                        (N170)? mem[2837] : 
                        (N172)? mem[2917] : 
                        (N174)? mem[2997] : 
                        (N176)? mem[3077] : 
                        (N178)? mem[3157] : 
                        (N180)? mem[3237] : 
                        (N182)? mem[3317] : 
                        (N184)? mem[3397] : 
                        (N186)? mem[3477] : 
                        (N188)? mem[3557] : 
                        (N190)? mem[3637] : 
                        (N192)? mem[3717] : 
                        (N194)? mem[3797] : 
                        (N196)? mem[3877] : 
                        (N198)? mem[3957] : 
                        (N200)? mem[4037] : 
                        (N202)? mem[4117] : 
                        (N204)? mem[4197] : 
                        (N206)? mem[4277] : 
                        (N208)? mem[4357] : 
                        (N210)? mem[4437] : 
                        (N212)? mem[4517] : 
                        (N214)? mem[4597] : 
                        (N216)? mem[4677] : 
                        (N218)? mem[4757] : 
                        (N220)? mem[4837] : 
                        (N222)? mem[4917] : 
                        (N224)? mem[4997] : 
                        (N226)? mem[5077] : 1'b0;
  assign data_out[36] = (N163)? mem[36] : 
                        (N165)? mem[116] : 
                        (N167)? mem[196] : 
                        (N169)? mem[276] : 
                        (N171)? mem[356] : 
                        (N173)? mem[436] : 
                        (N175)? mem[516] : 
                        (N177)? mem[596] : 
                        (N179)? mem[676] : 
                        (N181)? mem[756] : 
                        (N183)? mem[836] : 
                        (N185)? mem[916] : 
                        (N187)? mem[996] : 
                        (N189)? mem[1076] : 
                        (N191)? mem[1156] : 
                        (N193)? mem[1236] : 
                        (N195)? mem[1316] : 
                        (N197)? mem[1396] : 
                        (N199)? mem[1476] : 
                        (N201)? mem[1556] : 
                        (N203)? mem[1636] : 
                        (N205)? mem[1716] : 
                        (N207)? mem[1796] : 
                        (N209)? mem[1876] : 
                        (N211)? mem[1956] : 
                        (N213)? mem[2036] : 
                        (N215)? mem[2116] : 
                        (N217)? mem[2196] : 
                        (N219)? mem[2276] : 
                        (N221)? mem[2356] : 
                        (N223)? mem[2436] : 
                        (N225)? mem[2516] : 
                        (N164)? mem[2596] : 
                        (N166)? mem[2676] : 
                        (N168)? mem[2756] : 
                        (N170)? mem[2836] : 
                        (N172)? mem[2916] : 
                        (N174)? mem[2996] : 
                        (N176)? mem[3076] : 
                        (N178)? mem[3156] : 
                        (N180)? mem[3236] : 
                        (N182)? mem[3316] : 
                        (N184)? mem[3396] : 
                        (N186)? mem[3476] : 
                        (N188)? mem[3556] : 
                        (N190)? mem[3636] : 
                        (N192)? mem[3716] : 
                        (N194)? mem[3796] : 
                        (N196)? mem[3876] : 
                        (N198)? mem[3956] : 
                        (N200)? mem[4036] : 
                        (N202)? mem[4116] : 
                        (N204)? mem[4196] : 
                        (N206)? mem[4276] : 
                        (N208)? mem[4356] : 
                        (N210)? mem[4436] : 
                        (N212)? mem[4516] : 
                        (N214)? mem[4596] : 
                        (N216)? mem[4676] : 
                        (N218)? mem[4756] : 
                        (N220)? mem[4836] : 
                        (N222)? mem[4916] : 
                        (N224)? mem[4996] : 
                        (N226)? mem[5076] : 1'b0;
  assign data_out[35] = (N163)? mem[35] : 
                        (N165)? mem[115] : 
                        (N167)? mem[195] : 
                        (N169)? mem[275] : 
                        (N171)? mem[355] : 
                        (N173)? mem[435] : 
                        (N175)? mem[515] : 
                        (N177)? mem[595] : 
                        (N179)? mem[675] : 
                        (N181)? mem[755] : 
                        (N183)? mem[835] : 
                        (N185)? mem[915] : 
                        (N187)? mem[995] : 
                        (N189)? mem[1075] : 
                        (N191)? mem[1155] : 
                        (N193)? mem[1235] : 
                        (N195)? mem[1315] : 
                        (N197)? mem[1395] : 
                        (N199)? mem[1475] : 
                        (N201)? mem[1555] : 
                        (N203)? mem[1635] : 
                        (N205)? mem[1715] : 
                        (N207)? mem[1795] : 
                        (N209)? mem[1875] : 
                        (N211)? mem[1955] : 
                        (N213)? mem[2035] : 
                        (N215)? mem[2115] : 
                        (N217)? mem[2195] : 
                        (N219)? mem[2275] : 
                        (N221)? mem[2355] : 
                        (N223)? mem[2435] : 
                        (N225)? mem[2515] : 
                        (N164)? mem[2595] : 
                        (N166)? mem[2675] : 
                        (N168)? mem[2755] : 
                        (N170)? mem[2835] : 
                        (N172)? mem[2915] : 
                        (N174)? mem[2995] : 
                        (N176)? mem[3075] : 
                        (N178)? mem[3155] : 
                        (N180)? mem[3235] : 
                        (N182)? mem[3315] : 
                        (N184)? mem[3395] : 
                        (N186)? mem[3475] : 
                        (N188)? mem[3555] : 
                        (N190)? mem[3635] : 
                        (N192)? mem[3715] : 
                        (N194)? mem[3795] : 
                        (N196)? mem[3875] : 
                        (N198)? mem[3955] : 
                        (N200)? mem[4035] : 
                        (N202)? mem[4115] : 
                        (N204)? mem[4195] : 
                        (N206)? mem[4275] : 
                        (N208)? mem[4355] : 
                        (N210)? mem[4435] : 
                        (N212)? mem[4515] : 
                        (N214)? mem[4595] : 
                        (N216)? mem[4675] : 
                        (N218)? mem[4755] : 
                        (N220)? mem[4835] : 
                        (N222)? mem[4915] : 
                        (N224)? mem[4995] : 
                        (N226)? mem[5075] : 1'b0;
  assign data_out[34] = (N163)? mem[34] : 
                        (N165)? mem[114] : 
                        (N167)? mem[194] : 
                        (N169)? mem[274] : 
                        (N171)? mem[354] : 
                        (N173)? mem[434] : 
                        (N175)? mem[514] : 
                        (N177)? mem[594] : 
                        (N179)? mem[674] : 
                        (N181)? mem[754] : 
                        (N183)? mem[834] : 
                        (N185)? mem[914] : 
                        (N187)? mem[994] : 
                        (N189)? mem[1074] : 
                        (N191)? mem[1154] : 
                        (N193)? mem[1234] : 
                        (N195)? mem[1314] : 
                        (N197)? mem[1394] : 
                        (N199)? mem[1474] : 
                        (N201)? mem[1554] : 
                        (N203)? mem[1634] : 
                        (N205)? mem[1714] : 
                        (N207)? mem[1794] : 
                        (N209)? mem[1874] : 
                        (N211)? mem[1954] : 
                        (N213)? mem[2034] : 
                        (N215)? mem[2114] : 
                        (N217)? mem[2194] : 
                        (N219)? mem[2274] : 
                        (N221)? mem[2354] : 
                        (N223)? mem[2434] : 
                        (N225)? mem[2514] : 
                        (N164)? mem[2594] : 
                        (N166)? mem[2674] : 
                        (N168)? mem[2754] : 
                        (N170)? mem[2834] : 
                        (N172)? mem[2914] : 
                        (N174)? mem[2994] : 
                        (N176)? mem[3074] : 
                        (N178)? mem[3154] : 
                        (N180)? mem[3234] : 
                        (N182)? mem[3314] : 
                        (N184)? mem[3394] : 
                        (N186)? mem[3474] : 
                        (N188)? mem[3554] : 
                        (N190)? mem[3634] : 
                        (N192)? mem[3714] : 
                        (N194)? mem[3794] : 
                        (N196)? mem[3874] : 
                        (N198)? mem[3954] : 
                        (N200)? mem[4034] : 
                        (N202)? mem[4114] : 
                        (N204)? mem[4194] : 
                        (N206)? mem[4274] : 
                        (N208)? mem[4354] : 
                        (N210)? mem[4434] : 
                        (N212)? mem[4514] : 
                        (N214)? mem[4594] : 
                        (N216)? mem[4674] : 
                        (N218)? mem[4754] : 
                        (N220)? mem[4834] : 
                        (N222)? mem[4914] : 
                        (N224)? mem[4994] : 
                        (N226)? mem[5074] : 1'b0;
  assign data_out[33] = (N163)? mem[33] : 
                        (N165)? mem[113] : 
                        (N167)? mem[193] : 
                        (N169)? mem[273] : 
                        (N171)? mem[353] : 
                        (N173)? mem[433] : 
                        (N175)? mem[513] : 
                        (N177)? mem[593] : 
                        (N179)? mem[673] : 
                        (N181)? mem[753] : 
                        (N183)? mem[833] : 
                        (N185)? mem[913] : 
                        (N187)? mem[993] : 
                        (N189)? mem[1073] : 
                        (N191)? mem[1153] : 
                        (N193)? mem[1233] : 
                        (N195)? mem[1313] : 
                        (N197)? mem[1393] : 
                        (N199)? mem[1473] : 
                        (N201)? mem[1553] : 
                        (N203)? mem[1633] : 
                        (N205)? mem[1713] : 
                        (N207)? mem[1793] : 
                        (N209)? mem[1873] : 
                        (N211)? mem[1953] : 
                        (N213)? mem[2033] : 
                        (N215)? mem[2113] : 
                        (N217)? mem[2193] : 
                        (N219)? mem[2273] : 
                        (N221)? mem[2353] : 
                        (N223)? mem[2433] : 
                        (N225)? mem[2513] : 
                        (N164)? mem[2593] : 
                        (N166)? mem[2673] : 
                        (N168)? mem[2753] : 
                        (N170)? mem[2833] : 
                        (N172)? mem[2913] : 
                        (N174)? mem[2993] : 
                        (N176)? mem[3073] : 
                        (N178)? mem[3153] : 
                        (N180)? mem[3233] : 
                        (N182)? mem[3313] : 
                        (N184)? mem[3393] : 
                        (N186)? mem[3473] : 
                        (N188)? mem[3553] : 
                        (N190)? mem[3633] : 
                        (N192)? mem[3713] : 
                        (N194)? mem[3793] : 
                        (N196)? mem[3873] : 
                        (N198)? mem[3953] : 
                        (N200)? mem[4033] : 
                        (N202)? mem[4113] : 
                        (N204)? mem[4193] : 
                        (N206)? mem[4273] : 
                        (N208)? mem[4353] : 
                        (N210)? mem[4433] : 
                        (N212)? mem[4513] : 
                        (N214)? mem[4593] : 
                        (N216)? mem[4673] : 
                        (N218)? mem[4753] : 
                        (N220)? mem[4833] : 
                        (N222)? mem[4913] : 
                        (N224)? mem[4993] : 
                        (N226)? mem[5073] : 1'b0;
  assign data_out[32] = (N163)? mem[32] : 
                        (N165)? mem[112] : 
                        (N167)? mem[192] : 
                        (N169)? mem[272] : 
                        (N171)? mem[352] : 
                        (N173)? mem[432] : 
                        (N175)? mem[512] : 
                        (N177)? mem[592] : 
                        (N179)? mem[672] : 
                        (N181)? mem[752] : 
                        (N183)? mem[832] : 
                        (N185)? mem[912] : 
                        (N187)? mem[992] : 
                        (N189)? mem[1072] : 
                        (N191)? mem[1152] : 
                        (N193)? mem[1232] : 
                        (N195)? mem[1312] : 
                        (N197)? mem[1392] : 
                        (N199)? mem[1472] : 
                        (N201)? mem[1552] : 
                        (N203)? mem[1632] : 
                        (N205)? mem[1712] : 
                        (N207)? mem[1792] : 
                        (N209)? mem[1872] : 
                        (N211)? mem[1952] : 
                        (N213)? mem[2032] : 
                        (N215)? mem[2112] : 
                        (N217)? mem[2192] : 
                        (N219)? mem[2272] : 
                        (N221)? mem[2352] : 
                        (N223)? mem[2432] : 
                        (N225)? mem[2512] : 
                        (N164)? mem[2592] : 
                        (N166)? mem[2672] : 
                        (N168)? mem[2752] : 
                        (N170)? mem[2832] : 
                        (N172)? mem[2912] : 
                        (N174)? mem[2992] : 
                        (N176)? mem[3072] : 
                        (N178)? mem[3152] : 
                        (N180)? mem[3232] : 
                        (N182)? mem[3312] : 
                        (N184)? mem[3392] : 
                        (N186)? mem[3472] : 
                        (N188)? mem[3552] : 
                        (N190)? mem[3632] : 
                        (N192)? mem[3712] : 
                        (N194)? mem[3792] : 
                        (N196)? mem[3872] : 
                        (N198)? mem[3952] : 
                        (N200)? mem[4032] : 
                        (N202)? mem[4112] : 
                        (N204)? mem[4192] : 
                        (N206)? mem[4272] : 
                        (N208)? mem[4352] : 
                        (N210)? mem[4432] : 
                        (N212)? mem[4512] : 
                        (N214)? mem[4592] : 
                        (N216)? mem[4672] : 
                        (N218)? mem[4752] : 
                        (N220)? mem[4832] : 
                        (N222)? mem[4912] : 
                        (N224)? mem[4992] : 
                        (N226)? mem[5072] : 1'b0;
  assign data_out[31] = (N163)? mem[31] : 
                        (N165)? mem[111] : 
                        (N167)? mem[191] : 
                        (N169)? mem[271] : 
                        (N171)? mem[351] : 
                        (N173)? mem[431] : 
                        (N175)? mem[511] : 
                        (N177)? mem[591] : 
                        (N179)? mem[671] : 
                        (N181)? mem[751] : 
                        (N183)? mem[831] : 
                        (N185)? mem[911] : 
                        (N187)? mem[991] : 
                        (N189)? mem[1071] : 
                        (N191)? mem[1151] : 
                        (N193)? mem[1231] : 
                        (N195)? mem[1311] : 
                        (N197)? mem[1391] : 
                        (N199)? mem[1471] : 
                        (N201)? mem[1551] : 
                        (N203)? mem[1631] : 
                        (N205)? mem[1711] : 
                        (N207)? mem[1791] : 
                        (N209)? mem[1871] : 
                        (N211)? mem[1951] : 
                        (N213)? mem[2031] : 
                        (N215)? mem[2111] : 
                        (N217)? mem[2191] : 
                        (N219)? mem[2271] : 
                        (N221)? mem[2351] : 
                        (N223)? mem[2431] : 
                        (N225)? mem[2511] : 
                        (N164)? mem[2591] : 
                        (N166)? mem[2671] : 
                        (N168)? mem[2751] : 
                        (N170)? mem[2831] : 
                        (N172)? mem[2911] : 
                        (N174)? mem[2991] : 
                        (N176)? mem[3071] : 
                        (N178)? mem[3151] : 
                        (N180)? mem[3231] : 
                        (N182)? mem[3311] : 
                        (N184)? mem[3391] : 
                        (N186)? mem[3471] : 
                        (N188)? mem[3551] : 
                        (N190)? mem[3631] : 
                        (N192)? mem[3711] : 
                        (N194)? mem[3791] : 
                        (N196)? mem[3871] : 
                        (N198)? mem[3951] : 
                        (N200)? mem[4031] : 
                        (N202)? mem[4111] : 
                        (N204)? mem[4191] : 
                        (N206)? mem[4271] : 
                        (N208)? mem[4351] : 
                        (N210)? mem[4431] : 
                        (N212)? mem[4511] : 
                        (N214)? mem[4591] : 
                        (N216)? mem[4671] : 
                        (N218)? mem[4751] : 
                        (N220)? mem[4831] : 
                        (N222)? mem[4911] : 
                        (N224)? mem[4991] : 
                        (N226)? mem[5071] : 1'b0;
  assign data_out[30] = (N163)? mem[30] : 
                        (N165)? mem[110] : 
                        (N167)? mem[190] : 
                        (N169)? mem[270] : 
                        (N171)? mem[350] : 
                        (N173)? mem[430] : 
                        (N175)? mem[510] : 
                        (N177)? mem[590] : 
                        (N179)? mem[670] : 
                        (N181)? mem[750] : 
                        (N183)? mem[830] : 
                        (N185)? mem[910] : 
                        (N187)? mem[990] : 
                        (N189)? mem[1070] : 
                        (N191)? mem[1150] : 
                        (N193)? mem[1230] : 
                        (N195)? mem[1310] : 
                        (N197)? mem[1390] : 
                        (N199)? mem[1470] : 
                        (N201)? mem[1550] : 
                        (N203)? mem[1630] : 
                        (N205)? mem[1710] : 
                        (N207)? mem[1790] : 
                        (N209)? mem[1870] : 
                        (N211)? mem[1950] : 
                        (N213)? mem[2030] : 
                        (N215)? mem[2110] : 
                        (N217)? mem[2190] : 
                        (N219)? mem[2270] : 
                        (N221)? mem[2350] : 
                        (N223)? mem[2430] : 
                        (N225)? mem[2510] : 
                        (N164)? mem[2590] : 
                        (N166)? mem[2670] : 
                        (N168)? mem[2750] : 
                        (N170)? mem[2830] : 
                        (N172)? mem[2910] : 
                        (N174)? mem[2990] : 
                        (N176)? mem[3070] : 
                        (N178)? mem[3150] : 
                        (N180)? mem[3230] : 
                        (N182)? mem[3310] : 
                        (N184)? mem[3390] : 
                        (N186)? mem[3470] : 
                        (N188)? mem[3550] : 
                        (N190)? mem[3630] : 
                        (N192)? mem[3710] : 
                        (N194)? mem[3790] : 
                        (N196)? mem[3870] : 
                        (N198)? mem[3950] : 
                        (N200)? mem[4030] : 
                        (N202)? mem[4110] : 
                        (N204)? mem[4190] : 
                        (N206)? mem[4270] : 
                        (N208)? mem[4350] : 
                        (N210)? mem[4430] : 
                        (N212)? mem[4510] : 
                        (N214)? mem[4590] : 
                        (N216)? mem[4670] : 
                        (N218)? mem[4750] : 
                        (N220)? mem[4830] : 
                        (N222)? mem[4910] : 
                        (N224)? mem[4990] : 
                        (N226)? mem[5070] : 1'b0;
  assign data_out[29] = (N163)? mem[29] : 
                        (N165)? mem[109] : 
                        (N167)? mem[189] : 
                        (N169)? mem[269] : 
                        (N171)? mem[349] : 
                        (N173)? mem[429] : 
                        (N175)? mem[509] : 
                        (N177)? mem[589] : 
                        (N179)? mem[669] : 
                        (N181)? mem[749] : 
                        (N183)? mem[829] : 
                        (N185)? mem[909] : 
                        (N187)? mem[989] : 
                        (N189)? mem[1069] : 
                        (N191)? mem[1149] : 
                        (N193)? mem[1229] : 
                        (N195)? mem[1309] : 
                        (N197)? mem[1389] : 
                        (N199)? mem[1469] : 
                        (N201)? mem[1549] : 
                        (N203)? mem[1629] : 
                        (N205)? mem[1709] : 
                        (N207)? mem[1789] : 
                        (N209)? mem[1869] : 
                        (N211)? mem[1949] : 
                        (N213)? mem[2029] : 
                        (N215)? mem[2109] : 
                        (N217)? mem[2189] : 
                        (N219)? mem[2269] : 
                        (N221)? mem[2349] : 
                        (N223)? mem[2429] : 
                        (N225)? mem[2509] : 
                        (N164)? mem[2589] : 
                        (N166)? mem[2669] : 
                        (N168)? mem[2749] : 
                        (N170)? mem[2829] : 
                        (N172)? mem[2909] : 
                        (N174)? mem[2989] : 
                        (N176)? mem[3069] : 
                        (N178)? mem[3149] : 
                        (N180)? mem[3229] : 
                        (N182)? mem[3309] : 
                        (N184)? mem[3389] : 
                        (N186)? mem[3469] : 
                        (N188)? mem[3549] : 
                        (N190)? mem[3629] : 
                        (N192)? mem[3709] : 
                        (N194)? mem[3789] : 
                        (N196)? mem[3869] : 
                        (N198)? mem[3949] : 
                        (N200)? mem[4029] : 
                        (N202)? mem[4109] : 
                        (N204)? mem[4189] : 
                        (N206)? mem[4269] : 
                        (N208)? mem[4349] : 
                        (N210)? mem[4429] : 
                        (N212)? mem[4509] : 
                        (N214)? mem[4589] : 
                        (N216)? mem[4669] : 
                        (N218)? mem[4749] : 
                        (N220)? mem[4829] : 
                        (N222)? mem[4909] : 
                        (N224)? mem[4989] : 
                        (N226)? mem[5069] : 1'b0;
  assign data_out[28] = (N163)? mem[28] : 
                        (N165)? mem[108] : 
                        (N167)? mem[188] : 
                        (N169)? mem[268] : 
                        (N171)? mem[348] : 
                        (N173)? mem[428] : 
                        (N175)? mem[508] : 
                        (N177)? mem[588] : 
                        (N179)? mem[668] : 
                        (N181)? mem[748] : 
                        (N183)? mem[828] : 
                        (N185)? mem[908] : 
                        (N187)? mem[988] : 
                        (N189)? mem[1068] : 
                        (N191)? mem[1148] : 
                        (N193)? mem[1228] : 
                        (N195)? mem[1308] : 
                        (N197)? mem[1388] : 
                        (N199)? mem[1468] : 
                        (N201)? mem[1548] : 
                        (N203)? mem[1628] : 
                        (N205)? mem[1708] : 
                        (N207)? mem[1788] : 
                        (N209)? mem[1868] : 
                        (N211)? mem[1948] : 
                        (N213)? mem[2028] : 
                        (N215)? mem[2108] : 
                        (N217)? mem[2188] : 
                        (N219)? mem[2268] : 
                        (N221)? mem[2348] : 
                        (N223)? mem[2428] : 
                        (N225)? mem[2508] : 
                        (N164)? mem[2588] : 
                        (N166)? mem[2668] : 
                        (N168)? mem[2748] : 
                        (N170)? mem[2828] : 
                        (N172)? mem[2908] : 
                        (N174)? mem[2988] : 
                        (N176)? mem[3068] : 
                        (N178)? mem[3148] : 
                        (N180)? mem[3228] : 
                        (N182)? mem[3308] : 
                        (N184)? mem[3388] : 
                        (N186)? mem[3468] : 
                        (N188)? mem[3548] : 
                        (N190)? mem[3628] : 
                        (N192)? mem[3708] : 
                        (N194)? mem[3788] : 
                        (N196)? mem[3868] : 
                        (N198)? mem[3948] : 
                        (N200)? mem[4028] : 
                        (N202)? mem[4108] : 
                        (N204)? mem[4188] : 
                        (N206)? mem[4268] : 
                        (N208)? mem[4348] : 
                        (N210)? mem[4428] : 
                        (N212)? mem[4508] : 
                        (N214)? mem[4588] : 
                        (N216)? mem[4668] : 
                        (N218)? mem[4748] : 
                        (N220)? mem[4828] : 
                        (N222)? mem[4908] : 
                        (N224)? mem[4988] : 
                        (N226)? mem[5068] : 1'b0;
  assign data_out[27] = (N163)? mem[27] : 
                        (N165)? mem[107] : 
                        (N167)? mem[187] : 
                        (N169)? mem[267] : 
                        (N171)? mem[347] : 
                        (N173)? mem[427] : 
                        (N175)? mem[507] : 
                        (N177)? mem[587] : 
                        (N179)? mem[667] : 
                        (N181)? mem[747] : 
                        (N183)? mem[827] : 
                        (N185)? mem[907] : 
                        (N187)? mem[987] : 
                        (N189)? mem[1067] : 
                        (N191)? mem[1147] : 
                        (N193)? mem[1227] : 
                        (N195)? mem[1307] : 
                        (N197)? mem[1387] : 
                        (N199)? mem[1467] : 
                        (N201)? mem[1547] : 
                        (N203)? mem[1627] : 
                        (N205)? mem[1707] : 
                        (N207)? mem[1787] : 
                        (N209)? mem[1867] : 
                        (N211)? mem[1947] : 
                        (N213)? mem[2027] : 
                        (N215)? mem[2107] : 
                        (N217)? mem[2187] : 
                        (N219)? mem[2267] : 
                        (N221)? mem[2347] : 
                        (N223)? mem[2427] : 
                        (N225)? mem[2507] : 
                        (N164)? mem[2587] : 
                        (N166)? mem[2667] : 
                        (N168)? mem[2747] : 
                        (N170)? mem[2827] : 
                        (N172)? mem[2907] : 
                        (N174)? mem[2987] : 
                        (N176)? mem[3067] : 
                        (N178)? mem[3147] : 
                        (N180)? mem[3227] : 
                        (N182)? mem[3307] : 
                        (N184)? mem[3387] : 
                        (N186)? mem[3467] : 
                        (N188)? mem[3547] : 
                        (N190)? mem[3627] : 
                        (N192)? mem[3707] : 
                        (N194)? mem[3787] : 
                        (N196)? mem[3867] : 
                        (N198)? mem[3947] : 
                        (N200)? mem[4027] : 
                        (N202)? mem[4107] : 
                        (N204)? mem[4187] : 
                        (N206)? mem[4267] : 
                        (N208)? mem[4347] : 
                        (N210)? mem[4427] : 
                        (N212)? mem[4507] : 
                        (N214)? mem[4587] : 
                        (N216)? mem[4667] : 
                        (N218)? mem[4747] : 
                        (N220)? mem[4827] : 
                        (N222)? mem[4907] : 
                        (N224)? mem[4987] : 
                        (N226)? mem[5067] : 1'b0;
  assign data_out[26] = (N163)? mem[26] : 
                        (N165)? mem[106] : 
                        (N167)? mem[186] : 
                        (N169)? mem[266] : 
                        (N171)? mem[346] : 
                        (N173)? mem[426] : 
                        (N175)? mem[506] : 
                        (N177)? mem[586] : 
                        (N179)? mem[666] : 
                        (N181)? mem[746] : 
                        (N183)? mem[826] : 
                        (N185)? mem[906] : 
                        (N187)? mem[986] : 
                        (N189)? mem[1066] : 
                        (N191)? mem[1146] : 
                        (N193)? mem[1226] : 
                        (N195)? mem[1306] : 
                        (N197)? mem[1386] : 
                        (N199)? mem[1466] : 
                        (N201)? mem[1546] : 
                        (N203)? mem[1626] : 
                        (N205)? mem[1706] : 
                        (N207)? mem[1786] : 
                        (N209)? mem[1866] : 
                        (N211)? mem[1946] : 
                        (N213)? mem[2026] : 
                        (N215)? mem[2106] : 
                        (N217)? mem[2186] : 
                        (N219)? mem[2266] : 
                        (N221)? mem[2346] : 
                        (N223)? mem[2426] : 
                        (N225)? mem[2506] : 
                        (N164)? mem[2586] : 
                        (N166)? mem[2666] : 
                        (N168)? mem[2746] : 
                        (N170)? mem[2826] : 
                        (N172)? mem[2906] : 
                        (N174)? mem[2986] : 
                        (N176)? mem[3066] : 
                        (N178)? mem[3146] : 
                        (N180)? mem[3226] : 
                        (N182)? mem[3306] : 
                        (N184)? mem[3386] : 
                        (N186)? mem[3466] : 
                        (N188)? mem[3546] : 
                        (N190)? mem[3626] : 
                        (N192)? mem[3706] : 
                        (N194)? mem[3786] : 
                        (N196)? mem[3866] : 
                        (N198)? mem[3946] : 
                        (N200)? mem[4026] : 
                        (N202)? mem[4106] : 
                        (N204)? mem[4186] : 
                        (N206)? mem[4266] : 
                        (N208)? mem[4346] : 
                        (N210)? mem[4426] : 
                        (N212)? mem[4506] : 
                        (N214)? mem[4586] : 
                        (N216)? mem[4666] : 
                        (N218)? mem[4746] : 
                        (N220)? mem[4826] : 
                        (N222)? mem[4906] : 
                        (N224)? mem[4986] : 
                        (N226)? mem[5066] : 1'b0;
  assign data_out[25] = (N163)? mem[25] : 
                        (N165)? mem[105] : 
                        (N167)? mem[185] : 
                        (N169)? mem[265] : 
                        (N171)? mem[345] : 
                        (N173)? mem[425] : 
                        (N175)? mem[505] : 
                        (N177)? mem[585] : 
                        (N179)? mem[665] : 
                        (N181)? mem[745] : 
                        (N183)? mem[825] : 
                        (N185)? mem[905] : 
                        (N187)? mem[985] : 
                        (N189)? mem[1065] : 
                        (N191)? mem[1145] : 
                        (N193)? mem[1225] : 
                        (N195)? mem[1305] : 
                        (N197)? mem[1385] : 
                        (N199)? mem[1465] : 
                        (N201)? mem[1545] : 
                        (N203)? mem[1625] : 
                        (N205)? mem[1705] : 
                        (N207)? mem[1785] : 
                        (N209)? mem[1865] : 
                        (N211)? mem[1945] : 
                        (N213)? mem[2025] : 
                        (N215)? mem[2105] : 
                        (N217)? mem[2185] : 
                        (N219)? mem[2265] : 
                        (N221)? mem[2345] : 
                        (N223)? mem[2425] : 
                        (N225)? mem[2505] : 
                        (N164)? mem[2585] : 
                        (N166)? mem[2665] : 
                        (N168)? mem[2745] : 
                        (N170)? mem[2825] : 
                        (N172)? mem[2905] : 
                        (N174)? mem[2985] : 
                        (N176)? mem[3065] : 
                        (N178)? mem[3145] : 
                        (N180)? mem[3225] : 
                        (N182)? mem[3305] : 
                        (N184)? mem[3385] : 
                        (N186)? mem[3465] : 
                        (N188)? mem[3545] : 
                        (N190)? mem[3625] : 
                        (N192)? mem[3705] : 
                        (N194)? mem[3785] : 
                        (N196)? mem[3865] : 
                        (N198)? mem[3945] : 
                        (N200)? mem[4025] : 
                        (N202)? mem[4105] : 
                        (N204)? mem[4185] : 
                        (N206)? mem[4265] : 
                        (N208)? mem[4345] : 
                        (N210)? mem[4425] : 
                        (N212)? mem[4505] : 
                        (N214)? mem[4585] : 
                        (N216)? mem[4665] : 
                        (N218)? mem[4745] : 
                        (N220)? mem[4825] : 
                        (N222)? mem[4905] : 
                        (N224)? mem[4985] : 
                        (N226)? mem[5065] : 1'b0;
  assign data_out[24] = (N163)? mem[24] : 
                        (N165)? mem[104] : 
                        (N167)? mem[184] : 
                        (N169)? mem[264] : 
                        (N171)? mem[344] : 
                        (N173)? mem[424] : 
                        (N175)? mem[504] : 
                        (N177)? mem[584] : 
                        (N179)? mem[664] : 
                        (N181)? mem[744] : 
                        (N183)? mem[824] : 
                        (N185)? mem[904] : 
                        (N187)? mem[984] : 
                        (N189)? mem[1064] : 
                        (N191)? mem[1144] : 
                        (N193)? mem[1224] : 
                        (N195)? mem[1304] : 
                        (N197)? mem[1384] : 
                        (N199)? mem[1464] : 
                        (N201)? mem[1544] : 
                        (N203)? mem[1624] : 
                        (N205)? mem[1704] : 
                        (N207)? mem[1784] : 
                        (N209)? mem[1864] : 
                        (N211)? mem[1944] : 
                        (N213)? mem[2024] : 
                        (N215)? mem[2104] : 
                        (N217)? mem[2184] : 
                        (N219)? mem[2264] : 
                        (N221)? mem[2344] : 
                        (N223)? mem[2424] : 
                        (N225)? mem[2504] : 
                        (N164)? mem[2584] : 
                        (N166)? mem[2664] : 
                        (N168)? mem[2744] : 
                        (N170)? mem[2824] : 
                        (N172)? mem[2904] : 
                        (N174)? mem[2984] : 
                        (N176)? mem[3064] : 
                        (N178)? mem[3144] : 
                        (N180)? mem[3224] : 
                        (N182)? mem[3304] : 
                        (N184)? mem[3384] : 
                        (N186)? mem[3464] : 
                        (N188)? mem[3544] : 
                        (N190)? mem[3624] : 
                        (N192)? mem[3704] : 
                        (N194)? mem[3784] : 
                        (N196)? mem[3864] : 
                        (N198)? mem[3944] : 
                        (N200)? mem[4024] : 
                        (N202)? mem[4104] : 
                        (N204)? mem[4184] : 
                        (N206)? mem[4264] : 
                        (N208)? mem[4344] : 
                        (N210)? mem[4424] : 
                        (N212)? mem[4504] : 
                        (N214)? mem[4584] : 
                        (N216)? mem[4664] : 
                        (N218)? mem[4744] : 
                        (N220)? mem[4824] : 
                        (N222)? mem[4904] : 
                        (N224)? mem[4984] : 
                        (N226)? mem[5064] : 1'b0;
  assign data_out[23] = (N163)? mem[23] : 
                        (N165)? mem[103] : 
                        (N167)? mem[183] : 
                        (N169)? mem[263] : 
                        (N171)? mem[343] : 
                        (N173)? mem[423] : 
                        (N175)? mem[503] : 
                        (N177)? mem[583] : 
                        (N179)? mem[663] : 
                        (N181)? mem[743] : 
                        (N183)? mem[823] : 
                        (N185)? mem[903] : 
                        (N187)? mem[983] : 
                        (N189)? mem[1063] : 
                        (N191)? mem[1143] : 
                        (N193)? mem[1223] : 
                        (N195)? mem[1303] : 
                        (N197)? mem[1383] : 
                        (N199)? mem[1463] : 
                        (N201)? mem[1543] : 
                        (N203)? mem[1623] : 
                        (N205)? mem[1703] : 
                        (N207)? mem[1783] : 
                        (N209)? mem[1863] : 
                        (N211)? mem[1943] : 
                        (N213)? mem[2023] : 
                        (N215)? mem[2103] : 
                        (N217)? mem[2183] : 
                        (N219)? mem[2263] : 
                        (N221)? mem[2343] : 
                        (N223)? mem[2423] : 
                        (N225)? mem[2503] : 
                        (N164)? mem[2583] : 
                        (N166)? mem[2663] : 
                        (N168)? mem[2743] : 
                        (N170)? mem[2823] : 
                        (N172)? mem[2903] : 
                        (N174)? mem[2983] : 
                        (N176)? mem[3063] : 
                        (N178)? mem[3143] : 
                        (N180)? mem[3223] : 
                        (N182)? mem[3303] : 
                        (N184)? mem[3383] : 
                        (N186)? mem[3463] : 
                        (N188)? mem[3543] : 
                        (N190)? mem[3623] : 
                        (N192)? mem[3703] : 
                        (N194)? mem[3783] : 
                        (N196)? mem[3863] : 
                        (N198)? mem[3943] : 
                        (N200)? mem[4023] : 
                        (N202)? mem[4103] : 
                        (N204)? mem[4183] : 
                        (N206)? mem[4263] : 
                        (N208)? mem[4343] : 
                        (N210)? mem[4423] : 
                        (N212)? mem[4503] : 
                        (N214)? mem[4583] : 
                        (N216)? mem[4663] : 
                        (N218)? mem[4743] : 
                        (N220)? mem[4823] : 
                        (N222)? mem[4903] : 
                        (N224)? mem[4983] : 
                        (N226)? mem[5063] : 1'b0;
  assign data_out[22] = (N163)? mem[22] : 
                        (N165)? mem[102] : 
                        (N167)? mem[182] : 
                        (N169)? mem[262] : 
                        (N171)? mem[342] : 
                        (N173)? mem[422] : 
                        (N175)? mem[502] : 
                        (N177)? mem[582] : 
                        (N179)? mem[662] : 
                        (N181)? mem[742] : 
                        (N183)? mem[822] : 
                        (N185)? mem[902] : 
                        (N187)? mem[982] : 
                        (N189)? mem[1062] : 
                        (N191)? mem[1142] : 
                        (N193)? mem[1222] : 
                        (N195)? mem[1302] : 
                        (N197)? mem[1382] : 
                        (N199)? mem[1462] : 
                        (N201)? mem[1542] : 
                        (N203)? mem[1622] : 
                        (N205)? mem[1702] : 
                        (N207)? mem[1782] : 
                        (N209)? mem[1862] : 
                        (N211)? mem[1942] : 
                        (N213)? mem[2022] : 
                        (N215)? mem[2102] : 
                        (N217)? mem[2182] : 
                        (N219)? mem[2262] : 
                        (N221)? mem[2342] : 
                        (N223)? mem[2422] : 
                        (N225)? mem[2502] : 
                        (N164)? mem[2582] : 
                        (N166)? mem[2662] : 
                        (N168)? mem[2742] : 
                        (N170)? mem[2822] : 
                        (N172)? mem[2902] : 
                        (N174)? mem[2982] : 
                        (N176)? mem[3062] : 
                        (N178)? mem[3142] : 
                        (N180)? mem[3222] : 
                        (N182)? mem[3302] : 
                        (N184)? mem[3382] : 
                        (N186)? mem[3462] : 
                        (N188)? mem[3542] : 
                        (N190)? mem[3622] : 
                        (N192)? mem[3702] : 
                        (N194)? mem[3782] : 
                        (N196)? mem[3862] : 
                        (N198)? mem[3942] : 
                        (N200)? mem[4022] : 
                        (N202)? mem[4102] : 
                        (N204)? mem[4182] : 
                        (N206)? mem[4262] : 
                        (N208)? mem[4342] : 
                        (N210)? mem[4422] : 
                        (N212)? mem[4502] : 
                        (N214)? mem[4582] : 
                        (N216)? mem[4662] : 
                        (N218)? mem[4742] : 
                        (N220)? mem[4822] : 
                        (N222)? mem[4902] : 
                        (N224)? mem[4982] : 
                        (N226)? mem[5062] : 1'b0;
  assign data_out[21] = (N163)? mem[21] : 
                        (N165)? mem[101] : 
                        (N167)? mem[181] : 
                        (N169)? mem[261] : 
                        (N171)? mem[341] : 
                        (N173)? mem[421] : 
                        (N175)? mem[501] : 
                        (N177)? mem[581] : 
                        (N179)? mem[661] : 
                        (N181)? mem[741] : 
                        (N183)? mem[821] : 
                        (N185)? mem[901] : 
                        (N187)? mem[981] : 
                        (N189)? mem[1061] : 
                        (N191)? mem[1141] : 
                        (N193)? mem[1221] : 
                        (N195)? mem[1301] : 
                        (N197)? mem[1381] : 
                        (N199)? mem[1461] : 
                        (N201)? mem[1541] : 
                        (N203)? mem[1621] : 
                        (N205)? mem[1701] : 
                        (N207)? mem[1781] : 
                        (N209)? mem[1861] : 
                        (N211)? mem[1941] : 
                        (N213)? mem[2021] : 
                        (N215)? mem[2101] : 
                        (N217)? mem[2181] : 
                        (N219)? mem[2261] : 
                        (N221)? mem[2341] : 
                        (N223)? mem[2421] : 
                        (N225)? mem[2501] : 
                        (N164)? mem[2581] : 
                        (N166)? mem[2661] : 
                        (N168)? mem[2741] : 
                        (N170)? mem[2821] : 
                        (N172)? mem[2901] : 
                        (N174)? mem[2981] : 
                        (N176)? mem[3061] : 
                        (N178)? mem[3141] : 
                        (N180)? mem[3221] : 
                        (N182)? mem[3301] : 
                        (N184)? mem[3381] : 
                        (N186)? mem[3461] : 
                        (N188)? mem[3541] : 
                        (N190)? mem[3621] : 
                        (N192)? mem[3701] : 
                        (N194)? mem[3781] : 
                        (N196)? mem[3861] : 
                        (N198)? mem[3941] : 
                        (N200)? mem[4021] : 
                        (N202)? mem[4101] : 
                        (N204)? mem[4181] : 
                        (N206)? mem[4261] : 
                        (N208)? mem[4341] : 
                        (N210)? mem[4421] : 
                        (N212)? mem[4501] : 
                        (N214)? mem[4581] : 
                        (N216)? mem[4661] : 
                        (N218)? mem[4741] : 
                        (N220)? mem[4821] : 
                        (N222)? mem[4901] : 
                        (N224)? mem[4981] : 
                        (N226)? mem[5061] : 1'b0;
  assign data_out[20] = (N163)? mem[20] : 
                        (N165)? mem[100] : 
                        (N167)? mem[180] : 
                        (N169)? mem[260] : 
                        (N171)? mem[340] : 
                        (N173)? mem[420] : 
                        (N175)? mem[500] : 
                        (N177)? mem[580] : 
                        (N179)? mem[660] : 
                        (N181)? mem[740] : 
                        (N183)? mem[820] : 
                        (N185)? mem[900] : 
                        (N187)? mem[980] : 
                        (N189)? mem[1060] : 
                        (N191)? mem[1140] : 
                        (N193)? mem[1220] : 
                        (N195)? mem[1300] : 
                        (N197)? mem[1380] : 
                        (N199)? mem[1460] : 
                        (N201)? mem[1540] : 
                        (N203)? mem[1620] : 
                        (N205)? mem[1700] : 
                        (N207)? mem[1780] : 
                        (N209)? mem[1860] : 
                        (N211)? mem[1940] : 
                        (N213)? mem[2020] : 
                        (N215)? mem[2100] : 
                        (N217)? mem[2180] : 
                        (N219)? mem[2260] : 
                        (N221)? mem[2340] : 
                        (N223)? mem[2420] : 
                        (N225)? mem[2500] : 
                        (N164)? mem[2580] : 
                        (N166)? mem[2660] : 
                        (N168)? mem[2740] : 
                        (N170)? mem[2820] : 
                        (N172)? mem[2900] : 
                        (N174)? mem[2980] : 
                        (N176)? mem[3060] : 
                        (N178)? mem[3140] : 
                        (N180)? mem[3220] : 
                        (N182)? mem[3300] : 
                        (N184)? mem[3380] : 
                        (N186)? mem[3460] : 
                        (N188)? mem[3540] : 
                        (N190)? mem[3620] : 
                        (N192)? mem[3700] : 
                        (N194)? mem[3780] : 
                        (N196)? mem[3860] : 
                        (N198)? mem[3940] : 
                        (N200)? mem[4020] : 
                        (N202)? mem[4100] : 
                        (N204)? mem[4180] : 
                        (N206)? mem[4260] : 
                        (N208)? mem[4340] : 
                        (N210)? mem[4420] : 
                        (N212)? mem[4500] : 
                        (N214)? mem[4580] : 
                        (N216)? mem[4660] : 
                        (N218)? mem[4740] : 
                        (N220)? mem[4820] : 
                        (N222)? mem[4900] : 
                        (N224)? mem[4980] : 
                        (N226)? mem[5060] : 1'b0;
  assign data_out[19] = (N163)? mem[19] : 
                        (N165)? mem[99] : 
                        (N167)? mem[179] : 
                        (N169)? mem[259] : 
                        (N171)? mem[339] : 
                        (N173)? mem[419] : 
                        (N175)? mem[499] : 
                        (N177)? mem[579] : 
                        (N179)? mem[659] : 
                        (N181)? mem[739] : 
                        (N183)? mem[819] : 
                        (N185)? mem[899] : 
                        (N187)? mem[979] : 
                        (N189)? mem[1059] : 
                        (N191)? mem[1139] : 
                        (N193)? mem[1219] : 
                        (N195)? mem[1299] : 
                        (N197)? mem[1379] : 
                        (N199)? mem[1459] : 
                        (N201)? mem[1539] : 
                        (N203)? mem[1619] : 
                        (N205)? mem[1699] : 
                        (N207)? mem[1779] : 
                        (N209)? mem[1859] : 
                        (N211)? mem[1939] : 
                        (N213)? mem[2019] : 
                        (N215)? mem[2099] : 
                        (N217)? mem[2179] : 
                        (N219)? mem[2259] : 
                        (N221)? mem[2339] : 
                        (N223)? mem[2419] : 
                        (N225)? mem[2499] : 
                        (N164)? mem[2579] : 
                        (N166)? mem[2659] : 
                        (N168)? mem[2739] : 
                        (N170)? mem[2819] : 
                        (N172)? mem[2899] : 
                        (N174)? mem[2979] : 
                        (N176)? mem[3059] : 
                        (N178)? mem[3139] : 
                        (N180)? mem[3219] : 
                        (N182)? mem[3299] : 
                        (N184)? mem[3379] : 
                        (N186)? mem[3459] : 
                        (N188)? mem[3539] : 
                        (N190)? mem[3619] : 
                        (N192)? mem[3699] : 
                        (N194)? mem[3779] : 
                        (N196)? mem[3859] : 
                        (N198)? mem[3939] : 
                        (N200)? mem[4019] : 
                        (N202)? mem[4099] : 
                        (N204)? mem[4179] : 
                        (N206)? mem[4259] : 
                        (N208)? mem[4339] : 
                        (N210)? mem[4419] : 
                        (N212)? mem[4499] : 
                        (N214)? mem[4579] : 
                        (N216)? mem[4659] : 
                        (N218)? mem[4739] : 
                        (N220)? mem[4819] : 
                        (N222)? mem[4899] : 
                        (N224)? mem[4979] : 
                        (N226)? mem[5059] : 1'b0;
  assign data_out[18] = (N163)? mem[18] : 
                        (N165)? mem[98] : 
                        (N167)? mem[178] : 
                        (N169)? mem[258] : 
                        (N171)? mem[338] : 
                        (N173)? mem[418] : 
                        (N175)? mem[498] : 
                        (N177)? mem[578] : 
                        (N179)? mem[658] : 
                        (N181)? mem[738] : 
                        (N183)? mem[818] : 
                        (N185)? mem[898] : 
                        (N187)? mem[978] : 
                        (N189)? mem[1058] : 
                        (N191)? mem[1138] : 
                        (N193)? mem[1218] : 
                        (N195)? mem[1298] : 
                        (N197)? mem[1378] : 
                        (N199)? mem[1458] : 
                        (N201)? mem[1538] : 
                        (N203)? mem[1618] : 
                        (N205)? mem[1698] : 
                        (N207)? mem[1778] : 
                        (N209)? mem[1858] : 
                        (N211)? mem[1938] : 
                        (N213)? mem[2018] : 
                        (N215)? mem[2098] : 
                        (N217)? mem[2178] : 
                        (N219)? mem[2258] : 
                        (N221)? mem[2338] : 
                        (N223)? mem[2418] : 
                        (N225)? mem[2498] : 
                        (N164)? mem[2578] : 
                        (N166)? mem[2658] : 
                        (N168)? mem[2738] : 
                        (N170)? mem[2818] : 
                        (N172)? mem[2898] : 
                        (N174)? mem[2978] : 
                        (N176)? mem[3058] : 
                        (N178)? mem[3138] : 
                        (N180)? mem[3218] : 
                        (N182)? mem[3298] : 
                        (N184)? mem[3378] : 
                        (N186)? mem[3458] : 
                        (N188)? mem[3538] : 
                        (N190)? mem[3618] : 
                        (N192)? mem[3698] : 
                        (N194)? mem[3778] : 
                        (N196)? mem[3858] : 
                        (N198)? mem[3938] : 
                        (N200)? mem[4018] : 
                        (N202)? mem[4098] : 
                        (N204)? mem[4178] : 
                        (N206)? mem[4258] : 
                        (N208)? mem[4338] : 
                        (N210)? mem[4418] : 
                        (N212)? mem[4498] : 
                        (N214)? mem[4578] : 
                        (N216)? mem[4658] : 
                        (N218)? mem[4738] : 
                        (N220)? mem[4818] : 
                        (N222)? mem[4898] : 
                        (N224)? mem[4978] : 
                        (N226)? mem[5058] : 1'b0;
  assign data_out[17] = (N163)? mem[17] : 
                        (N165)? mem[97] : 
                        (N167)? mem[177] : 
                        (N169)? mem[257] : 
                        (N171)? mem[337] : 
                        (N173)? mem[417] : 
                        (N175)? mem[497] : 
                        (N177)? mem[577] : 
                        (N179)? mem[657] : 
                        (N181)? mem[737] : 
                        (N183)? mem[817] : 
                        (N185)? mem[897] : 
                        (N187)? mem[977] : 
                        (N189)? mem[1057] : 
                        (N191)? mem[1137] : 
                        (N193)? mem[1217] : 
                        (N195)? mem[1297] : 
                        (N197)? mem[1377] : 
                        (N199)? mem[1457] : 
                        (N201)? mem[1537] : 
                        (N203)? mem[1617] : 
                        (N205)? mem[1697] : 
                        (N207)? mem[1777] : 
                        (N209)? mem[1857] : 
                        (N211)? mem[1937] : 
                        (N213)? mem[2017] : 
                        (N215)? mem[2097] : 
                        (N217)? mem[2177] : 
                        (N219)? mem[2257] : 
                        (N221)? mem[2337] : 
                        (N223)? mem[2417] : 
                        (N225)? mem[2497] : 
                        (N164)? mem[2577] : 
                        (N166)? mem[2657] : 
                        (N168)? mem[2737] : 
                        (N170)? mem[2817] : 
                        (N172)? mem[2897] : 
                        (N174)? mem[2977] : 
                        (N176)? mem[3057] : 
                        (N178)? mem[3137] : 
                        (N180)? mem[3217] : 
                        (N182)? mem[3297] : 
                        (N184)? mem[3377] : 
                        (N186)? mem[3457] : 
                        (N188)? mem[3537] : 
                        (N190)? mem[3617] : 
                        (N192)? mem[3697] : 
                        (N194)? mem[3777] : 
                        (N196)? mem[3857] : 
                        (N198)? mem[3937] : 
                        (N200)? mem[4017] : 
                        (N202)? mem[4097] : 
                        (N204)? mem[4177] : 
                        (N206)? mem[4257] : 
                        (N208)? mem[4337] : 
                        (N210)? mem[4417] : 
                        (N212)? mem[4497] : 
                        (N214)? mem[4577] : 
                        (N216)? mem[4657] : 
                        (N218)? mem[4737] : 
                        (N220)? mem[4817] : 
                        (N222)? mem[4897] : 
                        (N224)? mem[4977] : 
                        (N226)? mem[5057] : 1'b0;
  assign data_out[16] = (N163)? mem[16] : 
                        (N165)? mem[96] : 
                        (N167)? mem[176] : 
                        (N169)? mem[256] : 
                        (N171)? mem[336] : 
                        (N173)? mem[416] : 
                        (N175)? mem[496] : 
                        (N177)? mem[576] : 
                        (N179)? mem[656] : 
                        (N181)? mem[736] : 
                        (N183)? mem[816] : 
                        (N185)? mem[896] : 
                        (N187)? mem[976] : 
                        (N189)? mem[1056] : 
                        (N191)? mem[1136] : 
                        (N193)? mem[1216] : 
                        (N195)? mem[1296] : 
                        (N197)? mem[1376] : 
                        (N199)? mem[1456] : 
                        (N201)? mem[1536] : 
                        (N203)? mem[1616] : 
                        (N205)? mem[1696] : 
                        (N207)? mem[1776] : 
                        (N209)? mem[1856] : 
                        (N211)? mem[1936] : 
                        (N213)? mem[2016] : 
                        (N215)? mem[2096] : 
                        (N217)? mem[2176] : 
                        (N219)? mem[2256] : 
                        (N221)? mem[2336] : 
                        (N223)? mem[2416] : 
                        (N225)? mem[2496] : 
                        (N164)? mem[2576] : 
                        (N166)? mem[2656] : 
                        (N168)? mem[2736] : 
                        (N170)? mem[2816] : 
                        (N172)? mem[2896] : 
                        (N174)? mem[2976] : 
                        (N176)? mem[3056] : 
                        (N178)? mem[3136] : 
                        (N180)? mem[3216] : 
                        (N182)? mem[3296] : 
                        (N184)? mem[3376] : 
                        (N186)? mem[3456] : 
                        (N188)? mem[3536] : 
                        (N190)? mem[3616] : 
                        (N192)? mem[3696] : 
                        (N194)? mem[3776] : 
                        (N196)? mem[3856] : 
                        (N198)? mem[3936] : 
                        (N200)? mem[4016] : 
                        (N202)? mem[4096] : 
                        (N204)? mem[4176] : 
                        (N206)? mem[4256] : 
                        (N208)? mem[4336] : 
                        (N210)? mem[4416] : 
                        (N212)? mem[4496] : 
                        (N214)? mem[4576] : 
                        (N216)? mem[4656] : 
                        (N218)? mem[4736] : 
                        (N220)? mem[4816] : 
                        (N222)? mem[4896] : 
                        (N224)? mem[4976] : 
                        (N226)? mem[5056] : 1'b0;
  assign data_out[15] = (N163)? mem[15] : 
                        (N165)? mem[95] : 
                        (N167)? mem[175] : 
                        (N169)? mem[255] : 
                        (N171)? mem[335] : 
                        (N173)? mem[415] : 
                        (N175)? mem[495] : 
                        (N177)? mem[575] : 
                        (N179)? mem[655] : 
                        (N181)? mem[735] : 
                        (N183)? mem[815] : 
                        (N185)? mem[895] : 
                        (N187)? mem[975] : 
                        (N189)? mem[1055] : 
                        (N191)? mem[1135] : 
                        (N193)? mem[1215] : 
                        (N195)? mem[1295] : 
                        (N197)? mem[1375] : 
                        (N199)? mem[1455] : 
                        (N201)? mem[1535] : 
                        (N203)? mem[1615] : 
                        (N205)? mem[1695] : 
                        (N207)? mem[1775] : 
                        (N209)? mem[1855] : 
                        (N211)? mem[1935] : 
                        (N213)? mem[2015] : 
                        (N215)? mem[2095] : 
                        (N217)? mem[2175] : 
                        (N219)? mem[2255] : 
                        (N221)? mem[2335] : 
                        (N223)? mem[2415] : 
                        (N225)? mem[2495] : 
                        (N164)? mem[2575] : 
                        (N166)? mem[2655] : 
                        (N168)? mem[2735] : 
                        (N170)? mem[2815] : 
                        (N172)? mem[2895] : 
                        (N174)? mem[2975] : 
                        (N176)? mem[3055] : 
                        (N178)? mem[3135] : 
                        (N180)? mem[3215] : 
                        (N182)? mem[3295] : 
                        (N184)? mem[3375] : 
                        (N186)? mem[3455] : 
                        (N188)? mem[3535] : 
                        (N190)? mem[3615] : 
                        (N192)? mem[3695] : 
                        (N194)? mem[3775] : 
                        (N196)? mem[3855] : 
                        (N198)? mem[3935] : 
                        (N200)? mem[4015] : 
                        (N202)? mem[4095] : 
                        (N204)? mem[4175] : 
                        (N206)? mem[4255] : 
                        (N208)? mem[4335] : 
                        (N210)? mem[4415] : 
                        (N212)? mem[4495] : 
                        (N214)? mem[4575] : 
                        (N216)? mem[4655] : 
                        (N218)? mem[4735] : 
                        (N220)? mem[4815] : 
                        (N222)? mem[4895] : 
                        (N224)? mem[4975] : 
                        (N226)? mem[5055] : 1'b0;
  assign data_out[14] = (N163)? mem[14] : 
                        (N165)? mem[94] : 
                        (N167)? mem[174] : 
                        (N169)? mem[254] : 
                        (N171)? mem[334] : 
                        (N173)? mem[414] : 
                        (N175)? mem[494] : 
                        (N177)? mem[574] : 
                        (N179)? mem[654] : 
                        (N181)? mem[734] : 
                        (N183)? mem[814] : 
                        (N185)? mem[894] : 
                        (N187)? mem[974] : 
                        (N189)? mem[1054] : 
                        (N191)? mem[1134] : 
                        (N193)? mem[1214] : 
                        (N195)? mem[1294] : 
                        (N197)? mem[1374] : 
                        (N199)? mem[1454] : 
                        (N201)? mem[1534] : 
                        (N203)? mem[1614] : 
                        (N205)? mem[1694] : 
                        (N207)? mem[1774] : 
                        (N209)? mem[1854] : 
                        (N211)? mem[1934] : 
                        (N213)? mem[2014] : 
                        (N215)? mem[2094] : 
                        (N217)? mem[2174] : 
                        (N219)? mem[2254] : 
                        (N221)? mem[2334] : 
                        (N223)? mem[2414] : 
                        (N225)? mem[2494] : 
                        (N164)? mem[2574] : 
                        (N166)? mem[2654] : 
                        (N168)? mem[2734] : 
                        (N170)? mem[2814] : 
                        (N172)? mem[2894] : 
                        (N174)? mem[2974] : 
                        (N176)? mem[3054] : 
                        (N178)? mem[3134] : 
                        (N180)? mem[3214] : 
                        (N182)? mem[3294] : 
                        (N184)? mem[3374] : 
                        (N186)? mem[3454] : 
                        (N188)? mem[3534] : 
                        (N190)? mem[3614] : 
                        (N192)? mem[3694] : 
                        (N194)? mem[3774] : 
                        (N196)? mem[3854] : 
                        (N198)? mem[3934] : 
                        (N200)? mem[4014] : 
                        (N202)? mem[4094] : 
                        (N204)? mem[4174] : 
                        (N206)? mem[4254] : 
                        (N208)? mem[4334] : 
                        (N210)? mem[4414] : 
                        (N212)? mem[4494] : 
                        (N214)? mem[4574] : 
                        (N216)? mem[4654] : 
                        (N218)? mem[4734] : 
                        (N220)? mem[4814] : 
                        (N222)? mem[4894] : 
                        (N224)? mem[4974] : 
                        (N226)? mem[5054] : 1'b0;
  assign data_out[13] = (N163)? mem[13] : 
                        (N165)? mem[93] : 
                        (N167)? mem[173] : 
                        (N169)? mem[253] : 
                        (N171)? mem[333] : 
                        (N173)? mem[413] : 
                        (N175)? mem[493] : 
                        (N177)? mem[573] : 
                        (N179)? mem[653] : 
                        (N181)? mem[733] : 
                        (N183)? mem[813] : 
                        (N185)? mem[893] : 
                        (N187)? mem[973] : 
                        (N189)? mem[1053] : 
                        (N191)? mem[1133] : 
                        (N193)? mem[1213] : 
                        (N195)? mem[1293] : 
                        (N197)? mem[1373] : 
                        (N199)? mem[1453] : 
                        (N201)? mem[1533] : 
                        (N203)? mem[1613] : 
                        (N205)? mem[1693] : 
                        (N207)? mem[1773] : 
                        (N209)? mem[1853] : 
                        (N211)? mem[1933] : 
                        (N213)? mem[2013] : 
                        (N215)? mem[2093] : 
                        (N217)? mem[2173] : 
                        (N219)? mem[2253] : 
                        (N221)? mem[2333] : 
                        (N223)? mem[2413] : 
                        (N225)? mem[2493] : 
                        (N164)? mem[2573] : 
                        (N166)? mem[2653] : 
                        (N168)? mem[2733] : 
                        (N170)? mem[2813] : 
                        (N172)? mem[2893] : 
                        (N174)? mem[2973] : 
                        (N176)? mem[3053] : 
                        (N178)? mem[3133] : 
                        (N180)? mem[3213] : 
                        (N182)? mem[3293] : 
                        (N184)? mem[3373] : 
                        (N186)? mem[3453] : 
                        (N188)? mem[3533] : 
                        (N190)? mem[3613] : 
                        (N192)? mem[3693] : 
                        (N194)? mem[3773] : 
                        (N196)? mem[3853] : 
                        (N198)? mem[3933] : 
                        (N200)? mem[4013] : 
                        (N202)? mem[4093] : 
                        (N204)? mem[4173] : 
                        (N206)? mem[4253] : 
                        (N208)? mem[4333] : 
                        (N210)? mem[4413] : 
                        (N212)? mem[4493] : 
                        (N214)? mem[4573] : 
                        (N216)? mem[4653] : 
                        (N218)? mem[4733] : 
                        (N220)? mem[4813] : 
                        (N222)? mem[4893] : 
                        (N224)? mem[4973] : 
                        (N226)? mem[5053] : 1'b0;
  assign data_out[12] = (N163)? mem[12] : 
                        (N165)? mem[92] : 
                        (N167)? mem[172] : 
                        (N169)? mem[252] : 
                        (N171)? mem[332] : 
                        (N173)? mem[412] : 
                        (N175)? mem[492] : 
                        (N177)? mem[572] : 
                        (N179)? mem[652] : 
                        (N181)? mem[732] : 
                        (N183)? mem[812] : 
                        (N185)? mem[892] : 
                        (N187)? mem[972] : 
                        (N189)? mem[1052] : 
                        (N191)? mem[1132] : 
                        (N193)? mem[1212] : 
                        (N195)? mem[1292] : 
                        (N197)? mem[1372] : 
                        (N199)? mem[1452] : 
                        (N201)? mem[1532] : 
                        (N203)? mem[1612] : 
                        (N205)? mem[1692] : 
                        (N207)? mem[1772] : 
                        (N209)? mem[1852] : 
                        (N211)? mem[1932] : 
                        (N213)? mem[2012] : 
                        (N215)? mem[2092] : 
                        (N217)? mem[2172] : 
                        (N219)? mem[2252] : 
                        (N221)? mem[2332] : 
                        (N223)? mem[2412] : 
                        (N225)? mem[2492] : 
                        (N164)? mem[2572] : 
                        (N166)? mem[2652] : 
                        (N168)? mem[2732] : 
                        (N170)? mem[2812] : 
                        (N172)? mem[2892] : 
                        (N174)? mem[2972] : 
                        (N176)? mem[3052] : 
                        (N178)? mem[3132] : 
                        (N180)? mem[3212] : 
                        (N182)? mem[3292] : 
                        (N184)? mem[3372] : 
                        (N186)? mem[3452] : 
                        (N188)? mem[3532] : 
                        (N190)? mem[3612] : 
                        (N192)? mem[3692] : 
                        (N194)? mem[3772] : 
                        (N196)? mem[3852] : 
                        (N198)? mem[3932] : 
                        (N200)? mem[4012] : 
                        (N202)? mem[4092] : 
                        (N204)? mem[4172] : 
                        (N206)? mem[4252] : 
                        (N208)? mem[4332] : 
                        (N210)? mem[4412] : 
                        (N212)? mem[4492] : 
                        (N214)? mem[4572] : 
                        (N216)? mem[4652] : 
                        (N218)? mem[4732] : 
                        (N220)? mem[4812] : 
                        (N222)? mem[4892] : 
                        (N224)? mem[4972] : 
                        (N226)? mem[5052] : 1'b0;
  assign data_out[11] = (N163)? mem[11] : 
                        (N165)? mem[91] : 
                        (N167)? mem[171] : 
                        (N169)? mem[251] : 
                        (N171)? mem[331] : 
                        (N173)? mem[411] : 
                        (N175)? mem[491] : 
                        (N177)? mem[571] : 
                        (N179)? mem[651] : 
                        (N181)? mem[731] : 
                        (N183)? mem[811] : 
                        (N185)? mem[891] : 
                        (N187)? mem[971] : 
                        (N189)? mem[1051] : 
                        (N191)? mem[1131] : 
                        (N193)? mem[1211] : 
                        (N195)? mem[1291] : 
                        (N197)? mem[1371] : 
                        (N199)? mem[1451] : 
                        (N201)? mem[1531] : 
                        (N203)? mem[1611] : 
                        (N205)? mem[1691] : 
                        (N207)? mem[1771] : 
                        (N209)? mem[1851] : 
                        (N211)? mem[1931] : 
                        (N213)? mem[2011] : 
                        (N215)? mem[2091] : 
                        (N217)? mem[2171] : 
                        (N219)? mem[2251] : 
                        (N221)? mem[2331] : 
                        (N223)? mem[2411] : 
                        (N225)? mem[2491] : 
                        (N164)? mem[2571] : 
                        (N166)? mem[2651] : 
                        (N168)? mem[2731] : 
                        (N170)? mem[2811] : 
                        (N172)? mem[2891] : 
                        (N174)? mem[2971] : 
                        (N176)? mem[3051] : 
                        (N178)? mem[3131] : 
                        (N180)? mem[3211] : 
                        (N182)? mem[3291] : 
                        (N184)? mem[3371] : 
                        (N186)? mem[3451] : 
                        (N188)? mem[3531] : 
                        (N190)? mem[3611] : 
                        (N192)? mem[3691] : 
                        (N194)? mem[3771] : 
                        (N196)? mem[3851] : 
                        (N198)? mem[3931] : 
                        (N200)? mem[4011] : 
                        (N202)? mem[4091] : 
                        (N204)? mem[4171] : 
                        (N206)? mem[4251] : 
                        (N208)? mem[4331] : 
                        (N210)? mem[4411] : 
                        (N212)? mem[4491] : 
                        (N214)? mem[4571] : 
                        (N216)? mem[4651] : 
                        (N218)? mem[4731] : 
                        (N220)? mem[4811] : 
                        (N222)? mem[4891] : 
                        (N224)? mem[4971] : 
                        (N226)? mem[5051] : 1'b0;
  assign data_out[10] = (N163)? mem[10] : 
                        (N165)? mem[90] : 
                        (N167)? mem[170] : 
                        (N169)? mem[250] : 
                        (N171)? mem[330] : 
                        (N173)? mem[410] : 
                        (N175)? mem[490] : 
                        (N177)? mem[570] : 
                        (N179)? mem[650] : 
                        (N181)? mem[730] : 
                        (N183)? mem[810] : 
                        (N185)? mem[890] : 
                        (N187)? mem[970] : 
                        (N189)? mem[1050] : 
                        (N191)? mem[1130] : 
                        (N193)? mem[1210] : 
                        (N195)? mem[1290] : 
                        (N197)? mem[1370] : 
                        (N199)? mem[1450] : 
                        (N201)? mem[1530] : 
                        (N203)? mem[1610] : 
                        (N205)? mem[1690] : 
                        (N207)? mem[1770] : 
                        (N209)? mem[1850] : 
                        (N211)? mem[1930] : 
                        (N213)? mem[2010] : 
                        (N215)? mem[2090] : 
                        (N217)? mem[2170] : 
                        (N219)? mem[2250] : 
                        (N221)? mem[2330] : 
                        (N223)? mem[2410] : 
                        (N225)? mem[2490] : 
                        (N164)? mem[2570] : 
                        (N166)? mem[2650] : 
                        (N168)? mem[2730] : 
                        (N170)? mem[2810] : 
                        (N172)? mem[2890] : 
                        (N174)? mem[2970] : 
                        (N176)? mem[3050] : 
                        (N178)? mem[3130] : 
                        (N180)? mem[3210] : 
                        (N182)? mem[3290] : 
                        (N184)? mem[3370] : 
                        (N186)? mem[3450] : 
                        (N188)? mem[3530] : 
                        (N190)? mem[3610] : 
                        (N192)? mem[3690] : 
                        (N194)? mem[3770] : 
                        (N196)? mem[3850] : 
                        (N198)? mem[3930] : 
                        (N200)? mem[4010] : 
                        (N202)? mem[4090] : 
                        (N204)? mem[4170] : 
                        (N206)? mem[4250] : 
                        (N208)? mem[4330] : 
                        (N210)? mem[4410] : 
                        (N212)? mem[4490] : 
                        (N214)? mem[4570] : 
                        (N216)? mem[4650] : 
                        (N218)? mem[4730] : 
                        (N220)? mem[4810] : 
                        (N222)? mem[4890] : 
                        (N224)? mem[4970] : 
                        (N226)? mem[5050] : 1'b0;
  assign data_out[9] = (N163)? mem[9] : 
                       (N165)? mem[89] : 
                       (N167)? mem[169] : 
                       (N169)? mem[249] : 
                       (N171)? mem[329] : 
                       (N173)? mem[409] : 
                       (N175)? mem[489] : 
                       (N177)? mem[569] : 
                       (N179)? mem[649] : 
                       (N181)? mem[729] : 
                       (N183)? mem[809] : 
                       (N185)? mem[889] : 
                       (N187)? mem[969] : 
                       (N189)? mem[1049] : 
                       (N191)? mem[1129] : 
                       (N193)? mem[1209] : 
                       (N195)? mem[1289] : 
                       (N197)? mem[1369] : 
                       (N199)? mem[1449] : 
                       (N201)? mem[1529] : 
                       (N203)? mem[1609] : 
                       (N205)? mem[1689] : 
                       (N207)? mem[1769] : 
                       (N209)? mem[1849] : 
                       (N211)? mem[1929] : 
                       (N213)? mem[2009] : 
                       (N215)? mem[2089] : 
                       (N217)? mem[2169] : 
                       (N219)? mem[2249] : 
                       (N221)? mem[2329] : 
                       (N223)? mem[2409] : 
                       (N225)? mem[2489] : 
                       (N164)? mem[2569] : 
                       (N166)? mem[2649] : 
                       (N168)? mem[2729] : 
                       (N170)? mem[2809] : 
                       (N172)? mem[2889] : 
                       (N174)? mem[2969] : 
                       (N176)? mem[3049] : 
                       (N178)? mem[3129] : 
                       (N180)? mem[3209] : 
                       (N182)? mem[3289] : 
                       (N184)? mem[3369] : 
                       (N186)? mem[3449] : 
                       (N188)? mem[3529] : 
                       (N190)? mem[3609] : 
                       (N192)? mem[3689] : 
                       (N194)? mem[3769] : 
                       (N196)? mem[3849] : 
                       (N198)? mem[3929] : 
                       (N200)? mem[4009] : 
                       (N202)? mem[4089] : 
                       (N204)? mem[4169] : 
                       (N206)? mem[4249] : 
                       (N208)? mem[4329] : 
                       (N210)? mem[4409] : 
                       (N212)? mem[4489] : 
                       (N214)? mem[4569] : 
                       (N216)? mem[4649] : 
                       (N218)? mem[4729] : 
                       (N220)? mem[4809] : 
                       (N222)? mem[4889] : 
                       (N224)? mem[4969] : 
                       (N226)? mem[5049] : 1'b0;
  assign data_out[8] = (N163)? mem[8] : 
                       (N165)? mem[88] : 
                       (N167)? mem[168] : 
                       (N169)? mem[248] : 
                       (N171)? mem[328] : 
                       (N173)? mem[408] : 
                       (N175)? mem[488] : 
                       (N177)? mem[568] : 
                       (N179)? mem[648] : 
                       (N181)? mem[728] : 
                       (N183)? mem[808] : 
                       (N185)? mem[888] : 
                       (N187)? mem[968] : 
                       (N189)? mem[1048] : 
                       (N191)? mem[1128] : 
                       (N193)? mem[1208] : 
                       (N195)? mem[1288] : 
                       (N197)? mem[1368] : 
                       (N199)? mem[1448] : 
                       (N201)? mem[1528] : 
                       (N203)? mem[1608] : 
                       (N205)? mem[1688] : 
                       (N207)? mem[1768] : 
                       (N209)? mem[1848] : 
                       (N211)? mem[1928] : 
                       (N213)? mem[2008] : 
                       (N215)? mem[2088] : 
                       (N217)? mem[2168] : 
                       (N219)? mem[2248] : 
                       (N221)? mem[2328] : 
                       (N223)? mem[2408] : 
                       (N225)? mem[2488] : 
                       (N164)? mem[2568] : 
                       (N166)? mem[2648] : 
                       (N168)? mem[2728] : 
                       (N170)? mem[2808] : 
                       (N172)? mem[2888] : 
                       (N174)? mem[2968] : 
                       (N176)? mem[3048] : 
                       (N178)? mem[3128] : 
                       (N180)? mem[3208] : 
                       (N182)? mem[3288] : 
                       (N184)? mem[3368] : 
                       (N186)? mem[3448] : 
                       (N188)? mem[3528] : 
                       (N190)? mem[3608] : 
                       (N192)? mem[3688] : 
                       (N194)? mem[3768] : 
                       (N196)? mem[3848] : 
                       (N198)? mem[3928] : 
                       (N200)? mem[4008] : 
                       (N202)? mem[4088] : 
                       (N204)? mem[4168] : 
                       (N206)? mem[4248] : 
                       (N208)? mem[4328] : 
                       (N210)? mem[4408] : 
                       (N212)? mem[4488] : 
                       (N214)? mem[4568] : 
                       (N216)? mem[4648] : 
                       (N218)? mem[4728] : 
                       (N220)? mem[4808] : 
                       (N222)? mem[4888] : 
                       (N224)? mem[4968] : 
                       (N226)? mem[5048] : 1'b0;
  assign data_out[7] = (N163)? mem[7] : 
                       (N165)? mem[87] : 
                       (N167)? mem[167] : 
                       (N169)? mem[247] : 
                       (N171)? mem[327] : 
                       (N173)? mem[407] : 
                       (N175)? mem[487] : 
                       (N177)? mem[567] : 
                       (N179)? mem[647] : 
                       (N181)? mem[727] : 
                       (N183)? mem[807] : 
                       (N185)? mem[887] : 
                       (N187)? mem[967] : 
                       (N189)? mem[1047] : 
                       (N191)? mem[1127] : 
                       (N193)? mem[1207] : 
                       (N195)? mem[1287] : 
                       (N197)? mem[1367] : 
                       (N199)? mem[1447] : 
                       (N201)? mem[1527] : 
                       (N203)? mem[1607] : 
                       (N205)? mem[1687] : 
                       (N207)? mem[1767] : 
                       (N209)? mem[1847] : 
                       (N211)? mem[1927] : 
                       (N213)? mem[2007] : 
                       (N215)? mem[2087] : 
                       (N217)? mem[2167] : 
                       (N219)? mem[2247] : 
                       (N221)? mem[2327] : 
                       (N223)? mem[2407] : 
                       (N225)? mem[2487] : 
                       (N164)? mem[2567] : 
                       (N166)? mem[2647] : 
                       (N168)? mem[2727] : 
                       (N170)? mem[2807] : 
                       (N172)? mem[2887] : 
                       (N174)? mem[2967] : 
                       (N176)? mem[3047] : 
                       (N178)? mem[3127] : 
                       (N180)? mem[3207] : 
                       (N182)? mem[3287] : 
                       (N184)? mem[3367] : 
                       (N186)? mem[3447] : 
                       (N188)? mem[3527] : 
                       (N190)? mem[3607] : 
                       (N192)? mem[3687] : 
                       (N194)? mem[3767] : 
                       (N196)? mem[3847] : 
                       (N198)? mem[3927] : 
                       (N200)? mem[4007] : 
                       (N202)? mem[4087] : 
                       (N204)? mem[4167] : 
                       (N206)? mem[4247] : 
                       (N208)? mem[4327] : 
                       (N210)? mem[4407] : 
                       (N212)? mem[4487] : 
                       (N214)? mem[4567] : 
                       (N216)? mem[4647] : 
                       (N218)? mem[4727] : 
                       (N220)? mem[4807] : 
                       (N222)? mem[4887] : 
                       (N224)? mem[4967] : 
                       (N226)? mem[5047] : 1'b0;
  assign data_out[6] = (N163)? mem[6] : 
                       (N165)? mem[86] : 
                       (N167)? mem[166] : 
                       (N169)? mem[246] : 
                       (N171)? mem[326] : 
                       (N173)? mem[406] : 
                       (N175)? mem[486] : 
                       (N177)? mem[566] : 
                       (N179)? mem[646] : 
                       (N181)? mem[726] : 
                       (N183)? mem[806] : 
                       (N185)? mem[886] : 
                       (N187)? mem[966] : 
                       (N189)? mem[1046] : 
                       (N191)? mem[1126] : 
                       (N193)? mem[1206] : 
                       (N195)? mem[1286] : 
                       (N197)? mem[1366] : 
                       (N199)? mem[1446] : 
                       (N201)? mem[1526] : 
                       (N203)? mem[1606] : 
                       (N205)? mem[1686] : 
                       (N207)? mem[1766] : 
                       (N209)? mem[1846] : 
                       (N211)? mem[1926] : 
                       (N213)? mem[2006] : 
                       (N215)? mem[2086] : 
                       (N217)? mem[2166] : 
                       (N219)? mem[2246] : 
                       (N221)? mem[2326] : 
                       (N223)? mem[2406] : 
                       (N225)? mem[2486] : 
                       (N164)? mem[2566] : 
                       (N166)? mem[2646] : 
                       (N168)? mem[2726] : 
                       (N170)? mem[2806] : 
                       (N172)? mem[2886] : 
                       (N174)? mem[2966] : 
                       (N176)? mem[3046] : 
                       (N178)? mem[3126] : 
                       (N180)? mem[3206] : 
                       (N182)? mem[3286] : 
                       (N184)? mem[3366] : 
                       (N186)? mem[3446] : 
                       (N188)? mem[3526] : 
                       (N190)? mem[3606] : 
                       (N192)? mem[3686] : 
                       (N194)? mem[3766] : 
                       (N196)? mem[3846] : 
                       (N198)? mem[3926] : 
                       (N200)? mem[4006] : 
                       (N202)? mem[4086] : 
                       (N204)? mem[4166] : 
                       (N206)? mem[4246] : 
                       (N208)? mem[4326] : 
                       (N210)? mem[4406] : 
                       (N212)? mem[4486] : 
                       (N214)? mem[4566] : 
                       (N216)? mem[4646] : 
                       (N218)? mem[4726] : 
                       (N220)? mem[4806] : 
                       (N222)? mem[4886] : 
                       (N224)? mem[4966] : 
                       (N226)? mem[5046] : 1'b0;
  assign data_out[5] = (N163)? mem[5] : 
                       (N165)? mem[85] : 
                       (N167)? mem[165] : 
                       (N169)? mem[245] : 
                       (N171)? mem[325] : 
                       (N173)? mem[405] : 
                       (N175)? mem[485] : 
                       (N177)? mem[565] : 
                       (N179)? mem[645] : 
                       (N181)? mem[725] : 
                       (N183)? mem[805] : 
                       (N185)? mem[885] : 
                       (N187)? mem[965] : 
                       (N189)? mem[1045] : 
                       (N191)? mem[1125] : 
                       (N193)? mem[1205] : 
                       (N195)? mem[1285] : 
                       (N197)? mem[1365] : 
                       (N199)? mem[1445] : 
                       (N201)? mem[1525] : 
                       (N203)? mem[1605] : 
                       (N205)? mem[1685] : 
                       (N207)? mem[1765] : 
                       (N209)? mem[1845] : 
                       (N211)? mem[1925] : 
                       (N213)? mem[2005] : 
                       (N215)? mem[2085] : 
                       (N217)? mem[2165] : 
                       (N219)? mem[2245] : 
                       (N221)? mem[2325] : 
                       (N223)? mem[2405] : 
                       (N225)? mem[2485] : 
                       (N164)? mem[2565] : 
                       (N166)? mem[2645] : 
                       (N168)? mem[2725] : 
                       (N170)? mem[2805] : 
                       (N172)? mem[2885] : 
                       (N174)? mem[2965] : 
                       (N176)? mem[3045] : 
                       (N178)? mem[3125] : 
                       (N180)? mem[3205] : 
                       (N182)? mem[3285] : 
                       (N184)? mem[3365] : 
                       (N186)? mem[3445] : 
                       (N188)? mem[3525] : 
                       (N190)? mem[3605] : 
                       (N192)? mem[3685] : 
                       (N194)? mem[3765] : 
                       (N196)? mem[3845] : 
                       (N198)? mem[3925] : 
                       (N200)? mem[4005] : 
                       (N202)? mem[4085] : 
                       (N204)? mem[4165] : 
                       (N206)? mem[4245] : 
                       (N208)? mem[4325] : 
                       (N210)? mem[4405] : 
                       (N212)? mem[4485] : 
                       (N214)? mem[4565] : 
                       (N216)? mem[4645] : 
                       (N218)? mem[4725] : 
                       (N220)? mem[4805] : 
                       (N222)? mem[4885] : 
                       (N224)? mem[4965] : 
                       (N226)? mem[5045] : 1'b0;
  assign data_out[4] = (N163)? mem[4] : 
                       (N165)? mem[84] : 
                       (N167)? mem[164] : 
                       (N169)? mem[244] : 
                       (N171)? mem[324] : 
                       (N173)? mem[404] : 
                       (N175)? mem[484] : 
                       (N177)? mem[564] : 
                       (N179)? mem[644] : 
                       (N181)? mem[724] : 
                       (N183)? mem[804] : 
                       (N185)? mem[884] : 
                       (N187)? mem[964] : 
                       (N189)? mem[1044] : 
                       (N191)? mem[1124] : 
                       (N193)? mem[1204] : 
                       (N195)? mem[1284] : 
                       (N197)? mem[1364] : 
                       (N199)? mem[1444] : 
                       (N201)? mem[1524] : 
                       (N203)? mem[1604] : 
                       (N205)? mem[1684] : 
                       (N207)? mem[1764] : 
                       (N209)? mem[1844] : 
                       (N211)? mem[1924] : 
                       (N213)? mem[2004] : 
                       (N215)? mem[2084] : 
                       (N217)? mem[2164] : 
                       (N219)? mem[2244] : 
                       (N221)? mem[2324] : 
                       (N223)? mem[2404] : 
                       (N225)? mem[2484] : 
                       (N164)? mem[2564] : 
                       (N166)? mem[2644] : 
                       (N168)? mem[2724] : 
                       (N170)? mem[2804] : 
                       (N172)? mem[2884] : 
                       (N174)? mem[2964] : 
                       (N176)? mem[3044] : 
                       (N178)? mem[3124] : 
                       (N180)? mem[3204] : 
                       (N182)? mem[3284] : 
                       (N184)? mem[3364] : 
                       (N186)? mem[3444] : 
                       (N188)? mem[3524] : 
                       (N190)? mem[3604] : 
                       (N192)? mem[3684] : 
                       (N194)? mem[3764] : 
                       (N196)? mem[3844] : 
                       (N198)? mem[3924] : 
                       (N200)? mem[4004] : 
                       (N202)? mem[4084] : 
                       (N204)? mem[4164] : 
                       (N206)? mem[4244] : 
                       (N208)? mem[4324] : 
                       (N210)? mem[4404] : 
                       (N212)? mem[4484] : 
                       (N214)? mem[4564] : 
                       (N216)? mem[4644] : 
                       (N218)? mem[4724] : 
                       (N220)? mem[4804] : 
                       (N222)? mem[4884] : 
                       (N224)? mem[4964] : 
                       (N226)? mem[5044] : 1'b0;
  assign data_out[3] = (N163)? mem[3] : 
                       (N165)? mem[83] : 
                       (N167)? mem[163] : 
                       (N169)? mem[243] : 
                       (N171)? mem[323] : 
                       (N173)? mem[403] : 
                       (N175)? mem[483] : 
                       (N177)? mem[563] : 
                       (N179)? mem[643] : 
                       (N181)? mem[723] : 
                       (N183)? mem[803] : 
                       (N185)? mem[883] : 
                       (N187)? mem[963] : 
                       (N189)? mem[1043] : 
                       (N191)? mem[1123] : 
                       (N193)? mem[1203] : 
                       (N195)? mem[1283] : 
                       (N197)? mem[1363] : 
                       (N199)? mem[1443] : 
                       (N201)? mem[1523] : 
                       (N203)? mem[1603] : 
                       (N205)? mem[1683] : 
                       (N207)? mem[1763] : 
                       (N209)? mem[1843] : 
                       (N211)? mem[1923] : 
                       (N213)? mem[2003] : 
                       (N215)? mem[2083] : 
                       (N217)? mem[2163] : 
                       (N219)? mem[2243] : 
                       (N221)? mem[2323] : 
                       (N223)? mem[2403] : 
                       (N225)? mem[2483] : 
                       (N164)? mem[2563] : 
                       (N166)? mem[2643] : 
                       (N168)? mem[2723] : 
                       (N170)? mem[2803] : 
                       (N172)? mem[2883] : 
                       (N174)? mem[2963] : 
                       (N176)? mem[3043] : 
                       (N178)? mem[3123] : 
                       (N180)? mem[3203] : 
                       (N182)? mem[3283] : 
                       (N184)? mem[3363] : 
                       (N186)? mem[3443] : 
                       (N188)? mem[3523] : 
                       (N190)? mem[3603] : 
                       (N192)? mem[3683] : 
                       (N194)? mem[3763] : 
                       (N196)? mem[3843] : 
                       (N198)? mem[3923] : 
                       (N200)? mem[4003] : 
                       (N202)? mem[4083] : 
                       (N204)? mem[4163] : 
                       (N206)? mem[4243] : 
                       (N208)? mem[4323] : 
                       (N210)? mem[4403] : 
                       (N212)? mem[4483] : 
                       (N214)? mem[4563] : 
                       (N216)? mem[4643] : 
                       (N218)? mem[4723] : 
                       (N220)? mem[4803] : 
                       (N222)? mem[4883] : 
                       (N224)? mem[4963] : 
                       (N226)? mem[5043] : 1'b0;
  assign data_out[2] = (N163)? mem[2] : 
                       (N165)? mem[82] : 
                       (N167)? mem[162] : 
                       (N169)? mem[242] : 
                       (N171)? mem[322] : 
                       (N173)? mem[402] : 
                       (N175)? mem[482] : 
                       (N177)? mem[562] : 
                       (N179)? mem[642] : 
                       (N181)? mem[722] : 
                       (N183)? mem[802] : 
                       (N185)? mem[882] : 
                       (N187)? mem[962] : 
                       (N189)? mem[1042] : 
                       (N191)? mem[1122] : 
                       (N193)? mem[1202] : 
                       (N195)? mem[1282] : 
                       (N197)? mem[1362] : 
                       (N199)? mem[1442] : 
                       (N201)? mem[1522] : 
                       (N203)? mem[1602] : 
                       (N205)? mem[1682] : 
                       (N207)? mem[1762] : 
                       (N209)? mem[1842] : 
                       (N211)? mem[1922] : 
                       (N213)? mem[2002] : 
                       (N215)? mem[2082] : 
                       (N217)? mem[2162] : 
                       (N219)? mem[2242] : 
                       (N221)? mem[2322] : 
                       (N223)? mem[2402] : 
                       (N225)? mem[2482] : 
                       (N164)? mem[2562] : 
                       (N166)? mem[2642] : 
                       (N168)? mem[2722] : 
                       (N170)? mem[2802] : 
                       (N172)? mem[2882] : 
                       (N174)? mem[2962] : 
                       (N176)? mem[3042] : 
                       (N178)? mem[3122] : 
                       (N180)? mem[3202] : 
                       (N182)? mem[3282] : 
                       (N184)? mem[3362] : 
                       (N186)? mem[3442] : 
                       (N188)? mem[3522] : 
                       (N190)? mem[3602] : 
                       (N192)? mem[3682] : 
                       (N194)? mem[3762] : 
                       (N196)? mem[3842] : 
                       (N198)? mem[3922] : 
                       (N200)? mem[4002] : 
                       (N202)? mem[4082] : 
                       (N204)? mem[4162] : 
                       (N206)? mem[4242] : 
                       (N208)? mem[4322] : 
                       (N210)? mem[4402] : 
                       (N212)? mem[4482] : 
                       (N214)? mem[4562] : 
                       (N216)? mem[4642] : 
                       (N218)? mem[4722] : 
                       (N220)? mem[4802] : 
                       (N222)? mem[4882] : 
                       (N224)? mem[4962] : 
                       (N226)? mem[5042] : 1'b0;
  assign data_out[1] = (N163)? mem[1] : 
                       (N165)? mem[81] : 
                       (N167)? mem[161] : 
                       (N169)? mem[241] : 
                       (N171)? mem[321] : 
                       (N173)? mem[401] : 
                       (N175)? mem[481] : 
                       (N177)? mem[561] : 
                       (N179)? mem[641] : 
                       (N181)? mem[721] : 
                       (N183)? mem[801] : 
                       (N185)? mem[881] : 
                       (N187)? mem[961] : 
                       (N189)? mem[1041] : 
                       (N191)? mem[1121] : 
                       (N193)? mem[1201] : 
                       (N195)? mem[1281] : 
                       (N197)? mem[1361] : 
                       (N199)? mem[1441] : 
                       (N201)? mem[1521] : 
                       (N203)? mem[1601] : 
                       (N205)? mem[1681] : 
                       (N207)? mem[1761] : 
                       (N209)? mem[1841] : 
                       (N211)? mem[1921] : 
                       (N213)? mem[2001] : 
                       (N215)? mem[2081] : 
                       (N217)? mem[2161] : 
                       (N219)? mem[2241] : 
                       (N221)? mem[2321] : 
                       (N223)? mem[2401] : 
                       (N225)? mem[2481] : 
                       (N164)? mem[2561] : 
                       (N166)? mem[2641] : 
                       (N168)? mem[2721] : 
                       (N170)? mem[2801] : 
                       (N172)? mem[2881] : 
                       (N174)? mem[2961] : 
                       (N176)? mem[3041] : 
                       (N178)? mem[3121] : 
                       (N180)? mem[3201] : 
                       (N182)? mem[3281] : 
                       (N184)? mem[3361] : 
                       (N186)? mem[3441] : 
                       (N188)? mem[3521] : 
                       (N190)? mem[3601] : 
                       (N192)? mem[3681] : 
                       (N194)? mem[3761] : 
                       (N196)? mem[3841] : 
                       (N198)? mem[3921] : 
                       (N200)? mem[4001] : 
                       (N202)? mem[4081] : 
                       (N204)? mem[4161] : 
                       (N206)? mem[4241] : 
                       (N208)? mem[4321] : 
                       (N210)? mem[4401] : 
                       (N212)? mem[4481] : 
                       (N214)? mem[4561] : 
                       (N216)? mem[4641] : 
                       (N218)? mem[4721] : 
                       (N220)? mem[4801] : 
                       (N222)? mem[4881] : 
                       (N224)? mem[4961] : 
                       (N226)? mem[5041] : 1'b0;
  assign data_out[0] = (N163)? mem[0] : 
                       (N165)? mem[80] : 
                       (N167)? mem[160] : 
                       (N169)? mem[240] : 
                       (N171)? mem[320] : 
                       (N173)? mem[400] : 
                       (N175)? mem[480] : 
                       (N177)? mem[560] : 
                       (N179)? mem[640] : 
                       (N181)? mem[720] : 
                       (N183)? mem[800] : 
                       (N185)? mem[880] : 
                       (N187)? mem[960] : 
                       (N189)? mem[1040] : 
                       (N191)? mem[1120] : 
                       (N193)? mem[1200] : 
                       (N195)? mem[1280] : 
                       (N197)? mem[1360] : 
                       (N199)? mem[1440] : 
                       (N201)? mem[1520] : 
                       (N203)? mem[1600] : 
                       (N205)? mem[1680] : 
                       (N207)? mem[1760] : 
                       (N209)? mem[1840] : 
                       (N211)? mem[1920] : 
                       (N213)? mem[2000] : 
                       (N215)? mem[2080] : 
                       (N217)? mem[2160] : 
                       (N219)? mem[2240] : 
                       (N221)? mem[2320] : 
                       (N223)? mem[2400] : 
                       (N225)? mem[2480] : 
                       (N164)? mem[2560] : 
                       (N166)? mem[2640] : 
                       (N168)? mem[2720] : 
                       (N170)? mem[2800] : 
                       (N172)? mem[2880] : 
                       (N174)? mem[2960] : 
                       (N176)? mem[3040] : 
                       (N178)? mem[3120] : 
                       (N180)? mem[3200] : 
                       (N182)? mem[3280] : 
                       (N184)? mem[3360] : 
                       (N186)? mem[3440] : 
                       (N188)? mem[3520] : 
                       (N190)? mem[3600] : 
                       (N192)? mem[3680] : 
                       (N194)? mem[3760] : 
                       (N196)? mem[3840] : 
                       (N198)? mem[3920] : 
                       (N200)? mem[4000] : 
                       (N202)? mem[4080] : 
                       (N204)? mem[4160] : 
                       (N206)? mem[4240] : 
                       (N208)? mem[4320] : 
                       (N210)? mem[4400] : 
                       (N212)? mem[4480] : 
                       (N214)? mem[4560] : 
                       (N216)? mem[4640] : 
                       (N218)? mem[4720] : 
                       (N220)? mem[4800] : 
                       (N222)? mem[4880] : 
                       (N224)? mem[4960] : 
                       (N226)? mem[5040] : 1'b0;

  bsg_dff_width_p1
  llr_read_en_dff
  (
    .clk_i(clk_i),
    .data_i(read_en),
    .data_o(llr_read_en_r)
  );


  bsg_dff_en_bypass_width_p80
  llr_dff_bypass
  (
    .clk_i(clk_i),
    .en_i(llr_read_en_r),
    .data_i(data_out),
    .data_o(data_o)
  );

  assign N11497 = ~addr_i[5];
  assign N11498 = N11497 & N11539;
  assign N11499 = N11497 & N11540;
  assign N11500 = N11497 & N11541;
  assign N11501 = N11497 & N11542;
  assign N11502 = ~addr_i[2];
  assign N11503 = N11502 & N11551;
  assign N11504 = N11502 & N11552;
  assign N11505 = N11502 & N11553;
  assign N11506 = N11502 & N11554;
  assign N537 = N11507 & N11503;
  assign N536 = N11507 & N11504;
  assign N535 = N11507 & N11505;
  assign N534 = N11507 & N11506;
  assign N533 = N11508 & N11503;
  assign N532 = N11508 & N11504;
  assign N531 = N11508 & N11505;
  assign N530 = N11508 & N11506;
  assign N529 = N11509 & N11503;
  assign N528 = N11509 & N11504;
  assign N527 = N11509 & N11505;
  assign N526 = N11509 & N11506;
  assign N525 = N11546 & N11503;
  assign N524 = N11546 & N11504;
  assign N523 = N11546 & N11505;
  assign N522 = N11546 & N11506;
  assign N521 = N11498 & N11510;
  assign N520 = N11498 & N11511;
  assign N519 = N11498 & N11512;
  assign N518 = N11498 & N11558;
  assign N517 = N11498 & N11503;
  assign N516 = N11498 & N11504;
  assign N515 = N11498 & N11505;
  assign N514 = N11498 & N11506;
  assign N513 = N11499 & N11510;
  assign N512 = N11499 & N11511;
  assign N511 = N11499 & N11512;
  assign N510 = N11499 & N11558;
  assign N509 = N11499 & N11503;
  assign N508 = N11499 & N11504;
  assign N507 = N11499 & N11505;
  assign N506 = N11499 & N11506;
  assign N505 = N11500 & N11510;
  assign N504 = N11500 & N11511;
  assign N503 = N11500 & N11512;
  assign N502 = N11500 & N11558;
  assign N501 = N11500 & N11503;
  assign N500 = N11500 & N11504;
  assign N499 = N11500 & N11505;
  assign N498 = N11500 & N11506;
  assign N497 = N11501 & N11510;
  assign N496 = N11501 & N11511;
  assign N495 = N11501 & N11512;
  assign N494 = N11501 & N11558;
  assign N493 = N11501 & N11503;
  assign N492 = N11501 & N11504;
  assign N491 = N11501 & N11505;
  assign N490 = N11501 & N11506;
  assign N11507 = addr_i[5] & N11539;
  assign N11508 = addr_i[5] & N11540;
  assign N11509 = addr_i[5] & N11541;
  assign N11510 = addr_i[2] & N11551;
  assign N11511 = addr_i[2] & N11552;
  assign N11512 = addr_i[2] & N11553;
  assign N641 = N11507 & N11510;
  assign N640 = N11507 & N11511;
  assign N639 = N11507 & N11512;
  assign N638 = N11507 & N11558;
  assign N637 = N11507 & N11559;
  assign N636 = N11507 & N11560;
  assign N635 = N11507 & N11561;
  assign N634 = N11507 & N11562;
  assign N633 = N11508 & N11510;
  assign N632 = N11508 & N11511;
  assign N631 = N11508 & N11512;
  assign N630 = N11508 & N11558;
  assign N629 = N11508 & N11559;
  assign N628 = N11508 & N11560;
  assign N627 = N11508 & N11561;
  assign N626 = N11508 & N11562;
  assign N625 = N11509 & N11510;
  assign N624 = N11509 & N11511;
  assign N623 = N11509 & N11512;
  assign N622 = N11509 & N11558;
  assign N621 = N11509 & N11559;
  assign N620 = N11509 & N11560;
  assign N619 = N11509 & N11561;
  assign N618 = N11509 & N11562;
  assign N617 = N11546 & N11510;
  assign N616 = N11546 & N11511;
  assign N615 = N11546 & N11512;
  assign N614 = N11547 & N11510;
  assign N613 = N11547 & N11511;
  assign N612 = N11547 & N11512;
  assign N611 = N11548 & N11510;
  assign N610 = N11548 & N11511;
  assign N609 = N11548 & N11512;
  assign N608 = N11549 & N11510;
  assign N607 = N11549 & N11511;
  assign N606 = N11549 & N11512;
  assign N605 = N11550 & N11510;
  assign N604 = N11550 & N11511;
  assign N603 = N11550 & N11512;
  assign N972 = N11513 & N11558;
  assign N971 = N11514 & N11558;
  assign N970 = N11515 & N11558;
  assign N969 = N11546 & N11516;
  assign N968 = N11546 & N11517;
  assign N967 = N11546 & N11518;
  assign N1329 = N11513 & N11559;
  assign N1328 = N11513 & N11560;
  assign N1327 = N11513 & N11561;
  assign N1326 = N11513 & N11562;
  assign N1325 = N11514 & N11559;
  assign N1324 = N11514 & N11560;
  assign N1323 = N11514 & N11561;
  assign N1322 = N11514 & N11562;
  assign N1321 = N11515 & N11559;
  assign N1320 = N11515 & N11560;
  assign N1319 = N11515 & N11561;
  assign N1318 = N11515 & N11562;
  assign N1317 = N11529 & N11559;
  assign N1316 = N11529 & N11560;
  assign N1315 = N11529 & N11561;
  assign N1314 = N11529 & N11562;
  assign N1313 = N11547 & N11516;
  assign N1312 = N11547 & N11517;
  assign N1311 = N11547 & N11518;
  assign N1310 = N11547 & N11534;
  assign N1309 = N11548 & N11516;
  assign N1308 = N11548 & N11517;
  assign N1307 = N11548 & N11518;
  assign N1306 = N11548 & N11534;
  assign N1305 = N11549 & N11516;
  assign N1304 = N11549 & N11517;
  assign N1303 = N11549 & N11518;
  assign N1302 = N11549 & N11534;
  assign N1301 = N11550 & N11516;
  assign N1300 = N11550 & N11517;
  assign N1299 = N11550 & N11518;
  assign N1298 = N11550 & N11534;
  assign N11513 = addr_i[5] & N11539;
  assign N11514 = addr_i[5] & N11540;
  assign N11515 = addr_i[5] & N11541;
  assign N11516 = addr_i[2] & N11551;
  assign N11517 = addr_i[2] & N11552;
  assign N11518 = addr_i[2] & N11553;
  assign N1498 = N11513 & N11516;
  assign N1497 = N11513 & N11517;
  assign N1496 = N11513 & N11518;
  assign N1495 = N11513 & N11534;
  assign N1494 = N11513 & N11535;
  assign N1493 = N11513 & N11536;
  assign N1492 = N11513 & N11537;
  assign N1491 = N11513 & N11538;
  assign N1490 = N11514 & N11516;
  assign N1489 = N11514 & N11517;
  assign N1488 = N11514 & N11518;
  assign N1487 = N11514 & N11534;
  assign N1486 = N11514 & N11535;
  assign N1485 = N11514 & N11536;
  assign N1484 = N11514 & N11537;
  assign N1483 = N11514 & N11538;
  assign N1482 = N11515 & N11516;
  assign N1481 = N11515 & N11517;
  assign N1480 = N11515 & N11518;
  assign N1479 = N11515 & N11534;
  assign N1478 = N11515 & N11535;
  assign N1477 = N11515 & N11536;
  assign N1476 = N11515 & N11537;
  assign N1475 = N11515 & N11538;
  assign N1474 = N11529 & N11516;
  assign N1473 = N11529 & N11517;
  assign N1472 = N11529 & N11518;
  assign N1471 = N11530 & N11516;
  assign N1470 = N11530 & N11517;
  assign N1469 = N11530 & N11518;
  assign N1468 = N11531 & N11516;
  assign N1467 = N11531 & N11517;
  assign N1466 = N11531 & N11518;
  assign N1465 = N11532 & N11516;
  assign N1464 = N11532 & N11517;
  assign N1463 = N11532 & N11518;
  assign N1462 = N11533 & N11516;
  assign N1461 = N11533 & N11517;
  assign N1460 = N11533 & N11518;
  assign N2091 = N11519 & N11535;
  assign N2090 = N11519 & N11536;
  assign N2089 = N11519 & N11537;
  assign N2088 = N11519 & N11538;
  assign N2087 = N11530 & N11524;
  assign N2086 = N11531 & N11524;
  assign N2085 = N11532 & N11524;
  assign N2084 = N11533 & N11524;
  assign N11519 = addr_i[5] & N11542;
  assign N11520 = N11497 & N11539;
  assign N11521 = N11497 & N11540;
  assign N11522 = N11497 & N11541;
  assign N11523 = N11497 & N11542;
  assign N11524 = addr_i[2] & N11554;
  assign N11525 = N11502 & N11551;
  assign N11526 = N11502 & N11552;
  assign N11527 = N11502 & N11553;
  assign N11528 = N11502 & N11554;
  assign N2211 = N11543 & N11524;
  assign N2210 = N11543 & N11525;
  assign N2209 = N11543 & N11526;
  assign N2208 = N11543 & N11527;
  assign N2207 = N11543 & N11528;
  assign N2206 = N11544 & N11524;
  assign N2205 = N11544 & N11525;
  assign N2204 = N11544 & N11526;
  assign N2203 = N11544 & N11527;
  assign N2202 = N11544 & N11528;
  assign N2201 = N11545 & N11524;
  assign N2200 = N11545 & N11525;
  assign N2199 = N11545 & N11526;
  assign N2198 = N11545 & N11527;
  assign N2197 = N11545 & N11528;
  assign N2196 = N11519 & N11555;
  assign N2195 = N11519 & N11556;
  assign N2194 = N11519 & N11557;
  assign N2193 = N11519 & N11524;
  assign N2192 = N11519 & N11525;
  assign N2191 = N11519 & N11526;
  assign N2190 = N11519 & N11527;
  assign N2189 = N11519 & N11528;
  assign N2188 = N11520 & N11555;
  assign N2187 = N11520 & N11556;
  assign N2186 = N11520 & N11557;
  assign N2185 = N11520 & N11524;
  assign N2184 = N11520 & N11525;
  assign N2183 = N11520 & N11526;
  assign N2182 = N11520 & N11527;
  assign N2181 = N11520 & N11528;
  assign N2180 = N11521 & N11555;
  assign N2179 = N11521 & N11556;
  assign N2178 = N11521 & N11557;
  assign N2177 = N11521 & N11524;
  assign N2176 = N11521 & N11525;
  assign N2175 = N11521 & N11526;
  assign N2174 = N11521 & N11527;
  assign N2173 = N11521 & N11528;
  assign N2172 = N11522 & N11555;
  assign N2171 = N11522 & N11556;
  assign N2170 = N11522 & N11557;
  assign N2169 = N11522 & N11524;
  assign N2168 = N11522 & N11525;
  assign N2167 = N11522 & N11526;
  assign N2166 = N11522 & N11527;
  assign N2165 = N11522 & N11528;
  assign N2164 = N11523 & N11555;
  assign N2163 = N11523 & N11556;
  assign N2162 = N11523 & N11557;
  assign N2161 = N11523 & N11524;
  assign N2160 = N11523 & N11525;
  assign N2159 = N11523 & N11526;
  assign N2158 = N11523 & N11527;
  assign N2157 = N11523 & N11528;
  assign N11529 = addr_i[5] & N11542;
  assign N11530 = N11497 & N11539;
  assign N11531 = N11497 & N11540;
  assign N11532 = N11497 & N11541;
  assign N11533 = N11497 & N11542;
  assign N11534 = addr_i[2] & N11554;
  assign N11535 = N11502 & N11551;
  assign N11536 = N11502 & N11552;
  assign N11537 = N11502 & N11553;
  assign N11538 = N11502 & N11554;
  assign N2331 = N11543 & N11534;
  assign N2330 = N11543 & N11535;
  assign N2329 = N11543 & N11536;
  assign N2328 = N11543 & N11537;
  assign N2327 = N11543 & N11538;
  assign N2326 = N11544 & N11534;
  assign N2325 = N11544 & N11535;
  assign N2324 = N11544 & N11536;
  assign N2323 = N11544 & N11537;
  assign N2322 = N11544 & N11538;
  assign N2321 = N11545 & N11534;
  assign N2320 = N11545 & N11535;
  assign N2319 = N11545 & N11536;
  assign N2318 = N11545 & N11537;
  assign N2317 = N11545 & N11538;
  assign N2316 = N11529 & N11555;
  assign N2315 = N11529 & N11556;
  assign N2314 = N11529 & N11557;
  assign N2313 = N11529 & N11534;
  assign N2312 = N11529 & N11535;
  assign N2311 = N11529 & N11536;
  assign N2310 = N11529 & N11537;
  assign N2309 = N11529 & N11538;
  assign N2308 = N11530 & N11555;
  assign N2307 = N11530 & N11556;
  assign N2306 = N11530 & N11557;
  assign N2305 = N11530 & N11534;
  assign N2304 = N11530 & N11535;
  assign N2303 = N11530 & N11536;
  assign N2302 = N11530 & N11537;
  assign N2301 = N11530 & N11538;
  assign N2300 = N11531 & N11555;
  assign N2299 = N11531 & N11556;
  assign N2298 = N11531 & N11557;
  assign N2297 = N11531 & N11534;
  assign N2296 = N11531 & N11535;
  assign N2295 = N11531 & N11536;
  assign N2294 = N11531 & N11537;
  assign N2293 = N11531 & N11538;
  assign N2292 = N11532 & N11555;
  assign N2291 = N11532 & N11556;
  assign N2290 = N11532 & N11557;
  assign N2289 = N11532 & N11534;
  assign N2288 = N11532 & N11535;
  assign N2287 = N11532 & N11536;
  assign N2286 = N11532 & N11537;
  assign N2285 = N11532 & N11538;
  assign N2284 = N11533 & N11555;
  assign N2283 = N11533 & N11556;
  assign N2282 = N11533 & N11557;
  assign N2281 = N11533 & N11534;
  assign N2280 = N11533 & N11535;
  assign N2279 = N11533 & N11536;
  assign N2278 = N11533 & N11537;
  assign N2277 = N11533 & N11538;
  assign N11539 = addr_i[3] & addr_i[4];
  assign N11540 = N0 & addr_i[4];
  assign N0 = ~addr_i[3];
  assign N11541 = addr_i[3] & N1;
  assign N1 = ~addr_i[4];
  assign N11542 = N2 & N3;
  assign N2 = ~addr_i[3];
  assign N3 = ~addr_i[4];
  assign N11543 = addr_i[5] & N11539;
  assign N11544 = addr_i[5] & N11540;
  assign N11545 = addr_i[5] & N11541;
  assign N11546 = addr_i[5] & N11542;
  assign N11547 = N11497 & N11539;
  assign N11548 = N11497 & N11540;
  assign N11549 = N11497 & N11541;
  assign N11550 = N11497 & N11542;
  assign N11551 = addr_i[0] & addr_i[1];
  assign N11552 = N4 & addr_i[1];
  assign N4 = ~addr_i[0];
  assign N11553 = addr_i[0] & N5;
  assign N5 = ~addr_i[1];
  assign N11554 = N6 & N7;
  assign N6 = ~addr_i[0];
  assign N7 = ~addr_i[1];
  assign N11555 = addr_i[2] & N11551;
  assign N11556 = addr_i[2] & N11552;
  assign N11557 = addr_i[2] & N11553;
  assign N11558 = addr_i[2] & N11554;
  assign N11559 = N11502 & N11551;
  assign N11560 = N11502 & N11552;
  assign N11561 = N11502 & N11553;
  assign N11562 = N11502 & N11554;
  assign N2460 = N11543 & N11555;
  assign N2459 = N11543 & N11556;
  assign N2458 = N11543 & N11557;
  assign N2457 = N11543 & N11558;
  assign N2456 = N11543 & N11559;
  assign N2455 = N11543 & N11560;
  assign N2454 = N11543 & N11561;
  assign N2453 = N11543 & N11562;
  assign N2452 = N11544 & N11555;
  assign N2451 = N11544 & N11556;
  assign N2450 = N11544 & N11557;
  assign N2449 = N11544 & N11558;
  assign N2448 = N11544 & N11559;
  assign N2447 = N11544 & N11560;
  assign N2446 = N11544 & N11561;
  assign N2445 = N11544 & N11562;
  assign N2444 = N11545 & N11555;
  assign N2443 = N11545 & N11556;
  assign N2442 = N11545 & N11557;
  assign N2441 = N11545 & N11558;
  assign N2440 = N11545 & N11559;
  assign N2439 = N11545 & N11560;
  assign N2438 = N11545 & N11561;
  assign N2437 = N11545 & N11562;
  assign N2436 = N11546 & N11555;
  assign N2435 = N11546 & N11556;
  assign N2434 = N11546 & N11557;
  assign N2433 = N11546 & N11558;
  assign N2432 = N11546 & N11559;
  assign N2431 = N11546 & N11560;
  assign N2430 = N11546 & N11561;
  assign N2429 = N11546 & N11562;
  assign N2428 = N11547 & N11555;
  assign N2427 = N11547 & N11556;
  assign N2426 = N11547 & N11557;
  assign N2425 = N11547 & N11558;
  assign N2424 = N11547 & N11559;
  assign N2423 = N11547 & N11560;
  assign N2422 = N11547 & N11561;
  assign N2421 = N11547 & N11562;
  assign N2420 = N11548 & N11555;
  assign N2419 = N11548 & N11556;
  assign N2418 = N11548 & N11557;
  assign N2417 = N11548 & N11558;
  assign N2416 = N11548 & N11559;
  assign N2415 = N11548 & N11560;
  assign N2414 = N11548 & N11561;
  assign N2413 = N11548 & N11562;
  assign N2412 = N11549 & N11555;
  assign N2411 = N11549 & N11556;
  assign N2410 = N11549 & N11557;
  assign N2409 = N11549 & N11558;
  assign N2408 = N11549 & N11559;
  assign N2407 = N11549 & N11560;
  assign N2406 = N11549 & N11561;
  assign N2405 = N11549 & N11562;
  assign N2404 = N11550 & N11555;
  assign N2403 = N11550 & N11556;
  assign N2402 = N11550 & N11557;
  assign N2401 = N11550 & N11558;
  assign N2400 = N11550 & N11559;
  assign N2399 = N11550 & N11560;
  assign N2398 = N11550 & N11561;
  assign N2397 = N11550 & N11562;
  assign N11563 = addr_i[5] & N11635;
  assign N11564 = addr_i[5] & N11636;
  assign N11565 = addr_i[5] & N11637;
  assign N11566 = addr_i[2] & N11647;
  assign N11567 = addr_i[2] & N11648;
  assign N11568 = addr_i[2] & N11649;
  assign N2629 = N11563 & N11566;
  assign N2628 = N11563 & N11567;
  assign N2627 = N11563 & N11568;
  assign N2626 = N11563 & N11654;
  assign N2625 = N11563 & N11595;
  assign N2624 = N11563 & N11596;
  assign N2623 = N11563 & N11597;
  assign N2622 = N11563 & N11598;
  assign N2621 = N11564 & N11566;
  assign N2620 = N11564 & N11567;
  assign N2619 = N11564 & N11568;
  assign N2618 = N11564 & N11654;
  assign N2617 = N11564 & N11595;
  assign N2616 = N11564 & N11596;
  assign N2615 = N11564 & N11597;
  assign N2614 = N11564 & N11598;
  assign N2613 = N11565 & N11566;
  assign N2612 = N11565 & N11567;
  assign N2611 = N11565 & N11568;
  assign N2610 = N11565 & N11654;
  assign N2609 = N11565 & N11595;
  assign N2608 = N11565 & N11596;
  assign N2607 = N11565 & N11597;
  assign N2606 = N11565 & N11598;
  assign N2605 = N11642 & N11566;
  assign N2604 = N11642 & N11567;
  assign N2603 = N11642 & N11568;
  assign N2602 = N11591 & N11566;
  assign N2601 = N11591 & N11567;
  assign N2600 = N11591 & N11568;
  assign N2599 = N11592 & N11566;
  assign N2598 = N11592 & N11567;
  assign N2597 = N11592 & N11568;
  assign N2596 = N11593 & N11566;
  assign N2595 = N11593 & N11567;
  assign N2594 = N11593 & N11568;
  assign N2593 = N11594 & N11566;
  assign N2592 = N11594 & N11567;
  assign N2591 = N11594 & N11568;
  assign N3252 = N11569 & N11654;
  assign N3251 = N11569 & N11595;
  assign N3250 = N11569 & N11596;
  assign N3249 = N11569 & N11597;
  assign N3248 = N11569 & N11598;
  assign N3247 = N11570 & N11654;
  assign N3246 = N11570 & N11595;
  assign N3245 = N11570 & N11596;
  assign N3244 = N11570 & N11597;
  assign N3243 = N11570 & N11598;
  assign N3242 = N11571 & N11654;
  assign N3241 = N11571 & N11595;
  assign N3240 = N11571 & N11596;
  assign N3239 = N11571 & N11597;
  assign N3238 = N11571 & N11598;
  assign N3237 = N11642 & N11572;
  assign N3236 = N11642 & N11573;
  assign N3235 = N11642 & N11574;
  assign N3234 = N11642 & N11595;
  assign N3233 = N11642 & N11596;
  assign N3232 = N11642 & N11597;
  assign N3231 = N11642 & N11598;
  assign N3230 = N11591 & N11572;
  assign N3229 = N11591 & N11573;
  assign N3228 = N11591 & N11574;
  assign N3227 = N11591 & N11654;
  assign N3226 = N11592 & N11572;
  assign N3225 = N11592 & N11573;
  assign N3224 = N11592 & N11574;
  assign N3223 = N11592 & N11654;
  assign N3222 = N11593 & N11572;
  assign N3221 = N11593 & N11573;
  assign N3220 = N11593 & N11574;
  assign N3219 = N11593 & N11654;
  assign N3218 = N11594 & N11572;
  assign N3217 = N11594 & N11573;
  assign N3216 = N11594 & N11574;
  assign N3215 = N11594 & N11654;
  assign N11569 = addr_i[5] & N11635;
  assign N11570 = addr_i[5] & N11636;
  assign N11571 = addr_i[5] & N11637;
  assign N11572 = addr_i[2] & N11647;
  assign N11573 = addr_i[2] & N11648;
  assign N11574 = addr_i[2] & N11649;
  assign N3486 = N11569 & N11572;
  assign N3485 = N11569 & N11573;
  assign N3484 = N11569 & N11574;
  assign N3483 = N11569 & N11630;
  assign N3482 = N11569 & N11587;
  assign N3481 = N11569 & N11588;
  assign N3480 = N11569 & N11589;
  assign N3479 = N11569 & N11590;
  assign N3478 = N11570 & N11572;
  assign N3477 = N11570 & N11573;
  assign N3476 = N11570 & N11574;
  assign N3475 = N11570 & N11630;
  assign N3474 = N11570 & N11587;
  assign N3473 = N11570 & N11588;
  assign N3472 = N11570 & N11589;
  assign N3471 = N11570 & N11590;
  assign N3470 = N11571 & N11572;
  assign N3469 = N11571 & N11573;
  assign N3468 = N11571 & N11574;
  assign N3467 = N11571 & N11630;
  assign N3466 = N11571 & N11587;
  assign N3465 = N11571 & N11588;
  assign N3464 = N11571 & N11589;
  assign N3463 = N11571 & N11590;
  assign N3462 = N11625 & N11572;
  assign N3461 = N11625 & N11573;
  assign N3460 = N11625 & N11574;
  assign N3459 = N11583 & N11572;
  assign N3458 = N11583 & N11573;
  assign N3457 = N11583 & N11574;
  assign N3456 = N11584 & N11572;
  assign N3455 = N11584 & N11573;
  assign N3454 = N11584 & N11574;
  assign N3453 = N11585 & N11572;
  assign N3452 = N11585 & N11573;
  assign N3451 = N11585 & N11574;
  assign N3450 = N11586 & N11572;
  assign N3449 = N11586 & N11573;
  assign N3448 = N11586 & N11574;
  assign N4020 = N11599 & N11630;
  assign N4019 = N11600 & N11630;
  assign N4018 = N11601 & N11630;
  assign N4017 = N11625 & N11602;
  assign N4016 = N11625 & N11603;
  assign N4015 = N11625 & N11604;
  assign N4014 = N11625 & N11587;
  assign N4013 = N11625 & N11588;
  assign N4012 = N11625 & N11589;
  assign N4011 = N11625 & N11590;
  assign N4010 = N11583 & N11630;
  assign N4009 = N11584 & N11630;
  assign N4008 = N11585 & N11630;
  assign N4007 = N11586 & N11630;
  assign N11575 = N11497 & N11635;
  assign N11576 = N11497 & N11636;
  assign N11577 = N11497 & N11637;
  assign N11578 = N11497 & N11638;
  assign N11579 = N11502 & N11647;
  assign N11580 = N11502 & N11648;
  assign N11581 = N11502 & N11649;
  assign N11582 = N11502 & N11650;
  assign N4133 = N11599 & N11579;
  assign N4132 = N11599 & N11580;
  assign N4131 = N11599 & N11581;
  assign N4130 = N11599 & N11582;
  assign N4129 = N11600 & N11579;
  assign N4128 = N11600 & N11580;
  assign N4127 = N11600 & N11581;
  assign N4126 = N11600 & N11582;
  assign N4125 = N11601 & N11579;
  assign N4124 = N11601 & N11580;
  assign N4123 = N11601 & N11581;
  assign N4122 = N11601 & N11582;
  assign N4121 = N11615 & N11579;
  assign N4120 = N11615 & N11580;
  assign N4119 = N11615 & N11581;
  assign N4118 = N11615 & N11582;
  assign N4117 = N11575 & N11602;
  assign N4116 = N11575 & N11603;
  assign N4115 = N11575 & N11604;
  assign N4114 = N11575 & N11620;
  assign N4113 = N11575 & N11579;
  assign N4112 = N11575 & N11580;
  assign N4111 = N11575 & N11581;
  assign N4110 = N11575 & N11582;
  assign N4109 = N11576 & N11602;
  assign N4108 = N11576 & N11603;
  assign N4107 = N11576 & N11604;
  assign N4106 = N11576 & N11620;
  assign N4105 = N11576 & N11579;
  assign N4104 = N11576 & N11580;
  assign N4103 = N11576 & N11581;
  assign N4102 = N11576 & N11582;
  assign N4101 = N11577 & N11602;
  assign N4100 = N11577 & N11603;
  assign N4099 = N11577 & N11604;
  assign N4098 = N11577 & N11620;
  assign N4097 = N11577 & N11579;
  assign N4096 = N11577 & N11580;
  assign N4095 = N11577 & N11581;
  assign N4094 = N11577 & N11582;
  assign N4093 = N11578 & N11602;
  assign N4092 = N11578 & N11603;
  assign N4091 = N11578 & N11604;
  assign N4090 = N11578 & N11620;
  assign N4089 = N11578 & N11579;
  assign N4088 = N11578 & N11580;
  assign N4087 = N11578 & N11581;
  assign N4086 = N11578 & N11582;
  assign N11583 = N11497 & N11635;
  assign N11584 = N11497 & N11636;
  assign N11585 = N11497 & N11637;
  assign N11586 = N11497 & N11638;
  assign N11587 = N11502 & N11647;
  assign N11588 = N11502 & N11648;
  assign N11589 = N11502 & N11649;
  assign N11590 = N11502 & N11650;
  assign N4246 = N11599 & N11587;
  assign N4245 = N11599 & N11588;
  assign N4244 = N11599 & N11589;
  assign N4243 = N11599 & N11590;
  assign N4242 = N11600 & N11587;
  assign N4241 = N11600 & N11588;
  assign N4240 = N11600 & N11589;
  assign N4239 = N11600 & N11590;
  assign N4238 = N11601 & N11587;
  assign N4237 = N11601 & N11588;
  assign N4236 = N11601 & N11589;
  assign N4235 = N11601 & N11590;
  assign N4234 = N11615 & N11587;
  assign N4233 = N11615 & N11588;
  assign N4232 = N11615 & N11589;
  assign N4231 = N11615 & N11590;
  assign N4230 = N11583 & N11602;
  assign N4229 = N11583 & N11603;
  assign N4228 = N11583 & N11604;
  assign N4227 = N11583 & N11620;
  assign N4226 = N11583 & N11587;
  assign N4225 = N11583 & N11588;
  assign N4224 = N11583 & N11589;
  assign N4223 = N11583 & N11590;
  assign N4222 = N11584 & N11602;
  assign N4221 = N11584 & N11603;
  assign N4220 = N11584 & N11604;
  assign N4219 = N11584 & N11620;
  assign N4218 = N11584 & N11587;
  assign N4217 = N11584 & N11588;
  assign N4216 = N11584 & N11589;
  assign N4215 = N11584 & N11590;
  assign N4214 = N11585 & N11602;
  assign N4213 = N11585 & N11603;
  assign N4212 = N11585 & N11604;
  assign N4211 = N11585 & N11620;
  assign N4210 = N11585 & N11587;
  assign N4209 = N11585 & N11588;
  assign N4208 = N11585 & N11589;
  assign N4207 = N11585 & N11590;
  assign N4206 = N11586 & N11602;
  assign N4205 = N11586 & N11603;
  assign N4204 = N11586 & N11604;
  assign N4203 = N11586 & N11620;
  assign N4202 = N11586 & N11587;
  assign N4201 = N11586 & N11588;
  assign N4200 = N11586 & N11589;
  assign N4199 = N11586 & N11590;
  assign N11591 = N11497 & N11635;
  assign N11592 = N11497 & N11636;
  assign N11593 = N11497 & N11637;
  assign N11594 = N11497 & N11638;
  assign N11595 = N11502 & N11647;
  assign N11596 = N11502 & N11648;
  assign N11597 = N11502 & N11649;
  assign N11598 = N11502 & N11650;
  assign N4359 = N11599 & N11595;
  assign N4358 = N11599 & N11596;
  assign N4357 = N11599 & N11597;
  assign N4356 = N11599 & N11598;
  assign N4355 = N11600 & N11595;
  assign N4354 = N11600 & N11596;
  assign N4353 = N11600 & N11597;
  assign N4352 = N11600 & N11598;
  assign N4351 = N11601 & N11595;
  assign N4350 = N11601 & N11596;
  assign N4349 = N11601 & N11597;
  assign N4348 = N11601 & N11598;
  assign N4347 = N11615 & N11595;
  assign N4346 = N11615 & N11596;
  assign N4345 = N11615 & N11597;
  assign N4344 = N11615 & N11598;
  assign N4343 = N11591 & N11602;
  assign N4342 = N11591 & N11603;
  assign N4341 = N11591 & N11604;
  assign N4340 = N11591 & N11620;
  assign N4339 = N11591 & N11595;
  assign N4338 = N11591 & N11596;
  assign N4337 = N11591 & N11597;
  assign N4336 = N11591 & N11598;
  assign N4335 = N11592 & N11602;
  assign N4334 = N11592 & N11603;
  assign N4333 = N11592 & N11604;
  assign N4332 = N11592 & N11620;
  assign N4331 = N11592 & N11595;
  assign N4330 = N11592 & N11596;
  assign N4329 = N11592 & N11597;
  assign N4328 = N11592 & N11598;
  assign N4327 = N11593 & N11602;
  assign N4326 = N11593 & N11603;
  assign N4325 = N11593 & N11604;
  assign N4324 = N11593 & N11620;
  assign N4323 = N11593 & N11595;
  assign N4322 = N11593 & N11596;
  assign N4321 = N11593 & N11597;
  assign N4320 = N11593 & N11598;
  assign N4319 = N11594 & N11602;
  assign N4318 = N11594 & N11603;
  assign N4317 = N11594 & N11604;
  assign N4316 = N11594 & N11620;
  assign N4315 = N11594 & N11595;
  assign N4314 = N11594 & N11596;
  assign N4313 = N11594 & N11597;
  assign N4312 = N11594 & N11598;
  assign N11599 = addr_i[5] & N11635;
  assign N11600 = addr_i[5] & N11636;
  assign N11601 = addr_i[5] & N11637;
  assign N11602 = addr_i[2] & N11647;
  assign N11603 = addr_i[2] & N11648;
  assign N11604 = addr_i[2] & N11649;
  assign N4463 = N11599 & N11602;
  assign N4462 = N11599 & N11603;
  assign N4461 = N11599 & N11604;
  assign N4460 = N11599 & N11620;
  assign N4459 = N11599 & N11655;
  assign N4458 = N11599 & N11656;
  assign N4457 = N11599 & N11657;
  assign N4456 = N11599 & N11658;
  assign N4455 = N11600 & N11602;
  assign N4454 = N11600 & N11603;
  assign N4453 = N11600 & N11604;
  assign N4452 = N11600 & N11620;
  assign N4451 = N11600 & N11655;
  assign N4450 = N11600 & N11656;
  assign N4449 = N11600 & N11657;
  assign N4448 = N11600 & N11658;
  assign N4447 = N11601 & N11602;
  assign N4446 = N11601 & N11603;
  assign N4445 = N11601 & N11604;
  assign N4444 = N11601 & N11620;
  assign N4443 = N11601 & N11655;
  assign N4442 = N11601 & N11656;
  assign N4441 = N11601 & N11657;
  assign N4440 = N11601 & N11658;
  assign N4439 = N11615 & N11602;
  assign N4438 = N11615 & N11603;
  assign N4437 = N11615 & N11604;
  assign N4436 = N11643 & N11602;
  assign N4435 = N11643 & N11603;
  assign N4434 = N11643 & N11604;
  assign N4433 = N11644 & N11602;
  assign N4432 = N11644 & N11603;
  assign N4431 = N11644 & N11604;
  assign N4430 = N11645 & N11602;
  assign N4429 = N11645 & N11603;
  assign N4428 = N11645 & N11604;
  assign N4427 = N11646 & N11602;
  assign N4426 = N11646 & N11603;
  assign N4425 = N11646 & N11604;
  assign N4932 = N11605 & N11620;
  assign N4931 = N11606 & N11620;
  assign N4930 = N11607 & N11620;
  assign N4929 = N11615 & N11608;
  assign N4928 = N11615 & N11609;
  assign N4927 = N11615 & N11610;
  assign N4926 = N11615 & N11655;
  assign N4925 = N11615 & N11656;
  assign N4924 = N11615 & N11657;
  assign N4923 = N11615 & N11658;
  assign N4922 = N11643 & N11620;
  assign N4921 = N11644 & N11620;
  assign N4920 = N11645 & N11620;
  assign N4919 = N11646 & N11620;
  assign N5159 = N11605 & N11655;
  assign N5158 = N11605 & N11656;
  assign N5157 = N11605 & N11657;
  assign N5156 = N11605 & N11658;
  assign N5155 = N11606 & N11655;
  assign N5154 = N11606 & N11656;
  assign N5153 = N11606 & N11657;
  assign N5152 = N11606 & N11658;
  assign N5151 = N11607 & N11655;
  assign N5150 = N11607 & N11656;
  assign N5149 = N11607 & N11657;
  assign N5148 = N11607 & N11658;
  assign N5147 = N11613 & N11655;
  assign N5146 = N11613 & N11656;
  assign N5145 = N11613 & N11657;
  assign N5144 = N11613 & N11658;
  assign N5143 = N11643 & N11608;
  assign N5142 = N11643 & N11609;
  assign N5141 = N11643 & N11610;
  assign N5140 = N11643 & N11614;
  assign N5139 = N11644 & N11608;
  assign N5138 = N11644 & N11609;
  assign N5137 = N11644 & N11610;
  assign N5136 = N11644 & N11614;
  assign N5135 = N11645 & N11608;
  assign N5134 = N11645 & N11609;
  assign N5133 = N11645 & N11610;
  assign N5132 = N11645 & N11614;
  assign N5131 = N11646 & N11608;
  assign N5130 = N11646 & N11609;
  assign N5129 = N11646 & N11610;
  assign N5128 = N11646 & N11614;
  assign N11605 = addr_i[5] & N11635;
  assign N11606 = addr_i[5] & N11636;
  assign N11607 = addr_i[5] & N11637;
  assign N11608 = addr_i[2] & N11647;
  assign N11609 = addr_i[2] & N11648;
  assign N11610 = addr_i[2] & N11649;
  assign N5328 = N11605 & N11608;
  assign N5327 = N11605 & N11609;
  assign N5326 = N11605 & N11610;
  assign N5325 = N11605 & N11614;
  assign N5324 = N11605 & N11631;
  assign N5323 = N11605 & N11632;
  assign N5322 = N11605 & N11633;
  assign N5321 = N11605 & N11634;
  assign N5320 = N11606 & N11608;
  assign N5319 = N11606 & N11609;
  assign N5318 = N11606 & N11610;
  assign N5317 = N11606 & N11614;
  assign N5316 = N11606 & N11631;
  assign N5315 = N11606 & N11632;
  assign N5314 = N11606 & N11633;
  assign N5313 = N11606 & N11634;
  assign N5312 = N11607 & N11608;
  assign N5311 = N11607 & N11609;
  assign N5310 = N11607 & N11610;
  assign N5309 = N11607 & N11614;
  assign N5308 = N11607 & N11631;
  assign N5307 = N11607 & N11632;
  assign N5306 = N11607 & N11633;
  assign N5305 = N11607 & N11634;
  assign N5304 = N11613 & N11608;
  assign N5303 = N11613 & N11609;
  assign N5302 = N11613 & N11610;
  assign N5301 = N11626 & N11608;
  assign N5300 = N11626 & N11609;
  assign N5299 = N11626 & N11610;
  assign N5298 = N11627 & N11608;
  assign N5297 = N11627 & N11609;
  assign N5296 = N11627 & N11610;
  assign N5295 = N11628 & N11608;
  assign N5294 = N11628 & N11609;
  assign N5293 = N11628 & N11610;
  assign N5292 = N11629 & N11608;
  assign N5291 = N11629 & N11609;
  assign N5290 = N11629 & N11610;
  assign N11611 = addr_i[5] & N11638;
  assign N11612 = addr_i[2] & N11650;
  assign N5863 = N11639 & N11612;
  assign N5862 = N11640 & N11612;
  assign N5861 = N11641 & N11612;
  assign N5860 = N11611 & N11651;
  assign N5859 = N11611 & N11652;
  assign N5858 = N11611 & N11653;
  assign N5857 = N11611 & N11612;
  assign N5856 = N11611 & N11631;
  assign N5855 = N11611 & N11632;
  assign N5854 = N11611 & N11633;
  assign N5853 = N11611 & N11634;
  assign N5852 = N11626 & N11612;
  assign N5851 = N11627 & N11612;
  assign N5850 = N11628 & N11612;
  assign N5849 = N11629 & N11612;
  assign N11613 = addr_i[5] & N11638;
  assign N11614 = addr_i[2] & N11650;
  assign N5943 = N11639 & N11614;
  assign N5942 = N11640 & N11614;
  assign N5941 = N11641 & N11614;
  assign N5940 = N11613 & N11651;
  assign N5939 = N11613 & N11652;
  assign N5938 = N11613 & N11653;
  assign N5937 = N11613 & N11614;
  assign N5936 = N11613 & N11631;
  assign N5935 = N11613 & N11632;
  assign N5934 = N11613 & N11633;
  assign N5933 = N11613 & N11634;
  assign N5932 = N11626 & N11614;
  assign N5931 = N11627 & N11614;
  assign N5930 = N11628 & N11614;
  assign N5929 = N11629 & N11614;
  assign N11615 = addr_i[5] & N11638;
  assign N11616 = N11497 & N11635;
  assign N11617 = N11497 & N11636;
  assign N11618 = N11497 & N11637;
  assign N11619 = N11497 & N11638;
  assign N11620 = addr_i[2] & N11650;
  assign N11621 = N11502 & N11647;
  assign N11622 = N11502 & N11648;
  assign N11623 = N11502 & N11649;
  assign N11624 = N11502 & N11650;
  assign N6063 = N11639 & N11620;
  assign N6062 = N11639 & N11621;
  assign N6061 = N11639 & N11622;
  assign N6060 = N11639 & N11623;
  assign N6059 = N11639 & N11624;
  assign N6058 = N11640 & N11620;
  assign N6057 = N11640 & N11621;
  assign N6056 = N11640 & N11622;
  assign N6055 = N11640 & N11623;
  assign N6054 = N11640 & N11624;
  assign N6053 = N11641 & N11620;
  assign N6052 = N11641 & N11621;
  assign N6051 = N11641 & N11622;
  assign N6050 = N11641 & N11623;
  assign N6049 = N11641 & N11624;
  assign N6048 = N11615 & N11651;
  assign N6047 = N11615 & N11652;
  assign N6046 = N11615 & N11653;
  assign N6045 = N11615 & N11620;
  assign N6044 = N11615 & N11621;
  assign N6043 = N11615 & N11622;
  assign N6042 = N11615 & N11623;
  assign N6041 = N11615 & N11624;
  assign N6040 = N11616 & N11651;
  assign N6039 = N11616 & N11652;
  assign N6038 = N11616 & N11653;
  assign N6037 = N11616 & N11620;
  assign N6036 = N11616 & N11621;
  assign N6035 = N11616 & N11622;
  assign N6034 = N11616 & N11623;
  assign N6033 = N11616 & N11624;
  assign N6032 = N11617 & N11651;
  assign N6031 = N11617 & N11652;
  assign N6030 = N11617 & N11653;
  assign N6029 = N11617 & N11620;
  assign N6028 = N11617 & N11621;
  assign N6027 = N11617 & N11622;
  assign N6026 = N11617 & N11623;
  assign N6025 = N11617 & N11624;
  assign N6024 = N11618 & N11651;
  assign N6023 = N11618 & N11652;
  assign N6022 = N11618 & N11653;
  assign N6021 = N11618 & N11620;
  assign N6020 = N11618 & N11621;
  assign N6019 = N11618 & N11622;
  assign N6018 = N11618 & N11623;
  assign N6017 = N11618 & N11624;
  assign N6016 = N11619 & N11651;
  assign N6015 = N11619 & N11652;
  assign N6014 = N11619 & N11653;
  assign N6013 = N11619 & N11620;
  assign N6012 = N11619 & N11621;
  assign N6011 = N11619 & N11622;
  assign N6010 = N11619 & N11623;
  assign N6009 = N11619 & N11624;
  assign N11625 = addr_i[5] & N11638;
  assign N11626 = N11497 & N11635;
  assign N11627 = N11497 & N11636;
  assign N11628 = N11497 & N11637;
  assign N11629 = N11497 & N11638;
  assign N11630 = addr_i[2] & N11650;
  assign N11631 = N11502 & N11647;
  assign N11632 = N11502 & N11648;
  assign N11633 = N11502 & N11649;
  assign N11634 = N11502 & N11650;
  assign N6183 = N11639 & N11630;
  assign N6182 = N11639 & N11631;
  assign N6181 = N11639 & N11632;
  assign N6180 = N11639 & N11633;
  assign N6179 = N11639 & N11634;
  assign N6178 = N11640 & N11630;
  assign N6177 = N11640 & N11631;
  assign N6176 = N11640 & N11632;
  assign N6175 = N11640 & N11633;
  assign N6174 = N11640 & N11634;
  assign N6173 = N11641 & N11630;
  assign N6172 = N11641 & N11631;
  assign N6171 = N11641 & N11632;
  assign N6170 = N11641 & N11633;
  assign N6169 = N11641 & N11634;
  assign N6168 = N11625 & N11651;
  assign N6167 = N11625 & N11652;
  assign N6166 = N11625 & N11653;
  assign N6165 = N11625 & N11630;
  assign N6164 = N11625 & N11631;
  assign N6163 = N11625 & N11632;
  assign N6162 = N11625 & N11633;
  assign N6161 = N11625 & N11634;
  assign N6160 = N11626 & N11651;
  assign N6159 = N11626 & N11652;
  assign N6158 = N11626 & N11653;
  assign N6157 = N11626 & N11630;
  assign N6156 = N11626 & N11631;
  assign N6155 = N11626 & N11632;
  assign N6154 = N11626 & N11633;
  assign N6153 = N11626 & N11634;
  assign N6152 = N11627 & N11651;
  assign N6151 = N11627 & N11652;
  assign N6150 = N11627 & N11653;
  assign N6149 = N11627 & N11630;
  assign N6148 = N11627 & N11631;
  assign N6147 = N11627 & N11632;
  assign N6146 = N11627 & N11633;
  assign N6145 = N11627 & N11634;
  assign N6144 = N11628 & N11651;
  assign N6143 = N11628 & N11652;
  assign N6142 = N11628 & N11653;
  assign N6141 = N11628 & N11630;
  assign N6140 = N11628 & N11631;
  assign N6139 = N11628 & N11632;
  assign N6138 = N11628 & N11633;
  assign N6137 = N11628 & N11634;
  assign N6136 = N11629 & N11651;
  assign N6135 = N11629 & N11652;
  assign N6134 = N11629 & N11653;
  assign N6133 = N11629 & N11630;
  assign N6132 = N11629 & N11631;
  assign N6131 = N11629 & N11632;
  assign N6130 = N11629 & N11633;
  assign N6129 = N11629 & N11634;
  assign N11635 = addr_i[3] & addr_i[4];
  assign N11636 = N8 & addr_i[4];
  assign N8 = ~addr_i[3];
  assign N11637 = addr_i[3] & N9;
  assign N9 = ~addr_i[4];
  assign N11638 = N10 & N11;
  assign N10 = ~addr_i[3];
  assign N11 = ~addr_i[4];
  assign N11639 = addr_i[5] & N11635;
  assign N11640 = addr_i[5] & N11636;
  assign N11641 = addr_i[5] & N11637;
  assign N11642 = addr_i[5] & N11638;
  assign N11643 = N11497 & N11635;
  assign N11644 = N11497 & N11636;
  assign N11645 = N11497 & N11637;
  assign N11646 = N11497 & N11638;
  assign N11647 = addr_i[0] & addr_i[1];
  assign N11648 = N12 & addr_i[1];
  assign N12 = ~addr_i[0];
  assign N11649 = addr_i[0] & N13;
  assign N13 = ~addr_i[1];
  assign N11650 = N14 & N15;
  assign N14 = ~addr_i[0];
  assign N15 = ~addr_i[1];
  assign N11651 = addr_i[2] & N11647;
  assign N11652 = addr_i[2] & N11648;
  assign N11653 = addr_i[2] & N11649;
  assign N11654 = addr_i[2] & N11650;
  assign N11655 = N11502 & N11647;
  assign N11656 = N11502 & N11648;
  assign N11657 = N11502 & N11649;
  assign N11658 = N11502 & N11650;
  assign N6312 = N11639 & N11651;
  assign N6311 = N11639 & N11652;
  assign N6310 = N11639 & N11653;
  assign N6309 = N11639 & N11654;
  assign N6308 = N11639 & N11655;
  assign N6307 = N11639 & N11656;
  assign N6306 = N11639 & N11657;
  assign N6305 = N11639 & N11658;
  assign N6304 = N11640 & N11651;
  assign N6303 = N11640 & N11652;
  assign N6302 = N11640 & N11653;
  assign N6301 = N11640 & N11654;
  assign N6300 = N11640 & N11655;
  assign N6299 = N11640 & N11656;
  assign N6298 = N11640 & N11657;
  assign N6297 = N11640 & N11658;
  assign N6296 = N11641 & N11651;
  assign N6295 = N11641 & N11652;
  assign N6294 = N11641 & N11653;
  assign N6293 = N11641 & N11654;
  assign N6292 = N11641 & N11655;
  assign N6291 = N11641 & N11656;
  assign N6290 = N11641 & N11657;
  assign N6289 = N11641 & N11658;
  assign N6288 = N11642 & N11651;
  assign N6287 = N11642 & N11652;
  assign N6286 = N11642 & N11653;
  assign N6285 = N11642 & N11654;
  assign N6284 = N11642 & N11655;
  assign N6283 = N11642 & N11656;
  assign N6282 = N11642 & N11657;
  assign N6281 = N11642 & N11658;
  assign N6280 = N11643 & N11651;
  assign N6279 = N11643 & N11652;
  assign N6278 = N11643 & N11653;
  assign N6277 = N11643 & N11654;
  assign N6276 = N11643 & N11655;
  assign N6275 = N11643 & N11656;
  assign N6274 = N11643 & N11657;
  assign N6273 = N11643 & N11658;
  assign N6272 = N11644 & N11651;
  assign N6271 = N11644 & N11652;
  assign N6270 = N11644 & N11653;
  assign N6269 = N11644 & N11654;
  assign N6268 = N11644 & N11655;
  assign N6267 = N11644 & N11656;
  assign N6266 = N11644 & N11657;
  assign N6265 = N11644 & N11658;
  assign N6264 = N11645 & N11651;
  assign N6263 = N11645 & N11652;
  assign N6262 = N11645 & N11653;
  assign N6261 = N11645 & N11654;
  assign N6260 = N11645 & N11655;
  assign N6259 = N11645 & N11656;
  assign N6258 = N11645 & N11657;
  assign N6257 = N11645 & N11658;
  assign N6256 = N11646 & N11651;
  assign N6255 = N11646 & N11652;
  assign N6254 = N11646 & N11653;
  assign N6253 = N11646 & N11654;
  assign N6252 = N11646 & N11655;
  assign N6251 = N11646 & N11656;
  assign N6250 = N11646 & N11657;
  assign N6249 = N11646 & N11658;
  assign { N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230 } = (N16)? { N641, N640, N639, N638, N537, N536, N535, N534, N633, N632, N631, N630, N533, N532, N531, N530, N625, N624, N623, N622, N529, N528, N527, N526, N617, N616, N615, N2433, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N229)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = w_mask_i[0];
  assign { N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295 } = (N17)? { N641, N640, N639, N638, N537, N536, N535, N534, N633, N632, N631, N630, N533, N532, N531, N530, N625, N624, N623, N622, N529, N528, N527, N526, N617, N616, N615, N2433, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N294)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N17 = w_mask_i[1];
  assign { N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360 } = (N18)? { N641, N640, N639, N638, N537, N536, N535, N534, N633, N632, N631, N630, N533, N532, N531, N530, N625, N624, N623, N622, N529, N528, N527, N526, N617, N616, N615, N2433, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N359)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N18 = w_mask_i[2];
  assign { N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425 } = (N19)? { N641, N640, N639, N638, N537, N536, N535, N534, N633, N632, N631, N630, N533, N532, N531, N530, N625, N624, N623, N622, N529, N528, N527, N526, N617, N616, N615, N2433, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N424)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N19 = w_mask_i[3];
  assign { N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538 } = (N20)? { N641, N640, N639, N638, N537, N536, N535, N534, N633, N632, N631, N630, N533, N532, N531, N530, N625, N624, N623, N622, N529, N528, N527, N526, N617, N616, N615, N2433, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N489)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N20 = w_mask_i[4];
  assign { N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642 } = (N21)? { N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N2433, N2432, N2431, N2430, N2429, N614, N613, N612, N2425, N2424, N2423, N2422, N2421, N611, N610, N609, N2417, N2416, N2415, N2414, N2413, N608, N607, N606, N2409, N2408, N2407, N2406, N2405, N605, N604, N603, N2401, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N602)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N21 = w_mask_i[5];
  assign { N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707 } = (N22)? { N1498, N1497, N1496, N972, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N971, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N970, N1321, N1320, N1319, N1318, N969, N968, N967, N2433, N2432, N2431, N2430, N2429, N1313, N1312, N1311, N2425, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N2417, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N2409, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N2401, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N706)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N22 = w_mask_i[6];
  assign { N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772 } = (N23)? { N1498, N1497, N1496, N972, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N971, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N970, N1321, N1320, N1319, N1318, N969, N968, N967, N2433, N2432, N2431, N2430, N2429, N1313, N1312, N1311, N2425, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N2417, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N2409, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N2401, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N771)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N23 = w_mask_i[7];
  assign { N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837 } = (N24)? { N1498, N1497, N1496, N972, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N971, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N970, N1321, N1320, N1319, N1318, N969, N968, N967, N2433, N2432, N2431, N2430, N2429, N1313, N1312, N1311, N2425, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N2417, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N2409, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N2401, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N836)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N24 = w_mask_i[8];
  assign { N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902 } = (N25)? { N1498, N1497, N1496, N972, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N971, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N970, N1321, N1320, N1319, N1318, N969, N968, N967, N2433, N2432, N2431, N2430, N2429, N1313, N1312, N1311, N2425, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N2417, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N2409, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N2401, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N901)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N25 = w_mask_i[9];
  assign { N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973 } = (N26)? { N1498, N1497, N1496, N972, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N971, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N970, N1321, N1320, N1319, N1318, N969, N968, N967, N2433, N2432, N2431, N2430, N2429, N1313, N1312, N1311, N2425, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N2417, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N2409, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N2401, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                   (N966)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N26 = w_mask_i[10];
  assign { N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038 } = (N27)? { N1498, N1497, N1496, N1495, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N1487, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N1479, N1321, N1320, N1319, N1318, N1474, N1473, N1472, N2313, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N1306, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N1302, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N1298, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1037)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N27 = w_mask_i[11];
  assign { N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103 } = (N28)? { N1498, N1497, N1496, N1495, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N1487, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N1479, N1321, N1320, N1319, N1318, N1474, N1473, N1472, N2313, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N1306, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N1302, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N1298, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1102)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N28 = w_mask_i[12];
  assign { N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168 } = (N29)? { N1498, N1497, N1496, N1495, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N1487, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N1479, N1321, N1320, N1319, N1318, N1474, N1473, N1472, N2313, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N1306, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N1302, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N1298, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1167)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N29 = w_mask_i[13];
  assign { N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233 } = (N30)? { N1498, N1497, N1496, N1495, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N1487, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N1479, N1321, N1320, N1319, N1318, N1474, N1473, N1472, N2313, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N1306, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N1302, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N1298, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1232)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N30 = w_mask_i[14];
  assign { N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330 } = (N31)? { N1498, N1497, N1496, N1495, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N1487, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N1479, N1321, N1320, N1319, N1318, N1474, N1473, N1472, N2313, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N1306, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N1302, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N1298, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1297)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N31 = w_mask_i[15];
  assign { N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395 } = (N32)? { N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N2313, N2312, N2311, N2310, N2309, N1471, N1470, N1469, N2305, N2304, N2303, N2302, N2301, N1468, N1467, N1466, N2297, N2296, N2295, N2294, N2293, N1465, N1464, N1463, N2289, N2288, N2287, N2286, N2285, N1462, N1461, N1460, N2281, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1394)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N32 = w_mask_i[16];
  assign { N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499 } = (N33)? { N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N2313, N2312, N2311, N2310, N2309, N1471, N1470, N1469, N2305, N2304, N2303, N2302, N2301, N1468, N1467, N1466, N2297, N2296, N2295, N2294, N2293, N1465, N1464, N1463, N2289, N2288, N2287, N2286, N2285, N1462, N1461, N1460, N2281, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1459)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N33 = w_mask_i[17];
  assign { N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564 } = (N34)? { N2460, N2459, N2458, N2331, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2326, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1563)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N34 = w_mask_i[18];
  assign { N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629 } = (N35)? { N2460, N2459, N2458, N2331, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2326, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1628)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N35 = w_mask_i[19];
  assign { N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694 } = (N36)? { N2460, N2459, N2458, N2331, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2326, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1693)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N36 = w_mask_i[20];
  assign { N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759 } = (N37)? { N2460, N2459, N2458, N2331, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2326, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1758)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N37 = w_mask_i[21];
  assign { N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824 } = (N38)? { N2460, N2459, N2458, N2211, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2206, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2201, N2320, N2319, N2318, N2317, N2196, N2195, N2194, N2193, N2091, N2090, N2089, N2088, N2308, N2307, N2306, N2087, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2086, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2085, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2084, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1823)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N38 = w_mask_i[22];
  assign { N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889 } = (N39)? { N2460, N2459, N2458, N2211, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2206, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2201, N2320, N2319, N2318, N2317, N2196, N2195, N2194, N2193, N2091, N2090, N2089, N2088, N2308, N2307, N2306, N2087, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2086, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2085, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2084, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1888)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N39 = w_mask_i[23];
  assign { N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954 } = (N40)? { N2460, N2459, N2458, N2211, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2206, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2201, N2320, N2319, N2318, N2317, N2196, N2195, N2194, N2193, N2091, N2090, N2089, N2088, N2308, N2307, N2306, N2087, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2086, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2085, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2084, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1953)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N40 = w_mask_i[24];
  assign { N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036, N2035, N2034, N2033, N2032, N2031, N2030, N2029, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019 } = (N41)? { N2460, N2459, N2458, N2211, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2206, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2201, N2320, N2319, N2318, N2317, N2196, N2195, N2194, N2193, N2091, N2090, N2089, N2088, N2308, N2307, N2306, N2087, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2086, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2085, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2084, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2018)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N41 = w_mask_i[25];
  assign { N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092 } = (N42)? { N2460, N2459, N2458, N2211, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2206, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2201, N2320, N2319, N2318, N2317, N2196, N2195, N2194, N2193, N2091, N2090, N2089, N2088, N2308, N2307, N2306, N2087, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2086, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2085, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2084, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2083)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N42 = w_mask_i[26];
  assign { N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248, N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229, N2228, N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215, N2214, N2213, N2212 } = (N43)? { N2460, N2459, N2458, N2211, N2210, N2209, N2208, N2207, N2452, N2451, N2450, N2206, N2205, N2204, N2203, N2202, N2444, N2443, N2442, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174, N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2156)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N43 = w_mask_i[27];
  assign { N2395, N2394, N2393, N2392, N2391, N2390, N2389, N2388, N2387, N2386, N2385, N2384, N2383, N2382, N2381, N2380, N2379, N2378, N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, N2368, N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, N2358, N2357, N2356, N2355, N2354, N2353, N2352, N2351, N2350, N2349, N2348, N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340, N2339, N2338, N2337, N2336, N2335, N2334, N2333, N2332 } = (N44)? { N2460, N2459, N2458, N2331, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2326, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2276)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N44 = w_mask_i[28];
  assign { N2524, N2523, N2522, N2521, N2520, N2519, N2518, N2517, N2516, N2515, N2514, N2513, N2512, N2511, N2510, N2509, N2508, N2507, N2506, N2505, N2504, N2503, N2502, N2501, N2500, N2499, N2498, N2497, N2496, N2495, N2494, N2493, N2492, N2491, N2490, N2489, N2488, N2487, N2486, N2485, N2484, N2483, N2482, N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471, N2470, N2469, N2468, N2467, N2466, N2465, N2464, N2463, N2462, N2461 } = (N45)? { N2460, N2459, N2458, N2457, N2456, N2455, N2454, N2453, N2452, N2451, N2450, N2449, N2448, N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, N2438, N2437, N2436, N2435, N2434, N2433, N2432, N2431, N2430, N2429, N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2396)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N45 = w_mask_i[29];
  assign { N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560, N2559, N2558, N2557, N2556, N2555, N2554, N2553, N2552, N2551, N2550, N2549, N2548, N2547, N2546, N2545, N2544, N2543, N2542, N2541, N2540, N2539, N2538, N2537, N2536, N2535, N2534, N2533, N2532, N2531, N2530, N2529, N2528, N2527, N2526 } = (N46)? { N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N6285, N3234, N3233, N3232, N3231, N2602, N2601, N2600, N3227, N4339, N4338, N4337, N4336, N2599, N2598, N2597, N3223, N4331, N4330, N4329, N4328, N2596, N2595, N2594, N3219, N4323, N4322, N4321, N4320, N2593, N2592, N2591, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2525)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N46 = w_mask_i[30];
  assign { N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, N2673, N2672, N2671, N2670, N2669, N2668, N2667, N2666, N2665, N2664, N2663, N2662, N2661, N2660, N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630 } = (N47)? { N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N6285, N3234, N3233, N3232, N3231, N2602, N2601, N2600, N3227, N4339, N4338, N4337, N4336, N2599, N2598, N2597, N3223, N4331, N4330, N4329, N4328, N2596, N2595, N2594, N3219, N4323, N4322, N4321, N4320, N2593, N2592, N2591, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2590)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N47 = w_mask_i[31];
  assign { N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, N2750, N2749, N2748, N2747, N2746, N2745, N2744, N2743, N2742, N2741, N2740, N2739, N2738, N2737, N2736, N2735, N2734, N2733, N2732, N2731, N2730, N2729, N2728, N2727, N2726, N2725, N2724, N2723, N2722, N2721, N2720, N2719, N2718, N2717, N2716, N2715, N2714, N2713, N2712, N2711, N2710, N2709, N2708, N2707, N2706, N2705, N2704, N2703, N2702, N2701, N2700, N2699, N2698, N2697, N2696, N2695 } = (N48)? { N3486, N3485, N3484, N3252, N3251, N3250, N3249, N3248, N3478, N3477, N3476, N3247, N3246, N3245, N3244, N3243, N3470, N3469, N3468, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N6285, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N4339, N4338, N4337, N4336, N3226, N3225, N3224, N3223, N4331, N4330, N4329, N4328, N3222, N3221, N3220, N3219, N4323, N4322, N4321, N4320, N3218, N3217, N3216, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2694)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N48 = w_mask_i[32];
  assign { N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N2806, N2805, N2804, N2803, N2802, N2801, N2800, N2799, N2798, N2797, N2796, N2795, N2794, N2793, N2792, N2791, N2790, N2789, N2788, N2787, N2786, N2785, N2784, N2783, N2782, N2781, N2780, N2779, N2778, N2777, N2776, N2775, N2774, N2773, N2772, N2771, N2770, N2769, N2768, N2767, N2766, N2765, N2764, N2763, N2762, N2761, N2760 } = (N49)? { N3486, N3485, N3484, N3252, N3251, N3250, N3249, N3248, N3478, N3477, N3476, N3247, N3246, N3245, N3244, N3243, N3470, N3469, N3468, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N6285, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N4339, N4338, N4337, N4336, N3226, N3225, N3224, N3223, N4331, N4330, N4329, N4328, N3222, N3221, N3220, N3219, N4323, N4322, N4321, N4320, N3218, N3217, N3216, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2759)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N49 = w_mask_i[33];
  assign { N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, N2878, N2877, N2876, N2875, N2874, N2873, N2872, N2871, N2870, N2869, N2868, N2867, N2866, N2865, N2864, N2863, N2862, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, N2848, N2847, N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838, N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, N2827, N2826, N2825 } = (N50)? { N3486, N3485, N3484, N3252, N3251, N3250, N3249, N3248, N3478, N3477, N3476, N3247, N3246, N3245, N3244, N3243, N3470, N3469, N3468, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N6285, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N4339, N4338, N4337, N4336, N3226, N3225, N3224, N3223, N4331, N4330, N4329, N4328, N3222, N3221, N3220, N3219, N4323, N4322, N4321, N4320, N3218, N3217, N3216, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2824)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N50 = w_mask_i[34];
  assign { N2953, N2952, N2951, N2950, N2949, N2948, N2947, N2946, N2945, N2944, N2943, N2942, N2941, N2940, N2939, N2938, N2937, N2936, N2935, N2934, N2933, N2932, N2931, N2930, N2929, N2928, N2927, N2926, N2925, N2924, N2923, N2922, N2921, N2920, N2919, N2918, N2917, N2916, N2915, N2914, N2913, N2912, N2911, N2910, N2909, N2908, N2907, N2906, N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898, N2897, N2896, N2895, N2894, N2893, N2892, N2891, N2890 } = (N51)? { N3486, N3485, N3484, N3252, N3251, N3250, N3249, N3248, N3478, N3477, N3476, N3247, N3246, N3245, N3244, N3243, N3470, N3469, N3468, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N6285, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N4339, N4338, N4337, N4336, N3226, N3225, N3224, N3223, N4331, N4330, N4329, N4328, N3222, N3221, N3220, N3219, N4323, N4322, N4321, N4320, N3218, N3217, N3216, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2889)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N51 = w_mask_i[35];
  assign { N3018, N3017, N3016, N3015, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N3007, N3006, N3005, N3004, N3003, N3002, N3001, N3000, N2999, N2998, N2997, N2996, N2995, N2994, N2993, N2992, N2991, N2990, N2989, N2988, N2987, N2986, N2985, N2984, N2983, N2982, N2981, N2980, N2979, N2978, N2977, N2976, N2975, N2974, N2973, N2972, N2971, N2970, N2969, N2968, N2967, N2966, N2965, N2964, N2963, N2962, N2961, N2960, N2959, N2958, N2957, N2956, N2955 } = (N52)? { N3486, N3485, N3484, N3252, N3251, N3250, N3249, N3248, N3478, N3477, N3476, N3247, N3246, N3245, N3244, N3243, N3470, N3469, N3468, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N6285, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N4339, N4338, N4337, N4336, N3226, N3225, N3224, N3223, N4331, N4330, N4329, N4328, N3222, N3221, N3220, N3219, N4323, N4322, N4321, N4320, N3218, N3217, N3216, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2954)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N52 = w_mask_i[36];
  assign { N3083, N3082, N3081, N3080, N3079, N3078, N3077, N3076, N3075, N3074, N3073, N3072, N3071, N3070, N3069, N3068, N3067, N3066, N3065, N3064, N3063, N3062, N3061, N3060, N3059, N3058, N3057, N3056, N3055, N3054, N3053, N3052, N3051, N3050, N3049, N3048, N3047, N3046, N3045, N3044, N3043, N3042, N3041, N3040, N3039, N3038, N3037, N3036, N3035, N3034, N3033, N3032, N3031, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N3023, N3022, N3021, N3020 } = (N53)? { N3486, N3485, N3484, N3252, N3251, N3250, N3249, N3248, N3478, N3477, N3476, N3247, N3246, N3245, N3244, N3243, N3470, N3469, N3468, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N6285, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N4339, N4338, N4337, N4336, N3226, N3225, N3224, N3223, N4331, N4330, N4329, N4328, N3222, N3221, N3220, N3219, N4323, N4322, N4321, N4320, N3218, N3217, N3216, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3019)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N53 = w_mask_i[37];
  assign { N3148, N3147, N3146, N3145, N3144, N3143, N3142, N3141, N3140, N3139, N3138, N3137, N3136, N3135, N3134, N3133, N3132, N3131, N3130, N3129, N3128, N3127, N3126, N3125, N3124, N3123, N3122, N3121, N3120, N3119, N3118, N3117, N3116, N3115, N3114, N3113, N3112, N3111, N3110, N3109, N3108, N3107, N3106, N3105, N3104, N3103, N3102, N3101, N3100, N3099, N3098, N3097, N3096, N3095, N3094, N3093, N3092, N3091, N3090, N3089, N3088, N3087, N3086, N3085 } = (N54)? { N3486, N3485, N3484, N3252, N3251, N3250, N3249, N3248, N3478, N3477, N3476, N3247, N3246, N3245, N3244, N3243, N3470, N3469, N3468, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N6285, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N4339, N4338, N4337, N4336, N3226, N3225, N3224, N3223, N4331, N4330, N4329, N4328, N3222, N3221, N3220, N3219, N4323, N4322, N4321, N4320, N3218, N3217, N3216, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3084)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N54 = w_mask_i[38];
  assign { N3213, N3212, N3211, N3210, N3209, N3208, N3207, N3206, N3205, N3204, N3203, N3202, N3201, N3200, N3199, N3198, N3197, N3196, N3195, N3194, N3193, N3192, N3191, N3190, N3189, N3188, N3187, N3186, N3185, N3184, N3183, N3182, N3181, N3180, N3179, N3178, N3177, N3176, N3175, N3174, N3173, N3172, N3171, N3170, N3169, N3168, N3167, N3166, N3165, N3164, N3163, N3162, N3161, N3160, N3159, N3158, N3157, N3156, N3155, N3154, N3153, N3152, N3151, N3150 } = (N55)? { N3486, N3485, N3484, N3252, N3251, N3250, N3249, N3248, N3478, N3477, N3476, N3247, N3246, N3245, N3244, N3243, N3470, N3469, N3468, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N6285, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N4339, N4338, N4337, N4336, N3226, N3225, N3224, N3223, N4331, N4330, N4329, N4328, N3222, N3221, N3220, N3219, N4323, N4322, N4321, N4320, N3218, N3217, N3216, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3149)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N55 = w_mask_i[39];
  assign { N3316, N3315, N3314, N3313, N3312, N3311, N3310, N3309, N3308, N3307, N3306, N3305, N3304, N3303, N3302, N3301, N3300, N3299, N3298, N3297, N3296, N3295, N3294, N3293, N3292, N3291, N3290, N3289, N3288, N3287, N3286, N3285, N3284, N3283, N3282, N3281, N3280, N3279, N3278, N3277, N3276, N3275, N3274, N3273, N3272, N3271, N3270, N3269, N3268, N3267, N3266, N3265, N3264, N3263, N3262, N3261, N3260, N3259, N3258, N3257, N3256, N3255, N3254, N3253 } = (N56)? { N3486, N3485, N3484, N3252, N3251, N3250, N3249, N3248, N3478, N3477, N3476, N3247, N3246, N3245, N3244, N3243, N3470, N3469, N3468, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N6285, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N4339, N4338, N4337, N4336, N3226, N3225, N3224, N3223, N4331, N4330, N4329, N4328, N3222, N3221, N3220, N3219, N4323, N4322, N4321, N4320, N3218, N3217, N3216, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3214)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N56 = w_mask_i[40];
  assign { N3381, N3380, N3379, N3378, N3377, N3376, N3375, N3374, N3373, N3372, N3371, N3370, N3369, N3368, N3367, N3366, N3365, N3364, N3363, N3362, N3361, N3360, N3359, N3358, N3357, N3356, N3355, N3354, N3353, N3352, N3351, N3350, N3349, N3348, N3347, N3346, N3345, N3344, N3343, N3342, N3341, N3340, N3339, N3338, N3337, N3336, N3335, N3334, N3333, N3332, N3331, N3330, N3329, N3328, N3327, N3326, N3325, N3324, N3323, N3322, N3321, N3320, N3319, N3318 } = (N57)? { N3486, N3485, N3484, N3483, N3482, N3481, N3480, N3479, N3478, N3477, N3476, N3475, N3474, N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N6165, N4014, N4013, N4012, N4011, N3459, N3458, N3457, N4010, N4226, N4225, N4224, N4223, N3456, N3455, N3454, N4009, N4218, N4217, N4216, N4215, N3453, N3452, N3451, N4008, N4210, N4209, N4208, N4207, N3450, N3449, N3448, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3317)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N57 = w_mask_i[41];
  assign { N3446, N3445, N3444, N3443, N3442, N3441, N3440, N3439, N3438, N3437, N3436, N3435, N3434, N3433, N3432, N3431, N3430, N3429, N3428, N3427, N3426, N3425, N3424, N3423, N3422, N3421, N3420, N3419, N3418, N3417, N3416, N3415, N3414, N3413, N3412, N3411, N3410, N3409, N3408, N3407, N3406, N3405, N3404, N3403, N3402, N3401, N3400, N3399, N3398, N3397, N3396, N3395, N3394, N3393, N3392, N3391, N3390, N3389, N3388, N3387, N3386, N3385, N3384, N3383 } = (N58)? { N3486, N3485, N3484, N3483, N3482, N3481, N3480, N3479, N3478, N3477, N3476, N3475, N3474, N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N6165, N4014, N4013, N4012, N4011, N3459, N3458, N3457, N4010, N4226, N4225, N4224, N4223, N3456, N3455, N3454, N4009, N4218, N4217, N4216, N4215, N3453, N3452, N3451, N4008, N4210, N4209, N4208, N4207, N3450, N3449, N3448, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3382)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N58 = w_mask_i[42];
  assign { N3550, N3549, N3548, N3547, N3546, N3545, N3544, N3543, N3542, N3541, N3540, N3539, N3538, N3537, N3536, N3535, N3534, N3533, N3532, N3531, N3530, N3529, N3528, N3527, N3526, N3525, N3524, N3523, N3522, N3521, N3520, N3519, N3518, N3517, N3516, N3515, N3514, N3513, N3512, N3511, N3510, N3509, N3508, N3507, N3506, N3505, N3504, N3503, N3502, N3501, N3500, N3499, N3498, N3497, N3496, N3495, N3494, N3493, N3492, N3491, N3490, N3489, N3488, N3487 } = (N59)? { N3486, N3485, N3484, N3483, N3482, N3481, N3480, N3479, N3478, N3477, N3476, N3475, N3474, N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N6165, N4014, N4013, N4012, N4011, N3459, N3458, N3457, N4010, N4226, N4225, N4224, N4223, N3456, N3455, N3454, N4009, N4218, N4217, N4216, N4215, N3453, N3452, N3451, N4008, N4210, N4209, N4208, N4207, N3450, N3449, N3448, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3447)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N59 = w_mask_i[43];
  assign { N3615, N3614, N3613, N3612, N3611, N3610, N3609, N3608, N3607, N3606, N3605, N3604, N3603, N3602, N3601, N3600, N3599, N3598, N3597, N3596, N3595, N3594, N3593, N3592, N3591, N3590, N3589, N3588, N3587, N3586, N3585, N3584, N3583, N3582, N3581, N3580, N3579, N3578, N3577, N3576, N3575, N3574, N3573, N3572, N3571, N3570, N3569, N3568, N3567, N3566, N3565, N3564, N3563, N3562, N3561, N3560, N3559, N3558, N3557, N3556, N3555, N3554, N3553, N3552 } = (N60)? { N4463, N4462, N4461, N4020, N4246, N4245, N4244, N4243, N4455, N4454, N4453, N4019, N4242, N4241, N4240, N4239, N4447, N4446, N4445, N4018, N4238, N4237, N4236, N4235, N4017, N4016, N4015, N6165, N4014, N4013, N4012, N4011, N4230, N4229, N4228, N4010, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4009, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4008, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3551)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N60 = w_mask_i[44];
  assign { N3680, N3679, N3678, N3677, N3676, N3675, N3674, N3673, N3672, N3671, N3670, N3669, N3668, N3667, N3666, N3665, N3664, N3663, N3662, N3661, N3660, N3659, N3658, N3657, N3656, N3655, N3654, N3653, N3652, N3651, N3650, N3649, N3648, N3647, N3646, N3645, N3644, N3643, N3642, N3641, N3640, N3639, N3638, N3637, N3636, N3635, N3634, N3633, N3632, N3631, N3630, N3629, N3628, N3627, N3626, N3625, N3624, N3623, N3622, N3621, N3620, N3619, N3618, N3617 } = (N61)? { N4463, N4462, N4461, N4020, N4246, N4245, N4244, N4243, N4455, N4454, N4453, N4019, N4242, N4241, N4240, N4239, N4447, N4446, N4445, N4018, N4238, N4237, N4236, N4235, N4017, N4016, N4015, N6165, N4014, N4013, N4012, N4011, N4230, N4229, N4228, N4010, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4009, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4008, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3616)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N61 = w_mask_i[45];
  assign { N3745, N3744, N3743, N3742, N3741, N3740, N3739, N3738, N3737, N3736, N3735, N3734, N3733, N3732, N3731, N3730, N3729, N3728, N3727, N3726, N3725, N3724, N3723, N3722, N3721, N3720, N3719, N3718, N3717, N3716, N3715, N3714, N3713, N3712, N3711, N3710, N3709, N3708, N3707, N3706, N3705, N3704, N3703, N3702, N3701, N3700, N3699, N3698, N3697, N3696, N3695, N3694, N3693, N3692, N3691, N3690, N3689, N3688, N3687, N3686, N3685, N3684, N3683, N3682 } = (N62)? { N4463, N4462, N4461, N4020, N4246, N4245, N4244, N4243, N4455, N4454, N4453, N4019, N4242, N4241, N4240, N4239, N4447, N4446, N4445, N4018, N4238, N4237, N4236, N4235, N4017, N4016, N4015, N6165, N4014, N4013, N4012, N4011, N4230, N4229, N4228, N4010, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4009, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4008, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3681)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N62 = w_mask_i[46];
  assign { N3810, N3809, N3808, N3807, N3806, N3805, N3804, N3803, N3802, N3801, N3800, N3799, N3798, N3797, N3796, N3795, N3794, N3793, N3792, N3791, N3790, N3789, N3788, N3787, N3786, N3785, N3784, N3783, N3782, N3781, N3780, N3779, N3778, N3777, N3776, N3775, N3774, N3773, N3772, N3771, N3770, N3769, N3768, N3767, N3766, N3765, N3764, N3763, N3762, N3761, N3760, N3759, N3758, N3757, N3756, N3755, N3754, N3753, N3752, N3751, N3750, N3749, N3748, N3747 } = (N63)? { N4463, N4462, N4461, N4020, N4246, N4245, N4244, N4243, N4455, N4454, N4453, N4019, N4242, N4241, N4240, N4239, N4447, N4446, N4445, N4018, N4238, N4237, N4236, N4235, N4017, N4016, N4015, N6165, N4014, N4013, N4012, N4011, N4230, N4229, N4228, N4010, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4009, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4008, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3746)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N63 = w_mask_i[47];
  assign { N3875, N3874, N3873, N3872, N3871, N3870, N3869, N3868, N3867, N3866, N3865, N3864, N3863, N3862, N3861, N3860, N3859, N3858, N3857, N3856, N3855, N3854, N3853, N3852, N3851, N3850, N3849, N3848, N3847, N3846, N3845, N3844, N3843, N3842, N3841, N3840, N3839, N3838, N3837, N3836, N3835, N3834, N3833, N3832, N3831, N3830, N3829, N3828, N3827, N3826, N3825, N3824, N3823, N3822, N3821, N3820, N3819, N3818, N3817, N3816, N3815, N3814, N3813, N3812 } = (N64)? { N4463, N4462, N4461, N4020, N4246, N4245, N4244, N4243, N4455, N4454, N4453, N4019, N4242, N4241, N4240, N4239, N4447, N4446, N4445, N4018, N4238, N4237, N4236, N4235, N4017, N4016, N4015, N6165, N4014, N4013, N4012, N4011, N4230, N4229, N4228, N4010, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4009, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4008, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3811)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N64 = w_mask_i[48];
  assign { N3940, N3939, N3938, N3937, N3936, N3935, N3934, N3933, N3932, N3931, N3930, N3929, N3928, N3927, N3926, N3925, N3924, N3923, N3922, N3921, N3920, N3919, N3918, N3917, N3916, N3915, N3914, N3913, N3912, N3911, N3910, N3909, N3908, N3907, N3906, N3905, N3904, N3903, N3902, N3901, N3900, N3899, N3898, N3897, N3896, N3895, N3894, N3893, N3892, N3891, N3890, N3889, N3888, N3887, N3886, N3885, N3884, N3883, N3882, N3881, N3880, N3879, N3878, N3877 } = (N65)? { N4463, N4462, N4461, N4020, N4246, N4245, N4244, N4243, N4455, N4454, N4453, N4019, N4242, N4241, N4240, N4239, N4447, N4446, N4445, N4018, N4238, N4237, N4236, N4235, N4017, N4016, N4015, N6165, N4014, N4013, N4012, N4011, N4230, N4229, N4228, N4010, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4009, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4008, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3876)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N65 = w_mask_i[49];
  assign { N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998, N3997, N3996, N3995, N3994, N3993, N3992, N3991, N3990, N3989, N3988, N3987, N3986, N3985, N3984, N3983, N3982, N3981, N3980, N3979, N3978, N3977, N3976, N3975, N3974, N3973, N3972, N3971, N3970, N3969, N3968, N3967, N3966, N3965, N3964, N3963, N3962, N3961, N3960, N3959, N3958, N3957, N3956, N3955, N3954, N3953, N3952, N3951, N3950, N3949, N3948, N3947, N3946, N3945, N3944, N3943, N3942 } = (N66)? { N4463, N4462, N4461, N4020, N4246, N4245, N4244, N4243, N4455, N4454, N4453, N4019, N4242, N4241, N4240, N4239, N4447, N4446, N4445, N4018, N4238, N4237, N4236, N4235, N4017, N4016, N4015, N6165, N4014, N4013, N4012, N4011, N4230, N4229, N4228, N4010, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4009, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4008, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3941)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N66 = w_mask_i[50];
  assign { N4084, N4083, N4082, N4081, N4080, N4079, N4078, N4077, N4076, N4075, N4074, N4073, N4072, N4071, N4070, N4069, N4068, N4067, N4066, N4065, N4064, N4063, N4062, N4061, N4060, N4059, N4058, N4057, N4056, N4055, N4054, N4053, N4052, N4051, N4050, N4049, N4048, N4047, N4046, N4045, N4044, N4043, N4042, N4041, N4040, N4039, N4038, N4037, N4036, N4035, N4034, N4033, N4032, N4031, N4030, N4029, N4028, N4027, N4026, N4025, N4024, N4023, N4022, N4021 } = (N67)? { N4463, N4462, N4461, N4020, N4246, N4245, N4244, N4243, N4455, N4454, N4453, N4019, N4242, N4241, N4240, N4239, N4447, N4446, N4445, N4018, N4238, N4237, N4236, N4235, N4017, N4016, N4015, N6165, N4014, N4013, N4012, N4011, N4230, N4229, N4228, N4010, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4009, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4008, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4006)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N67 = w_mask_i[51];
  assign { N4197, N4196, N4195, N4194, N4193, N4192, N4191, N4190, N4189, N4188, N4187, N4186, N4185, N4184, N4183, N4182, N4181, N4180, N4179, N4178, N4177, N4176, N4175, N4174, N4173, N4172, N4171, N4170, N4169, N4168, N4167, N4166, N4165, N4164, N4163, N4162, N4161, N4160, N4159, N4158, N4157, N4156, N4155, N4154, N4153, N4152, N4151, N4150, N4149, N4148, N4147, N4146, N4145, N4144, N4143, N4142, N4141, N4140, N4139, N4138, N4137, N4136, N4135, N4134 } = (N68)? { N4463, N4462, N4461, N4460, N4133, N4132, N4131, N4130, N4455, N4454, N4453, N4452, N4129, N4128, N4127, N4126, N4447, N4446, N4445, N4444, N4125, N4124, N4123, N4122, N4439, N4438, N4437, N6045, N4121, N4120, N4119, N4118, N4117, N4116, N4115, N4114, N4113, N4112, N4111, N4110, N4109, N4108, N4107, N4106, N4105, N4104, N4103, N4102, N4101, N4100, N4099, N4098, N4097, N4096, N4095, N4094, N4093, N4092, N4091, N4090, N4089, N4088, N4087, N4086 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4085)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N68 = w_mask_i[52];
  assign { N4310, N4309, N4308, N4307, N4306, N4305, N4304, N4303, N4302, N4301, N4300, N4299, N4298, N4297, N4296, N4295, N4294, N4293, N4292, N4291, N4290, N4289, N4288, N4287, N4286, N4285, N4284, N4283, N4282, N4281, N4280, N4279, N4278, N4277, N4276, N4275, N4274, N4273, N4272, N4271, N4270, N4269, N4268, N4267, N4266, N4265, N4264, N4263, N4262, N4261, N4260, N4259, N4258, N4257, N4256, N4255, N4254, N4253, N4252, N4251, N4250, N4249, N4248, N4247 } = (N69)? { N4463, N4462, N4461, N4460, N4246, N4245, N4244, N4243, N4455, N4454, N4453, N4452, N4242, N4241, N4240, N4239, N4447, N4446, N4445, N4444, N4238, N4237, N4236, N4235, N4439, N4438, N4437, N6045, N4234, N4233, N4232, N4231, N4230, N4229, N4228, N4227, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4219, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4211, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4203, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4198)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N69 = w_mask_i[53];
  assign { N4423, N4422, N4421, N4420, N4419, N4418, N4417, N4416, N4415, N4414, N4413, N4412, N4411, N4410, N4409, N4408, N4407, N4406, N4405, N4404, N4403, N4402, N4401, N4400, N4399, N4398, N4397, N4396, N4395, N4394, N4393, N4392, N4391, N4390, N4389, N4388, N4387, N4386, N4385, N4384, N4383, N4382, N4381, N4380, N4379, N4378, N4377, N4376, N4375, N4374, N4373, N4372, N4371, N4370, N4369, N4368, N4367, N4366, N4365, N4364, N4363, N4362, N4361, N4360 } = (N70)? { N4463, N4462, N4461, N4460, N4359, N4358, N4357, N4356, N4455, N4454, N4453, N4452, N4355, N4354, N4353, N4352, N4447, N4446, N4445, N4444, N4351, N4350, N4349, N4348, N4439, N4438, N4437, N6045, N4347, N4346, N4345, N4344, N4343, N4342, N4341, N4340, N4339, N4338, N4337, N4336, N4335, N4334, N4333, N4332, N4331, N4330, N4329, N4328, N4327, N4326, N4325, N4324, N4323, N4322, N4321, N4320, N4319, N4318, N4317, N4316, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4311)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N70 = w_mask_i[54];
  assign { N4527, N4526, N4525, N4524, N4523, N4522, N4521, N4520, N4519, N4518, N4517, N4516, N4515, N4514, N4513, N4512, N4511, N4510, N4509, N4508, N4507, N4506, N4505, N4504, N4503, N4502, N4501, N4500, N4499, N4498, N4497, N4496, N4495, N4494, N4493, N4492, N4491, N4490, N4489, N4488, N4487, N4486, N4485, N4484, N4483, N4482, N4481, N4480, N4479, N4478, N4477, N4476, N4475, N4474, N4473, N4472, N4471, N4470, N4469, N4468, N4467, N4466, N4465, N4464 } = (N71)? { N4463, N4462, N4461, N4460, N4459, N4458, N4457, N4456, N4455, N4454, N4453, N4452, N4451, N4450, N4449, N4448, N4447, N4446, N4445, N4444, N4443, N4442, N4441, N4440, N4439, N4438, N4437, N6045, N4926, N4925, N4924, N4923, N4436, N4435, N4434, N4922, N6276, N6275, N6274, N6273, N4433, N4432, N4431, N4921, N6268, N6267, N6266, N6265, N4430, N4429, N4428, N4920, N6260, N6259, N6258, N6257, N4427, N4426, N4425, N4919, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4424)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N71 = w_mask_i[55];
  assign { N4592, N4591, N4590, N4589, N4588, N4587, N4586, N4585, N4584, N4583, N4582, N4581, N4580, N4579, N4578, N4577, N4576, N4575, N4574, N4573, N4572, N4571, N4570, N4569, N4568, N4567, N4566, N4565, N4564, N4563, N4562, N4561, N4560, N4559, N4558, N4557, N4556, N4555, N4554, N4553, N4552, N4551, N4550, N4549, N4548, N4547, N4546, N4545, N4544, N4543, N4542, N4541, N4540, N4539, N4538, N4537, N4536, N4535, N4534, N4533, N4532, N4531, N4530, N4529 } = (N72)? { N5328, N5327, N5326, N4932, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N4931, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N4930, N5151, N5150, N5149, N5148, N4929, N4928, N4927, N6045, N4926, N4925, N4924, N4923, N5143, N5142, N5141, N4922, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N4921, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N4920, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N4919, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4528)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N72 = w_mask_i[56];
  assign { N4657, N4656, N4655, N4654, N4653, N4652, N4651, N4650, N4649, N4648, N4647, N4646, N4645, N4644, N4643, N4642, N4641, N4640, N4639, N4638, N4637, N4636, N4635, N4634, N4633, N4632, N4631, N4630, N4629, N4628, N4627, N4626, N4625, N4624, N4623, N4622, N4621, N4620, N4619, N4618, N4617, N4616, N4615, N4614, N4613, N4612, N4611, N4610, N4609, N4608, N4607, N4606, N4605, N4604, N4603, N4602, N4601, N4600, N4599, N4598, N4597, N4596, N4595, N4594 } = (N73)? { N5328, N5327, N5326, N4932, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N4931, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N4930, N5151, N5150, N5149, N5148, N4929, N4928, N4927, N6045, N4926, N4925, N4924, N4923, N5143, N5142, N5141, N4922, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N4921, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N4920, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N4919, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4593)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N73 = w_mask_i[57];
  assign { N4722, N4721, N4720, N4719, N4718, N4717, N4716, N4715, N4714, N4713, N4712, N4711, N4710, N4709, N4708, N4707, N4706, N4705, N4704, N4703, N4702, N4701, N4700, N4699, N4698, N4697, N4696, N4695, N4694, N4693, N4692, N4691, N4690, N4689, N4688, N4687, N4686, N4685, N4684, N4683, N4682, N4681, N4680, N4679, N4678, N4677, N4676, N4675, N4674, N4673, N4672, N4671, N4670, N4669, N4668, N4667, N4666, N4665, N4664, N4663, N4662, N4661, N4660, N4659 } = (N74)? { N5328, N5327, N5326, N4932, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N4931, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N4930, N5151, N5150, N5149, N5148, N4929, N4928, N4927, N6045, N4926, N4925, N4924, N4923, N5143, N5142, N5141, N4922, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N4921, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N4920, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N4919, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4658)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N74 = w_mask_i[58];
  assign { N4787, N4786, N4785, N4784, N4783, N4782, N4781, N4780, N4779, N4778, N4777, N4776, N4775, N4774, N4773, N4772, N4771, N4770, N4769, N4768, N4767, N4766, N4765, N4764, N4763, N4762, N4761, N4760, N4759, N4758, N4757, N4756, N4755, N4754, N4753, N4752, N4751, N4750, N4749, N4748, N4747, N4746, N4745, N4744, N4743, N4742, N4741, N4740, N4739, N4738, N4737, N4736, N4735, N4734, N4733, N4732, N4731, N4730, N4729, N4728, N4727, N4726, N4725, N4724 } = (N75)? { N5328, N5327, N5326, N4932, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N4931, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N4930, N5151, N5150, N5149, N5148, N4929, N4928, N4927, N6045, N4926, N4925, N4924, N4923, N5143, N5142, N5141, N4922, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N4921, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N4920, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N4919, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4723)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N75 = w_mask_i[59];
  assign { N4852, N4851, N4850, N4849, N4848, N4847, N4846, N4845, N4844, N4843, N4842, N4841, N4840, N4839, N4838, N4837, N4836, N4835, N4834, N4833, N4832, N4831, N4830, N4829, N4828, N4827, N4826, N4825, N4824, N4823, N4822, N4821, N4820, N4819, N4818, N4817, N4816, N4815, N4814, N4813, N4812, N4811, N4810, N4809, N4808, N4807, N4806, N4805, N4804, N4803, N4802, N4801, N4800, N4799, N4798, N4797, N4796, N4795, N4794, N4793, N4792, N4791, N4790, N4789 } = (N76)? { N5328, N5327, N5326, N4932, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N4931, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N4930, N5151, N5150, N5149, N5148, N4929, N4928, N4927, N6045, N4926, N4925, N4924, N4923, N5143, N5142, N5141, N4922, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N4921, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N4920, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N4919, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4788)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N76 = w_mask_i[60];
  assign { N4917, N4916, N4915, N4914, N4913, N4912, N4911, N4910, N4909, N4908, N4907, N4906, N4905, N4904, N4903, N4902, N4901, N4900, N4899, N4898, N4897, N4896, N4895, N4894, N4893, N4892, N4891, N4890, N4889, N4888, N4887, N4886, N4885, N4884, N4883, N4882, N4881, N4880, N4879, N4878, N4877, N4876, N4875, N4874, N4873, N4872, N4871, N4870, N4869, N4868, N4867, N4866, N4865, N4864, N4863, N4862, N4861, N4860, N4859, N4858, N4857, N4856, N4855, N4854 } = (N77)? { N5328, N5327, N5326, N4932, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N4931, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N4930, N5151, N5150, N5149, N5148, N4929, N4928, N4927, N6045, N4926, N4925, N4924, N4923, N5143, N5142, N5141, N4922, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N4921, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N4920, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N4919, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4853)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N77 = w_mask_i[61];
  assign { N4996, N4995, N4994, N4993, N4992, N4991, N4990, N4989, N4988, N4987, N4986, N4985, N4984, N4983, N4982, N4981, N4980, N4979, N4978, N4977, N4976, N4975, N4974, N4973, N4972, N4971, N4970, N4969, N4968, N4967, N4966, N4965, N4964, N4963, N4962, N4961, N4960, N4959, N4958, N4957, N4956, N4955, N4954, N4953, N4952, N4951, N4950, N4949, N4948, N4947, N4946, N4945, N4944, N4943, N4942, N4941, N4940, N4939, N4938, N4937, N4936, N4935, N4934, N4933 } = (N78)? { N5328, N5327, N5326, N4932, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N4931, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N4930, N5151, N5150, N5149, N5148, N4929, N4928, N4927, N6045, N4926, N4925, N4924, N4923, N5143, N5142, N5141, N4922, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N4921, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N4920, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N4919, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4918)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N78 = w_mask_i[62];
  assign { N5061, N5060, N5059, N5058, N5057, N5056, N5055, N5054, N5053, N5052, N5051, N5050, N5049, N5048, N5047, N5046, N5045, N5044, N5043, N5042, N5041, N5040, N5039, N5038, N5037, N5036, N5035, N5034, N5033, N5032, N5031, N5030, N5029, N5028, N5027, N5026, N5025, N5024, N5023, N5022, N5021, N5020, N5019, N5018, N5017, N5016, N5015, N5014, N5013, N5012, N5011, N5010, N5009, N5008, N5007, N5006, N5005, N5004, N5003, N5002, N5001, N5000, N4999, N4998 } = (N79)? { N5328, N5327, N5326, N5325, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N5317, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N5309, N5151, N5150, N5149, N5148, N5304, N5303, N5302, N5937, N5147, N5146, N5145, N5144, N5143, N5142, N5141, N5140, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N5136, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N5132, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N5128, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4997)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N79 = w_mask_i[63];
  assign { N5126, N5125, N5124, N5123, N5122, N5121, N5120, N5119, N5118, N5117, N5116, N5115, N5114, N5113, N5112, N5111, N5110, N5109, N5108, N5107, N5106, N5105, N5104, N5103, N5102, N5101, N5100, N5099, N5098, N5097, N5096, N5095, N5094, N5093, N5092, N5091, N5090, N5089, N5088, N5087, N5086, N5085, N5084, N5083, N5082, N5081, N5080, N5079, N5078, N5077, N5076, N5075, N5074, N5073, N5072, N5071, N5070, N5069, N5068, N5067, N5066, N5065, N5064, N5063 } = (N80)? { N5328, N5327, N5326, N5325, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N5317, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N5309, N5151, N5150, N5149, N5148, N5304, N5303, N5302, N5937, N5147, N5146, N5145, N5144, N5143, N5142, N5141, N5140, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N5136, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N5132, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N5128, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5062)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N80 = w_mask_i[64];
  assign { N5223, N5222, N5221, N5220, N5219, N5218, N5217, N5216, N5215, N5214, N5213, N5212, N5211, N5210, N5209, N5208, N5207, N5206, N5205, N5204, N5203, N5202, N5201, N5200, N5199, N5198, N5197, N5196, N5195, N5194, N5193, N5192, N5191, N5190, N5189, N5188, N5187, N5186, N5185, N5184, N5183, N5182, N5181, N5180, N5179, N5178, N5177, N5176, N5175, N5174, N5173, N5172, N5171, N5170, N5169, N5168, N5167, N5166, N5165, N5164, N5163, N5162, N5161, N5160 } = (N81)? { N5328, N5327, N5326, N5325, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N5317, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N5309, N5151, N5150, N5149, N5148, N5304, N5303, N5302, N5937, N5147, N5146, N5145, N5144, N5143, N5142, N5141, N5140, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N5136, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N5132, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N5128, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5127)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N81 = w_mask_i[65];
  assign { N5288, N5287, N5286, N5285, N5284, N5283, N5282, N5281, N5280, N5279, N5278, N5277, N5276, N5275, N5274, N5273, N5272, N5271, N5270, N5269, N5268, N5267, N5266, N5265, N5264, N5263, N5262, N5261, N5260, N5259, N5258, N5257, N5256, N5255, N5254, N5253, N5252, N5251, N5250, N5249, N5248, N5247, N5246, N5245, N5244, N5243, N5242, N5241, N5240, N5239, N5238, N5237, N5236, N5235, N5234, N5233, N5232, N5231, N5230, N5229, N5228, N5227, N5226, N5225 } = (N82)? { N5328, N5327, N5326, N5325, N5324, N5323, N5322, N5321, N5320, N5319, N5318, N5317, N5316, N5315, N5314, N5313, N5312, N5311, N5310, N5309, N5308, N5307, N5306, N5305, N5304, N5303, N5302, N5937, N5936, N5935, N5934, N5933, N5301, N5300, N5299, N5932, N6156, N6155, N6154, N6153, N5298, N5297, N5296, N5931, N6148, N6147, N6146, N6145, N5295, N5294, N5293, N5930, N6140, N6139, N6138, N6137, N5292, N5291, N5290, N5929, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5224)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N82 = w_mask_i[66];
  assign { N5392, N5391, N5390, N5389, N5388, N5387, N5386, N5385, N5384, N5383, N5382, N5381, N5380, N5379, N5378, N5377, N5376, N5375, N5374, N5373, N5372, N5371, N5370, N5369, N5368, N5367, N5366, N5365, N5364, N5363, N5362, N5361, N5360, N5359, N5358, N5357, N5356, N5355, N5354, N5353, N5352, N5351, N5350, N5349, N5348, N5347, N5346, N5345, N5344, N5343, N5342, N5341, N5340, N5339, N5338, N5337, N5336, N5335, N5334, N5333, N5332, N5331, N5330, N5329 } = (N83)? { N5328, N5327, N5326, N5325, N5324, N5323, N5322, N5321, N5320, N5319, N5318, N5317, N5316, N5315, N5314, N5313, N5312, N5311, N5310, N5309, N5308, N5307, N5306, N5305, N5304, N5303, N5302, N5937, N5936, N5935, N5934, N5933, N5301, N5300, N5299, N5932, N6156, N6155, N6154, N6153, N5298, N5297, N5296, N5931, N6148, N6147, N6146, N6145, N5295, N5294, N5293, N5930, N6140, N6139, N6138, N6137, N5292, N5291, N5290, N5929, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5289)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N83 = w_mask_i[67];
  assign { N5457, N5456, N5455, N5454, N5453, N5452, N5451, N5450, N5449, N5448, N5447, N5446, N5445, N5444, N5443, N5442, N5441, N5440, N5439, N5438, N5437, N5436, N5435, N5434, N5433, N5432, N5431, N5430, N5429, N5428, N5427, N5426, N5425, N5424, N5423, N5422, N5421, N5420, N5419, N5418, N5417, N5416, N5415, N5414, N5413, N5412, N5411, N5410, N5409, N5408, N5407, N5406, N5405, N5404, N5403, N5402, N5401, N5400, N5399, N5398, N5397, N5396, N5395, N5394 } = (N84)? { N6312, N6311, N6310, N5943, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N5942, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N5941, N6172, N6171, N6170, N6169, N5940, N5939, N5938, N5937, N5936, N5935, N5934, N5933, N6160, N6159, N6158, N5932, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N5931, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N5930, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N5929, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5393)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N84 = w_mask_i[68];
  assign { N5522, N5521, N5520, N5519, N5518, N5517, N5516, N5515, N5514, N5513, N5512, N5511, N5510, N5509, N5508, N5507, N5506, N5505, N5504, N5503, N5502, N5501, N5500, N5499, N5498, N5497, N5496, N5495, N5494, N5493, N5492, N5491, N5490, N5489, N5488, N5487, N5486, N5485, N5484, N5483, N5482, N5481, N5480, N5479, N5478, N5477, N5476, N5475, N5474, N5473, N5472, N5471, N5470, N5469, N5468, N5467, N5466, N5465, N5464, N5463, N5462, N5461, N5460, N5459 } = (N85)? { N6312, N6311, N6310, N5943, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N5942, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N5941, N6172, N6171, N6170, N6169, N5940, N5939, N5938, N5937, N5936, N5935, N5934, N5933, N6160, N6159, N6158, N5932, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N5931, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N5930, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N5929, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5458)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N85 = w_mask_i[69];
  assign { N5587, N5586, N5585, N5584, N5583, N5582, N5581, N5580, N5579, N5578, N5577, N5576, N5575, N5574, N5573, N5572, N5571, N5570, N5569, N5568, N5567, N5566, N5565, N5564, N5563, N5562, N5561, N5560, N5559, N5558, N5557, N5556, N5555, N5554, N5553, N5552, N5551, N5550, N5549, N5548, N5547, N5546, N5545, N5544, N5543, N5542, N5541, N5540, N5539, N5538, N5537, N5536, N5535, N5534, N5533, N5532, N5531, N5530, N5529, N5528, N5527, N5526, N5525, N5524 } = (N86)? { N6312, N6311, N6310, N5943, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N5942, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N5941, N6172, N6171, N6170, N6169, N5940, N5939, N5938, N5937, N5936, N5935, N5934, N5933, N6160, N6159, N6158, N5932, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N5931, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N5930, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N5929, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5523)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N86 = w_mask_i[70];
  assign { N5652, N5651, N5650, N5649, N5648, N5647, N5646, N5645, N5644, N5643, N5642, N5641, N5640, N5639, N5638, N5637, N5636, N5635, N5634, N5633, N5632, N5631, N5630, N5629, N5628, N5627, N5626, N5625, N5624, N5623, N5622, N5621, N5620, N5619, N5618, N5617, N5616, N5615, N5614, N5613, N5612, N5611, N5610, N5609, N5608, N5607, N5606, N5605, N5604, N5603, N5602, N5601, N5600, N5599, N5598, N5597, N5596, N5595, N5594, N5593, N5592, N5591, N5590, N5589 } = (N87)? { N6312, N6311, N6310, N5943, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N5942, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N5941, N6172, N6171, N6170, N6169, N5940, N5939, N5938, N5937, N5936, N5935, N5934, N5933, N6160, N6159, N6158, N5932, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N5931, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N5930, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N5929, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5588)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N87 = w_mask_i[71];
  assign { N5717, N5716, N5715, N5714, N5713, N5712, N5711, N5710, N5709, N5708, N5707, N5706, N5705, N5704, N5703, N5702, N5701, N5700, N5699, N5698, N5697, N5696, N5695, N5694, N5693, N5692, N5691, N5690, N5689, N5688, N5687, N5686, N5685, N5684, N5683, N5682, N5681, N5680, N5679, N5678, N5677, N5676, N5675, N5674, N5673, N5672, N5671, N5670, N5669, N5668, N5667, N5666, N5665, N5664, N5663, N5662, N5661, N5660, N5659, N5658, N5657, N5656, N5655, N5654 } = (N88)? { N6312, N6311, N6310, N5943, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N5942, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N5941, N6172, N6171, N6170, N6169, N5940, N5939, N5938, N5937, N5936, N5935, N5934, N5933, N6160, N6159, N6158, N5932, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N5931, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N5930, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N5929, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5653)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N88 = w_mask_i[72];
  assign { N5782, N5781, N5780, N5779, N5778, N5777, N5776, N5775, N5774, N5773, N5772, N5771, N5770, N5769, N5768, N5767, N5766, N5765, N5764, N5763, N5762, N5761, N5760, N5759, N5758, N5757, N5756, N5755, N5754, N5753, N5752, N5751, N5750, N5749, N5748, N5747, N5746, N5745, N5744, N5743, N5742, N5741, N5740, N5739, N5738, N5737, N5736, N5735, N5734, N5733, N5732, N5731, N5730, N5729, N5728, N5727, N5726, N5725, N5724, N5723, N5722, N5721, N5720, N5719 } = (N89)? { N6312, N6311, N6310, N5943, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N5942, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N5941, N6172, N6171, N6170, N6169, N5940, N5939, N5938, N5937, N5936, N5935, N5934, N5933, N6160, N6159, N6158, N5932, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N5931, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N5930, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N5929, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5718)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N89 = w_mask_i[73];
  assign { N5847, N5846, N5845, N5844, N5843, N5842, N5841, N5840, N5839, N5838, N5837, N5836, N5835, N5834, N5833, N5832, N5831, N5830, N5829, N5828, N5827, N5826, N5825, N5824, N5823, N5822, N5821, N5820, N5819, N5818, N5817, N5816, N5815, N5814, N5813, N5812, N5811, N5810, N5809, N5808, N5807, N5806, N5805, N5804, N5803, N5802, N5801, N5800, N5799, N5798, N5797, N5796, N5795, N5794, N5793, N5792, N5791, N5790, N5789, N5788, N5787, N5786, N5785, N5784 } = (N90)? { N6312, N6311, N6310, N5863, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N5862, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N5861, N6172, N6171, N6170, N6169, N5860, N5859, N5858, N5857, N5856, N5855, N5854, N5853, N6160, N6159, N6158, N5852, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N5851, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N5850, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N5849, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5783)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N90 = w_mask_i[74];
  assign { N5927, N5926, N5925, N5924, N5923, N5922, N5921, N5920, N5919, N5918, N5917, N5916, N5915, N5914, N5913, N5912, N5911, N5910, N5909, N5908, N5907, N5906, N5905, N5904, N5903, N5902, N5901, N5900, N5899, N5898, N5897, N5896, N5895, N5894, N5893, N5892, N5891, N5890, N5889, N5888, N5887, N5886, N5885, N5884, N5883, N5882, N5881, N5880, N5879, N5878, N5877, N5876, N5875, N5874, N5873, N5872, N5871, N5870, N5869, N5868, N5867, N5866, N5865, N5864 } = (N91)? { N6312, N6311, N6310, N5863, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N5862, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N5861, N6172, N6171, N6170, N6169, N5860, N5859, N5858, N5857, N5856, N5855, N5854, N5853, N6160, N6159, N6158, N5852, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N5851, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N5850, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N5849, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5848)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N91 = w_mask_i[75];
  assign { N6007, N6006, N6005, N6004, N6003, N6002, N6001, N6000, N5999, N5998, N5997, N5996, N5995, N5994, N5993, N5992, N5991, N5990, N5989, N5988, N5987, N5986, N5985, N5984, N5983, N5982, N5981, N5980, N5979, N5978, N5977, N5976, N5975, N5974, N5973, N5972, N5971, N5970, N5969, N5968, N5967, N5966, N5965, N5964, N5963, N5962, N5961, N5960, N5959, N5958, N5957, N5956, N5955, N5954, N5953, N5952, N5951, N5950, N5949, N5948, N5947, N5946, N5945, N5944 } = (N92)? { N6312, N6311, N6310, N5943, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N5942, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N5941, N6172, N6171, N6170, N6169, N5940, N5939, N5938, N5937, N5936, N5935, N5934, N5933, N6160, N6159, N6158, N5932, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N5931, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N5930, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N5929, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5928)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N92 = w_mask_i[76];
  assign { N6127, N6126, N6125, N6124, N6123, N6122, N6121, N6120, N6119, N6118, N6117, N6116, N6115, N6114, N6113, N6112, N6111, N6110, N6109, N6108, N6107, N6106, N6105, N6104, N6103, N6102, N6101, N6100, N6099, N6098, N6097, N6096, N6095, N6094, N6093, N6092, N6091, N6090, N6089, N6088, N6087, N6086, N6085, N6084, N6083, N6082, N6081, N6080, N6079, N6078, N6077, N6076, N6075, N6074, N6073, N6072, N6071, N6070, N6069, N6068, N6067, N6066, N6065, N6064 } = (N93)? { N6312, N6311, N6310, N6063, N6062, N6061, N6060, N6059, N6304, N6303, N6302, N6058, N6057, N6056, N6055, N6054, N6296, N6295, N6294, N6053, N6052, N6051, N6050, N6049, N6048, N6047, N6046, N6045, N6044, N6043, N6042, N6041, N6040, N6039, N6038, N6037, N6036, N6035, N6034, N6033, N6032, N6031, N6030, N6029, N6028, N6027, N6026, N6025, N6024, N6023, N6022, N6021, N6020, N6019, N6018, N6017, N6016, N6015, N6014, N6013, N6012, N6011, N6010, N6009 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6008)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N93 = w_mask_i[77];
  assign { N6247, N6246, N6245, N6244, N6243, N6242, N6241, N6240, N6239, N6238, N6237, N6236, N6235, N6234, N6233, N6232, N6231, N6230, N6229, N6228, N6227, N6226, N6225, N6224, N6223, N6222, N6221, N6220, N6219, N6218, N6217, N6216, N6215, N6214, N6213, N6212, N6211, N6210, N6209, N6208, N6207, N6206, N6205, N6204, N6203, N6202, N6201, N6200, N6199, N6198, N6197, N6196, N6195, N6194, N6193, N6192, N6191, N6190, N6189, N6188, N6187, N6186, N6185, N6184 } = (N94)? { N6312, N6311, N6310, N6183, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N6178, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N6173, N6172, N6171, N6170, N6169, N6168, N6167, N6166, N6165, N6164, N6163, N6162, N6161, N6160, N6159, N6158, N6157, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N6149, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N6141, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N6133, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6128)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N94 = w_mask_i[78];
  assign { N6376, N6375, N6374, N6373, N6372, N6371, N6370, N6369, N6368, N6367, N6366, N6365, N6364, N6363, N6362, N6361, N6360, N6359, N6358, N6357, N6356, N6355, N6354, N6353, N6352, N6351, N6350, N6349, N6348, N6347, N6346, N6345, N6344, N6343, N6342, N6341, N6340, N6339, N6338, N6337, N6336, N6335, N6334, N6333, N6332, N6331, N6330, N6329, N6328, N6327, N6326, N6325, N6324, N6323, N6322, N6321, N6320, N6319, N6318, N6317, N6316, N6315, N6314, N6313 } = (N95)? { N6312, N6311, N6310, N6309, N6308, N6307, N6306, N6305, N6304, N6303, N6302, N6301, N6300, N6299, N6298, N6297, N6296, N6295, N6294, N6293, N6292, N6291, N6290, N6289, N6288, N6287, N6286, N6285, N6284, N6283, N6282, N6281, N6280, N6279, N6278, N6277, N6276, N6275, N6274, N6273, N6272, N6271, N6270, N6269, N6268, N6267, N6266, N6265, N6264, N6263, N6262, N6261, N6260, N6259, N6258, N6257, N6256, N6255, N6254, N6253, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6248)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N95 = w_mask_i[79];
  assign { N11496, N11495, N11494, N11493, N11492, N11491, N11490, N11489, N11488, N11487, N11486, N11485, N11484, N11483, N11482, N11481, N11480, N11479, N11478, N11477, N11476, N11475, N11474, N11473, N11472, N11471, N11470, N11469, N11468, N11467, N11466, N11465, N11464, N11463, N11462, N11461, N11460, N11459, N11458, N11457, N11456, N11455, N11454, N11453, N11452, N11451, N11450, N11449, N11448, N11447, N11446, N11445, N11444, N11443, N11442, N11441, N11440, N11439, N11438, N11437, N11436, N11435, N11434, N11433, N11432, N11431, N11430, N11429, N11428, N11427, N11426, N11425, N11424, N11423, N11422, N11421, N11420, N11419, N11418, N11417, N11416, N11415, N11414, N11413, N11412, N11411, N11410, N11409, N11408, N11407, N11406, N11405, N11404, N11403, N11402, N11401, N11400, N11399, N11398, N11397, N11396, N11395, N11394, N11393, N11392, N11391, N11390, N11389, N11388, N11387, N11386, N11385, N11384, N11383, N11382, N11381, N11380, N11379, N11378, N11377, N11376, N11375, N11374, N11373, N11372, N11371, N11370, N11369, N11368, N11367, N11366, N11365, N11364, N11363, N11362, N11361, N11360, N11359, N11358, N11357, N11356, N11355, N11354, N11353, N11352, N11351, N11350, N11349, N11348, N11347, N11346, N11345, N11344, N11343, N11342, N11341, N11340, N11339, N11338, N11337, N11336, N11335, N11334, N11333, N11332, N11331, N11330, N11329, N11328, N11327, N11326, N11325, N11324, N11323, N11322, N11321, N11320, N11319, N11318, N11317, N11316, N11315, N11314, N11313, N11312, N11311, N11310, N11309, N11308, N11307, N11306, N11305, N11304, N11303, N11302, N11301, N11300, N11299, N11298, N11297, N11296, N11295, N11294, N11293, N11292, N11291, N11290, N11289, N11288, N11287, N11286, N11285, N11284, N11283, N11282, N11281, N11280, N11279, N11278, N11277, N11276, N11275, N11274, N11273, N11272, N11271, N11270, N11269, N11268, N11267, N11266, N11265, N11264, N11263, N11262, N11261, N11260, N11259, N11258, N11257, N11256, N11255, N11254, N11253, N11252, N11251, N11250, N11249, N11248, N11247, N11246, N11245, N11244, N11243, N11242, N11241, N11240, N11239, N11238, N11237, N11236, N11235, N11234, N11233, N11232, N11231, N11230, N11229, N11228, N11227, N11226, N11225, N11224, N11223, N11222, N11221, N11220, N11219, N11218, N11217, N11216, N11215, N11214, N11213, N11212, N11211, N11210, N11209, N11208, N11207, N11206, N11205, N11204, N11203, N11202, N11201, N11200, N11199, N11198, N11197, N11196, N11195, N11194, N11193, N11192, N11191, N11190, N11189, N11188, N11187, N11186, N11185, N11184, N11183, N11182, N11181, N11180, N11179, N11178, N11177, N11176, N11175, N11174, N11173, N11172, N11171, N11170, N11169, N11168, N11167, N11166, N11165, N11164, N11163, N11162, N11161, N11160, N11159, N11158, N11157, N11156, N11155, N11154, N11153, N11152, N11151, N11150, N11149, N11148, N11147, N11146, N11145, N11144, N11143, N11142, N11141, N11140, N11139, N11138, N11137, N11136, N11135, N11134, N11133, N11132, N11131, N11130, N11129, N11128, N11127, N11126, N11125, N11124, N11123, N11122, N11121, N11120, N11119, N11118, N11117, N11116, N11115, N11114, N11113, N11112, N11111, N11110, N11109, N11108, N11107, N11106, N11105, N11104, N11103, N11102, N11101, N11100, N11099, N11098, N11097, N11096, N11095, N11094, N11093, N11092, N11091, N11090, N11089, N11088, N11087, N11086, N11085, N11084, N11083, N11082, N11081, N11080, N11079, N11078, N11077, N11076, N11075, N11074, N11073, N11072, N11071, N11070, N11069, N11068, N11067, N11066, N11065, N11064, N11063, N11062, N11061, N11060, N11059, N11058, N11057, N11056, N11055, N11054, N11053, N11052, N11051, N11050, N11049, N11048, N11047, N11046, N11045, N11044, N11043, N11042, N11041, N11040, N11039, N11038, N11037, N11036, N11035, N11034, N11033, N11032, N11031, N11030, N11029, N11028, N11027, N11026, N11025, N11024, N11023, N11022, N11021, N11020, N11019, N11018, N11017, N11016, N11015, N11014, N11013, N11012, N11011, N11010, N11009, N11008, N11007, N11006, N11005, N11004, N11003, N11002, N11001, N11000, N10999, N10998, N10997, N10996, N10995, N10994, N10993, N10992, N10991, N10990, N10989, N10988, N10987, N10986, N10985, N10984, N10983, N10982, N10981, N10980, N10979, N10978, N10977, N10976, N10975, N10974, N10973, N10972, N10971, N10970, N10969, N10968, N10967, N10966, N10965, N10964, N10963, N10962, N10961, N10960, N10959, N10958, N10957, N10956, N10955, N10954, N10953, N10952, N10951, N10950, N10949, N10948, N10947, N10946, N10945, N10944, N10943, N10942, N10941, N10940, N10939, N10938, N10937, N10936, N10935, N10934, N10933, N10932, N10931, N10930, N10929, N10928, N10927, N10926, N10925, N10924, N10923, N10922, N10921, N10920, N10919, N10918, N10917, N10916, N10915, N10914, N10913, N10912, N10911, N10910, N10909, N10908, N10907, N10906, N10905, N10904, N10903, N10902, N10901, N10900, N10899, N10898, N10897, N10896, N10895, N10894, N10893, N10892, N10891, N10890, N10889, N10888, N10887, N10886, N10885, N10884, N10883, N10882, N10881, N10880, N10879, N10878, N10877, N10876, N10875, N10874, N10873, N10872, N10871, N10870, N10869, N10868, N10867, N10866, N10865, N10864, N10863, N10862, N10861, N10860, N10859, N10858, N10857, N10856, N10855, N10854, N10853, N10852, N10851, N10850, N10849, N10848, N10847, N10846, N10845, N10844, N10843, N10842, N10841, N10840, N10839, N10838, N10837, N10836, N10835, N10834, N10833, N10832, N10831, N10830, N10829, N10828, N10827, N10826, N10825, N10824, N10823, N10822, N10821, N10820, N10819, N10818, N10817, N10816, N10815, N10814, N10813, N10812, N10811, N10810, N10809, N10808, N10807, N10806, N10805, N10804, N10803, N10802, N10801, N10800, N10799, N10798, N10797, N10796, N10795, N10794, N10793, N10792, N10791, N10790, N10789, N10788, N10787, N10786, N10785, N10784, N10783, N10782, N10781, N10780, N10779, N10778, N10777, N10776, N10775, N10774, N10773, N10772, N10771, N10770, N10769, N10768, N10767, N10766, N10765, N10764, N10763, N10762, N10761, N10760, N10759, N10758, N10757, N10756, N10755, N10754, N10753, N10752, N10751, N10750, N10749, N10748, N10747, N10746, N10745, N10744, N10743, N10742, N10741, N10740, N10739, N10738, N10737, N10736, N10735, N10734, N10733, N10732, N10731, N10730, N10729, N10728, N10727, N10726, N10725, N10724, N10723, N10722, N10721, N10720, N10719, N10718, N10717, N10716, N10715, N10714, N10713, N10712, N10711, N10710, N10709, N10708, N10707, N10706, N10705, N10704, N10703, N10702, N10701, N10700, N10699, N10698, N10697, N10696, N10695, N10694, N10693, N10692, N10691, N10690, N10689, N10688, N10687, N10686, N10685, N10684, N10683, N10682, N10681, N10680, N10679, N10678, N10677, N10676, N10675, N10674, N10673, N10672, N10671, N10670, N10669, N10668, N10667, N10666, N10665, N10664, N10663, N10662, N10661, N10660, N10659, N10658, N10657, N10656, N10655, N10654, N10653, N10652, N10651, N10650, N10649, N10648, N10647, N10646, N10645, N10644, N10643, N10642, N10641, N10640, N10639, N10638, N10637, N10636, N10635, N10634, N10633, N10632, N10631, N10630, N10629, N10628, N10627, N10626, N10625, N10624, N10623, N10622, N10621, N10620, N10619, N10618, N10617, N10616, N10615, N10614, N10613, N10612, N10611, N10610, N10609, N10608, N10607, N10606, N10605, N10604, N10603, N10602, N10601, N10600, N10599, N10598, N10597, N10596, N10595, N10594, N10593, N10592, N10591, N10590, N10589, N10588, N10587, N10586, N10585, N10584, N10583, N10582, N10581, N10580, N10579, N10578, N10577, N10576, N10575, N10574, N10573, N10572, N10571, N10570, N10569, N10568, N10567, N10566, N10565, N10564, N10563, N10562, N10561, N10560, N10559, N10558, N10557, N10556, N10555, N10554, N10553, N10552, N10551, N10550, N10549, N10548, N10547, N10546, N10545, N10544, N10543, N10542, N10541, N10540, N10539, N10538, N10537, N10536, N10535, N10534, N10533, N10532, N10531, N10530, N10529, N10528, N10527, N10526, N10525, N10524, N10523, N10522, N10521, N10520, N10519, N10518, N10517, N10516, N10515, N10514, N10513, N10512, N10511, N10510, N10509, N10508, N10507, N10506, N10505, N10504, N10503, N10502, N10501, N10500, N10499, N10498, N10497, N10496, N10495, N10494, N10493, N10492, N10491, N10490, N10489, N10488, N10487, N10486, N10485, N10484, N10483, N10482, N10481, N10480, N10479, N10478, N10477, N10476, N10475, N10474, N10473, N10472, N10471, N10470, N10469, N10468, N10467, N10466, N10465, N10464, N10463, N10462, N10461, N10460, N10459, N10458, N10457, N10456, N10455, N10454, N10453, N10452, N10451, N10450, N10449, N10448, N10447, N10446, N10445, N10444, N10443, N10442, N10441, N10440, N10439, N10438, N10437, N10436, N10435, N10434, N10433, N10432, N10431, N10430, N10429, N10428, N10427, N10426, N10425, N10424, N10423, N10422, N10421, N10420, N10419, N10418, N10417, N10416, N10415, N10414, N10413, N10412, N10411, N10410, N10409, N10408, N10407, N10406, N10405, N10404, N10403, N10402, N10401, N10400, N10399, N10398, N10397, N10396, N10395, N10394, N10393, N10392, N10391, N10390, N10389, N10388, N10387, N10386, N10385, N10384, N10383, N10382, N10381, N10380, N10379, N10378, N10377, N10376, N10375, N10374, N10373, N10372, N10371, N10370, N10369, N10368, N10367, N10366, N10365, N10364, N10363, N10362, N10361, N10360, N10359, N10358, N10357, N10356, N10355, N10354, N10353, N10352, N10351, N10350, N10349, N10348, N10347, N10346, N10345, N10344, N10343, N10342, N10341, N10340, N10339, N10338, N10337, N10336, N10335, N10334, N10333, N10332, N10331, N10330, N10329, N10328, N10327, N10326, N10325, N10324, N10323, N10322, N10321, N10320, N10319, N10318, N10317, N10316, N10315, N10314, N10313, N10312, N10311, N10310, N10309, N10308, N10307, N10306, N10305, N10304, N10303, N10302, N10301, N10300, N10299, N10298, N10297, N10296, N10295, N10294, N10293, N10292, N10291, N10290, N10289, N10288, N10287, N10286, N10285, N10284, N10283, N10282, N10281, N10280, N10279, N10278, N10277, N10276, N10275, N10274, N10273, N10272, N10271, N10270, N10269, N10268, N10267, N10266, N10265, N10264, N10263, N10262, N10261, N10260, N10259, N10258, N10257, N10256, N10255, N10254, N10253, N10252, N10251, N10250, N10249, N10248, N10247, N10246, N10245, N10244, N10243, N10242, N10241, N10240, N10239, N10238, N10237, N10236, N10235, N10234, N10233, N10232, N10231, N10230, N10229, N10228, N10227, N10226, N10225, N10224, N10223, N10222, N10221, N10220, N10219, N10218, N10217, N10216, N10215, N10214, N10213, N10212, N10211, N10210, N10209, N10208, N10207, N10206, N10205, N10204, N10203, N10202, N10201, N10200, N10199, N10198, N10197, N10196, N10195, N10194, N10193, N10192, N10191, N10190, N10189, N10188, N10187, N10186, N10185, N10184, N10183, N10182, N10181, N10180, N10179, N10178, N10177, N10176, N10175, N10174, N10173, N10172, N10171, N10170, N10169, N10168, N10167, N10166, N10165, N10164, N10163, N10162, N10161, N10160, N10159, N10158, N10157, N10156, N10155, N10154, N10153, N10152, N10151, N10150, N10149, N10148, N10147, N10146, N10145, N10144, N10143, N10142, N10141, N10140, N10139, N10138, N10137, N10136, N10135, N10134, N10133, N10132, N10131, N10130, N10129, N10128, N10127, N10126, N10125, N10124, N10123, N10122, N10121, N10120, N10119, N10118, N10117, N10116, N10115, N10114, N10113, N10112, N10111, N10110, N10109, N10108, N10107, N10106, N10105, N10104, N10103, N10102, N10101, N10100, N10099, N10098, N10097, N10096, N10095, N10094, N10093, N10092, N10091, N10090, N10089, N10088, N10087, N10086, N10085, N10084, N10083, N10082, N10081, N10080, N10079, N10078, N10077, N10076, N10075, N10074, N10073, N10072, N10071, N10070, N10069, N10068, N10067, N10066, N10065, N10064, N10063, N10062, N10061, N10060, N10059, N10058, N10057, N10056, N10055, N10054, N10053, N10052, N10051, N10050, N10049, N10048, N10047, N10046, N10045, N10044, N10043, N10042, N10041, N10040, N10039, N10038, N10037, N10036, N10035, N10034, N10033, N10032, N10031, N10030, N10029, N10028, N10027, N10026, N10025, N10024, N10023, N10022, N10021, N10020, N10019, N10018, N10017, N10016, N10015, N10014, N10013, N10012, N10011, N10010, N10009, N10008, N10007, N10006, N10005, N10004, N10003, N10002, N10001, N10000, N9999, N9998, N9997, N9996, N9995, N9994, N9993, N9992, N9991, N9990, N9989, N9988, N9987, N9986, N9985, N9984, N9983, N9982, N9981, N9980, N9979, N9978, N9977, N9976, N9975, N9974, N9973, N9972, N9971, N9970, N9969, N9968, N9967, N9966, N9965, N9964, N9963, N9962, N9961, N9960, N9959, N9958, N9957, N9956, N9955, N9954, N9953, N9952, N9951, N9950, N9949, N9948, N9947, N9946, N9945, N9944, N9943, N9942, N9941, N9940, N9939, N9938, N9937, N9936, N9935, N9934, N9933, N9932, N9931, N9930, N9929, N9928, N9927, N9926, N9925, N9924, N9923, N9922, N9921, N9920, N9919, N9918, N9917, N9916, N9915, N9914, N9913, N9912, N9911, N9910, N9909, N9908, N9907, N9906, N9905, N9904, N9903, N9902, N9901, N9900, N9899, N9898, N9897, N9896, N9895, N9894, N9893, N9892, N9891, N9890, N9889, N9888, N9887, N9886, N9885, N9884, N9883, N9882, N9881, N9880, N9879, N9878, N9877, N9876, N9875, N9874, N9873, N9872, N9871, N9870, N9869, N9868, N9867, N9866, N9865, N9864, N9863, N9862, N9861, N9860, N9859, N9858, N9857, N9856, N9855, N9854, N9853, N9852, N9851, N9850, N9849, N9848, N9847, N9846, N9845, N9844, N9843, N9842, N9841, N9840, N9839, N9838, N9837, N9836, N9835, N9834, N9833, N9832, N9831, N9830, N9829, N9828, N9827, N9826, N9825, N9824, N9823, N9822, N9821, N9820, N9819, N9818, N9817, N9816, N9815, N9814, N9813, N9812, N9811, N9810, N9809, N9808, N9807, N9806, N9805, N9804, N9803, N9802, N9801, N9800, N9799, N9798, N9797, N9796, N9795, N9794, N9793, N9792, N9791, N9790, N9789, N9788, N9787, N9786, N9785, N9784, N9783, N9782, N9781, N9780, N9779, N9778, N9777, N9776, N9775, N9774, N9773, N9772, N9771, N9770, N9769, N9768, N9767, N9766, N9765, N9764, N9763, N9762, N9761, N9760, N9759, N9758, N9757, N9756, N9755, N9754, N9753, N9752, N9751, N9750, N9749, N9748, N9747, N9746, N9745, N9744, N9743, N9742, N9741, N9740, N9739, N9738, N9737, N9736, N9735, N9734, N9733, N9732, N9731, N9730, N9729, N9728, N9727, N9726, N9725, N9724, N9723, N9722, N9721, N9720, N9719, N9718, N9717, N9716, N9715, N9714, N9713, N9712, N9711, N9710, N9709, N9708, N9707, N9706, N9705, N9704, N9703, N9702, N9701, N9700, N9699, N9698, N9697, N9696, N9695, N9694, N9693, N9692, N9691, N9690, N9689, N9688, N9687, N9686, N9685, N9684, N9683, N9682, N9681, N9680, N9679, N9678, N9677, N9676, N9675, N9674, N9673, N9672, N9671, N9670, N9669, N9668, N9667, N9666, N9665, N9664, N9663, N9662, N9661, N9660, N9659, N9658, N9657, N9656, N9655, N9654, N9653, N9652, N9651, N9650, N9649, N9648, N9647, N9646, N9645, N9644, N9643, N9642, N9641, N9640, N9639, N9638, N9637, N9636, N9635, N9634, N9633, N9632, N9631, N9630, N9629, N9628, N9627, N9626, N9625, N9624, N9623, N9622, N9621, N9620, N9619, N9618, N9617, N9616, N9615, N9614, N9613, N9612, N9611, N9610, N9609, N9608, N9607, N9606, N9605, N9604, N9603, N9602, N9601, N9600, N9599, N9598, N9597, N9596, N9595, N9594, N9593, N9592, N9591, N9590, N9589, N9588, N9587, N9586, N9585, N9584, N9583, N9582, N9581, N9580, N9579, N9578, N9577, N9576, N9575, N9574, N9573, N9572, N9571, N9570, N9569, N9568, N9567, N9566, N9565, N9564, N9563, N9562, N9561, N9560, N9559, N9558, N9557, N9556, N9555, N9554, N9553, N9552, N9551, N9550, N9549, N9548, N9547, N9546, N9545, N9544, N9543, N9542, N9541, N9540, N9539, N9538, N9537, N9536, N9535, N9534, N9533, N9532, N9531, N9530, N9529, N9528, N9527, N9526, N9525, N9524, N9523, N9522, N9521, N9520, N9519, N9518, N9517, N9516, N9515, N9514, N9513, N9512, N9511, N9510, N9509, N9508, N9507, N9506, N9505, N9504, N9503, N9502, N9501, N9500, N9499, N9498, N9497, N9496, N9495, N9494, N9493, N9492, N9491, N9490, N9489, N9488, N9487, N9486, N9485, N9484, N9483, N9482, N9481, N9480, N9479, N9478, N9477, N9476, N9475, N9474, N9473, N9472, N9471, N9470, N9469, N9468, N9467, N9466, N9465, N9464, N9463, N9462, N9461, N9460, N9459, N9458, N9457, N9456, N9455, N9454, N9453, N9452, N9451, N9450, N9449, N9448, N9447, N9446, N9445, N9444, N9443, N9442, N9441, N9440, N9439, N9438, N9437, N9436, N9435, N9434, N9433, N9432, N9431, N9430, N9429, N9428, N9427, N9426, N9425, N9424, N9423, N9422, N9421, N9420, N9419, N9418, N9417, N9416, N9415, N9414, N9413, N9412, N9411, N9410, N9409, N9408, N9407, N9406, N9405, N9404, N9403, N9402, N9401, N9400, N9399, N9398, N9397, N9396, N9395, N9394, N9393, N9392, N9391, N9390, N9389, N9388, N9387, N9386, N9385, N9384, N9383, N9382, N9381, N9380, N9379, N9378, N9377, N9376, N9375, N9374, N9373, N9372, N9371, N9370, N9369, N9368, N9367, N9366, N9365, N9364, N9363, N9362, N9361, N9360, N9359, N9358, N9357, N9356, N9355, N9354, N9353, N9352, N9351, N9350, N9349, N9348, N9347, N9346, N9345, N9344, N9343, N9342, N9341, N9340, N9339, N9338, N9337, N9336, N9335, N9334, N9333, N9332, N9331, N9330, N9329, N9328, N9327, N9326, N9325, N9324, N9323, N9322, N9321, N9320, N9319, N9318, N9317, N9316, N9315, N9314, N9313, N9312, N9311, N9310, N9309, N9308, N9307, N9306, N9305, N9304, N9303, N9302, N9301, N9300, N9299, N9298, N9297, N9296, N9295, N9294, N9293, N9292, N9291, N9290, N9289, N9288, N9287, N9286, N9285, N9284, N9283, N9282, N9281, N9280, N9279, N9278, N9277, N9276, N9275, N9274, N9273, N9272, N9271, N9270, N9269, N9268, N9267, N9266, N9265, N9264, N9263, N9262, N9261, N9260, N9259, N9258, N9257, N9256, N9255, N9254, N9253, N9252, N9251, N9250, N9249, N9248, N9247, N9246, N9245, N9244, N9243, N9242, N9241, N9240, N9239, N9238, N9237, N9236, N9235, N9234, N9233, N9232, N9231, N9230, N9229, N9228, N9227, N9226, N9225, N9224, N9223, N9222, N9221, N9220, N9219, N9218, N9217, N9216, N9215, N9214, N9213, N9212, N9211, N9210, N9209, N9208, N9207, N9206, N9205, N9204, N9203, N9202, N9201, N9200, N9199, N9198, N9197, N9196, N9195, N9194, N9193, N9192, N9191, N9190, N9189, N9188, N9187, N9186, N9185, N9184, N9183, N9182, N9181, N9180, N9179, N9178, N9177, N9176, N9175, N9174, N9173, N9172, N9171, N9170, N9169, N9168, N9167, N9166, N9165, N9164, N9163, N9162, N9161, N9160, N9159, N9158, N9157, N9156, N9155, N9154, N9153, N9152, N9151, N9150, N9149, N9148, N9147, N9146, N9145, N9144, N9143, N9142, N9141, N9140, N9139, N9138, N9137, N9136, N9135, N9134, N9133, N9132, N9131, N9130, N9129, N9128, N9127, N9126, N9125, N9124, N9123, N9122, N9121, N9120, N9119, N9118, N9117, N9116, N9115, N9114, N9113, N9112, N9111, N9110, N9109, N9108, N9107, N9106, N9105, N9104, N9103, N9102, N9101, N9100, N9099, N9098, N9097, N9096, N9095, N9094, N9093, N9092, N9091, N9090, N9089, N9088, N9087, N9086, N9085, N9084, N9083, N9082, N9081, N9080, N9079, N9078, N9077, N9076, N9075, N9074, N9073, N9072, N9071, N9070, N9069, N9068, N9067, N9066, N9065, N9064, N9063, N9062, N9061, N9060, N9059, N9058, N9057, N9056, N9055, N9054, N9053, N9052, N9051, N9050, N9049, N9048, N9047, N9046, N9045, N9044, N9043, N9042, N9041, N9040, N9039, N9038, N9037, N9036, N9035, N9034, N9033, N9032, N9031, N9030, N9029, N9028, N9027, N9026, N9025, N9024, N9023, N9022, N9021, N9020, N9019, N9018, N9017, N9016, N9015, N9014, N9013, N9012, N9011, N9010, N9009, N9008, N9007, N9006, N9005, N9004, N9003, N9002, N9001, N9000, N8999, N8998, N8997, N8996, N8995, N8994, N8993, N8992, N8991, N8990, N8989, N8988, N8987, N8986, N8985, N8984, N8983, N8982, N8981, N8980, N8979, N8978, N8977, N8976, N8975, N8974, N8973, N8972, N8971, N8970, N8969, N8968, N8967, N8966, N8965, N8964, N8963, N8962, N8961, N8960, N8959, N8958, N8957, N8956, N8955, N8954, N8953, N8952, N8951, N8950, N8949, N8948, N8947, N8946, N8945, N8944, N8943, N8942, N8941, N8940, N8939, N8938, N8937, N8936, N8935, N8934, N8933, N8932, N8931, N8930, N8929, N8928, N8927, N8926, N8925, N8924, N8923, N8922, N8921, N8920, N8919, N8918, N8917, N8916, N8915, N8914, N8913, N8912, N8911, N8910, N8909, N8908, N8907, N8906, N8905, N8904, N8903, N8902, N8901, N8900, N8899, N8898, N8897, N8896, N8895, N8894, N8893, N8892, N8891, N8890, N8889, N8888, N8887, N8886, N8885, N8884, N8883, N8882, N8881, N8880, N8879, N8878, N8877, N8876, N8875, N8874, N8873, N8872, N8871, N8870, N8869, N8868, N8867, N8866, N8865, N8864, N8863, N8862, N8861, N8860, N8859, N8858, N8857, N8856, N8855, N8854, N8853, N8852, N8851, N8850, N8849, N8848, N8847, N8846, N8845, N8844, N8843, N8842, N8841, N8840, N8839, N8838, N8837, N8836, N8835, N8834, N8833, N8832, N8831, N8830, N8829, N8828, N8827, N8826, N8825, N8824, N8823, N8822, N8821, N8820, N8819, N8818, N8817, N8816, N8815, N8814, N8813, N8812, N8811, N8810, N8809, N8808, N8807, N8806, N8805, N8804, N8803, N8802, N8801, N8800, N8799, N8798, N8797, N8796, N8795, N8794, N8793, N8792, N8791, N8790, N8789, N8788, N8787, N8786, N8785, N8784, N8783, N8782, N8781, N8780, N8779, N8778, N8777, N8776, N8775, N8774, N8773, N8772, N8771, N8770, N8769, N8768, N8767, N8766, N8765, N8764, N8763, N8762, N8761, N8760, N8759, N8758, N8757, N8756, N8755, N8754, N8753, N8752, N8751, N8750, N8749, N8748, N8747, N8746, N8745, N8744, N8743, N8742, N8741, N8740, N8739, N8738, N8737, N8736, N8735, N8734, N8733, N8732, N8731, N8730, N8729, N8728, N8727, N8726, N8725, N8724, N8723, N8722, N8721, N8720, N8719, N8718, N8717, N8716, N8715, N8714, N8713, N8712, N8711, N8710, N8709, N8708, N8707, N8706, N8705, N8704, N8703, N8702, N8701, N8700, N8699, N8698, N8697, N8696, N8695, N8694, N8693, N8692, N8691, N8690, N8689, N8688, N8687, N8686, N8685, N8684, N8683, N8682, N8681, N8680, N8679, N8678, N8677, N8676, N8675, N8674, N8673, N8672, N8671, N8670, N8669, N8668, N8667, N8666, N8665, N8664, N8663, N8662, N8661, N8660, N8659, N8658, N8657, N8656, N8655, N8654, N8653, N8652, N8651, N8650, N8649, N8648, N8647, N8646, N8645, N8644, N8643, N8642, N8641, N8640, N8639, N8638, N8637, N8636, N8635, N8634, N8633, N8632, N8631, N8630, N8629, N8628, N8627, N8626, N8625, N8624, N8623, N8622, N8621, N8620, N8619, N8618, N8617, N8616, N8615, N8614, N8613, N8612, N8611, N8610, N8609, N8608, N8607, N8606, N8605, N8604, N8603, N8602, N8601, N8600, N8599, N8598, N8597, N8596, N8595, N8594, N8593, N8592, N8591, N8590, N8589, N8588, N8587, N8586, N8585, N8584, N8583, N8582, N8581, N8580, N8579, N8578, N8577, N8576, N8575, N8574, N8573, N8572, N8571, N8570, N8569, N8568, N8567, N8566, N8565, N8564, N8563, N8562, N8561, N8560, N8559, N8558, N8557, N8556, N8555, N8554, N8553, N8552, N8551, N8550, N8549, N8548, N8547, N8546, N8545, N8544, N8543, N8542, N8541, N8540, N8539, N8538, N8537, N8536, N8535, N8534, N8533, N8532, N8531, N8530, N8529, N8528, N8527, N8526, N8525, N8524, N8523, N8522, N8521, N8520, N8519, N8518, N8517, N8516, N8515, N8514, N8513, N8512, N8511, N8510, N8509, N8508, N8507, N8506, N8505, N8504, N8503, N8502, N8501, N8500, N8499, N8498, N8497, N8496, N8495, N8494, N8493, N8492, N8491, N8490, N8489, N8488, N8487, N8486, N8485, N8484, N8483, N8482, N8481, N8480, N8479, N8478, N8477, N8476, N8475, N8474, N8473, N8472, N8471, N8470, N8469, N8468, N8467, N8466, N8465, N8464, N8463, N8462, N8461, N8460, N8459, N8458, N8457, N8456, N8455, N8454, N8453, N8452, N8451, N8450, N8449, N8448, N8447, N8446, N8445, N8444, N8443, N8442, N8441, N8440, N8439, N8438, N8437, N8436, N8435, N8434, N8433, N8432, N8431, N8430, N8429, N8428, N8427, N8426, N8425, N8424, N8423, N8422, N8421, N8420, N8419, N8418, N8417, N8416, N8415, N8414, N8413, N8412, N8411, N8410, N8409, N8408, N8407, N8406, N8405, N8404, N8403, N8402, N8401, N8400, N8399, N8398, N8397, N8396, N8395, N8394, N8393, N8392, N8391, N8390, N8389, N8388, N8387, N8386, N8385, N8384, N8383, N8382, N8381, N8380, N8379, N8378, N8377, N8376, N8375, N8374, N8373, N8372, N8371, N8370, N8369, N8368, N8367, N8366, N8365, N8364, N8363, N8362, N8361, N8360, N8359, N8358, N8357, N8356, N8355, N8354, N8353, N8352, N8351, N8350, N8349, N8348, N8347, N8346, N8345, N8344, N8343, N8342, N8341, N8340, N8339, N8338, N8337, N8336, N8335, N8334, N8333, N8332, N8331, N8330, N8329, N8328, N8327, N8326, N8325, N8324, N8323, N8322, N8321, N8320, N8319, N8318, N8317, N8316, N8315, N8314, N8313, N8312, N8311, N8310, N8309, N8308, N8307, N8306, N8305, N8304, N8303, N8302, N8301, N8300, N8299, N8298, N8297, N8296, N8295, N8294, N8293, N8292, N8291, N8290, N8289, N8288, N8287, N8286, N8285, N8284, N8283, N8282, N8281, N8280, N8279, N8278, N8277, N8276, N8275, N8274, N8273, N8272, N8271, N8270, N8269, N8268, N8267, N8266, N8265, N8264, N8263, N8262, N8261, N8260, N8259, N8258, N8257, N8256, N8255, N8254, N8253, N8252, N8251, N8250, N8249, N8248, N8247, N8246, N8245, N8244, N8243, N8242, N8241, N8240, N8239, N8238, N8237, N8236, N8235, N8234, N8233, N8232, N8231, N8230, N8229, N8228, N8227, N8226, N8225, N8224, N8223, N8222, N8221, N8220, N8219, N8218, N8217, N8216, N8215, N8214, N8213, N8212, N8211, N8210, N8209, N8208, N8207, N8206, N8205, N8204, N8203, N8202, N8201, N8200, N8199, N8198, N8197, N8196, N8195, N8194, N8193, N8192, N8191, N8190, N8189, N8188, N8187, N8186, N8185, N8184, N8183, N8182, N8181, N8180, N8179, N8178, N8177, N8176, N8175, N8174, N8173, N8172, N8171, N8170, N8169, N8168, N8167, N8166, N8165, N8164, N8163, N8162, N8161, N8160, N8159, N8158, N8157, N8156, N8155, N8154, N8153, N8152, N8151, N8150, N8149, N8148, N8147, N8146, N8145, N8144, N8143, N8142, N8141, N8140, N8139, N8138, N8137, N8136, N8135, N8134, N8133, N8132, N8131, N8130, N8129, N8128, N8127, N8126, N8125, N8124, N8123, N8122, N8121, N8120, N8119, N8118, N8117, N8116, N8115, N8114, N8113, N8112, N8111, N8110, N8109, N8108, N8107, N8106, N8105, N8104, N8103, N8102, N8101, N8100, N8099, N8098, N8097, N8096, N8095, N8094, N8093, N8092, N8091, N8090, N8089, N8088, N8087, N8086, N8085, N8084, N8083, N8082, N8081, N8080, N8079, N8078, N8077, N8076, N8075, N8074, N8073, N8072, N8071, N8070, N8069, N8068, N8067, N8066, N8065, N8064, N8063, N8062, N8061, N8060, N8059, N8058, N8057, N8056, N8055, N8054, N8053, N8052, N8051, N8050, N8049, N8048, N8047, N8046, N8045, N8044, N8043, N8042, N8041, N8040, N8039, N8038, N8037, N8036, N8035, N8034, N8033, N8032, N8031, N8030, N8029, N8028, N8027, N8026, N8025, N8024, N8023, N8022, N8021, N8020, N8019, N8018, N8017, N8016, N8015, N8014, N8013, N8012, N8011, N8010, N8009, N8008, N8007, N8006, N8005, N8004, N8003, N8002, N8001, N8000, N7999, N7998, N7997, N7996, N7995, N7994, N7993, N7992, N7991, N7990, N7989, N7988, N7987, N7986, N7985, N7984, N7983, N7982, N7981, N7980, N7979, N7978, N7977, N7976, N7975, N7974, N7973, N7972, N7971, N7970, N7969, N7968, N7967, N7966, N7965, N7964, N7963, N7962, N7961, N7960, N7959, N7958, N7957, N7956, N7955, N7954, N7953, N7952, N7951, N7950, N7949, N7948, N7947, N7946, N7945, N7944, N7943, N7942, N7941, N7940, N7939, N7938, N7937, N7936, N7935, N7934, N7933, N7932, N7931, N7930, N7929, N7928, N7927, N7926, N7925, N7924, N7923, N7922, N7921, N7920, N7919, N7918, N7917, N7916, N7915, N7914, N7913, N7912, N7911, N7910, N7909, N7908, N7907, N7906, N7905, N7904, N7903, N7902, N7901, N7900, N7899, N7898, N7897, N7896, N7895, N7894, N7893, N7892, N7891, N7890, N7889, N7888, N7887, N7886, N7885, N7884, N7883, N7882, N7881, N7880, N7879, N7878, N7877, N7876, N7875, N7874, N7873, N7872, N7871, N7870, N7869, N7868, N7867, N7866, N7865, N7864, N7863, N7862, N7861, N7860, N7859, N7858, N7857, N7856, N7855, N7854, N7853, N7852, N7851, N7850, N7849, N7848, N7847, N7846, N7845, N7844, N7843, N7842, N7841, N7840, N7839, N7838, N7837, N7836, N7835, N7834, N7833, N7832, N7831, N7830, N7829, N7828, N7827, N7826, N7825, N7824, N7823, N7822, N7821, N7820, N7819, N7818, N7817, N7816, N7815, N7814, N7813, N7812, N7811, N7810, N7809, N7808, N7807, N7806, N7805, N7804, N7803, N7802, N7801, N7800, N7799, N7798, N7797, N7796, N7795, N7794, N7793, N7792, N7791, N7790, N7789, N7788, N7787, N7786, N7785, N7784, N7783, N7782, N7781, N7780, N7779, N7778, N7777, N7776, N7775, N7774, N7773, N7772, N7771, N7770, N7769, N7768, N7767, N7766, N7765, N7764, N7763, N7762, N7761, N7760, N7759, N7758, N7757, N7756, N7755, N7754, N7753, N7752, N7751, N7750, N7749, N7748, N7747, N7746, N7745, N7744, N7743, N7742, N7741, N7740, N7739, N7738, N7737, N7736, N7735, N7734, N7733, N7732, N7731, N7730, N7729, N7728, N7727, N7726, N7725, N7724, N7723, N7722, N7721, N7720, N7719, N7718, N7717, N7716, N7715, N7714, N7713, N7712, N7711, N7710, N7709, N7708, N7707, N7706, N7705, N7704, N7703, N7702, N7701, N7700, N7699, N7698, N7697, N7696, N7695, N7694, N7693, N7692, N7691, N7690, N7689, N7688, N7687, N7686, N7685, N7684, N7683, N7682, N7681, N7680, N7679, N7678, N7677, N7676, N7675, N7674, N7673, N7672, N7671, N7670, N7669, N7668, N7667, N7666, N7665, N7664, N7663, N7662, N7661, N7660, N7659, N7658, N7657, N7656, N7655, N7654, N7653, N7652, N7651, N7650, N7649, N7648, N7647, N7646, N7645, N7644, N7643, N7642, N7641, N7640, N7639, N7638, N7637, N7636, N7635, N7634, N7633, N7632, N7631, N7630, N7629, N7628, N7627, N7626, N7625, N7624, N7623, N7622, N7621, N7620, N7619, N7618, N7617, N7616, N7615, N7614, N7613, N7612, N7611, N7610, N7609, N7608, N7607, N7606, N7605, N7604, N7603, N7602, N7601, N7600, N7599, N7598, N7597, N7596, N7595, N7594, N7593, N7592, N7591, N7590, N7589, N7588, N7587, N7586, N7585, N7584, N7583, N7582, N7581, N7580, N7579, N7578, N7577, N7576, N7575, N7574, N7573, N7572, N7571, N7570, N7569, N7568, N7567, N7566, N7565, N7564, N7563, N7562, N7561, N7560, N7559, N7558, N7557, N7556, N7555, N7554, N7553, N7552, N7551, N7550, N7549, N7548, N7547, N7546, N7545, N7544, N7543, N7542, N7541, N7540, N7539, N7538, N7537, N7536, N7535, N7534, N7533, N7532, N7531, N7530, N7529, N7528, N7527, N7526, N7525, N7524, N7523, N7522, N7521, N7520, N7519, N7518, N7517, N7516, N7515, N7514, N7513, N7512, N7511, N7510, N7509, N7508, N7507, N7506, N7505, N7504, N7503, N7502, N7501, N7500, N7499, N7498, N7497, N7496, N7495, N7494, N7493, N7492, N7491, N7490, N7489, N7488, N7487, N7486, N7485, N7484, N7483, N7482, N7481, N7480, N7479, N7478, N7477, N7476, N7475, N7474, N7473, N7472, N7471, N7470, N7469, N7468, N7467, N7466, N7465, N7464, N7463, N7462, N7461, N7460, N7459, N7458, N7457, N7456, N7455, N7454, N7453, N7452, N7451, N7450, N7449, N7448, N7447, N7446, N7445, N7444, N7443, N7442, N7441, N7440, N7439, N7438, N7437, N7436, N7435, N7434, N7433, N7432, N7431, N7430, N7429, N7428, N7427, N7426, N7425, N7424, N7423, N7422, N7421, N7420, N7419, N7418, N7417, N7416, N7415, N7414, N7413, N7412, N7411, N7410, N7409, N7408, N7407, N7406, N7405, N7404, N7403, N7402, N7401, N7400, N7399, N7398, N7397, N7396, N7395, N7394, N7393, N7392, N7391, N7390, N7389, N7388, N7387, N7386, N7385, N7384, N7383, N7382, N7381, N7380, N7379, N7378, N7377, N7376, N7375, N7374, N7373, N7372, N7371, N7370, N7369, N7368, N7367, N7366, N7365, N7364, N7363, N7362, N7361, N7360, N7359, N7358, N7357, N7356, N7355, N7354, N7353, N7352, N7351, N7350, N7349, N7348, N7347, N7346, N7345, N7344, N7343, N7342, N7341, N7340, N7339, N7338, N7337, N7336, N7335, N7334, N7333, N7332, N7331, N7330, N7329, N7328, N7327, N7326, N7325, N7324, N7323, N7322, N7321, N7320, N7319, N7318, N7317, N7316, N7315, N7314, N7313, N7312, N7311, N7310, N7309, N7308, N7307, N7306, N7305, N7304, N7303, N7302, N7301, N7300, N7299, N7298, N7297, N7296, N7295, N7294, N7293, N7292, N7291, N7290, N7289, N7288, N7287, N7286, N7285, N7284, N7283, N7282, N7281, N7280, N7279, N7278, N7277, N7276, N7275, N7274, N7273, N7272, N7271, N7270, N7269, N7268, N7267, N7266, N7265, N7264, N7263, N7262, N7261, N7260, N7259, N7258, N7257, N7256, N7255, N7254, N7253, N7252, N7251, N7250, N7249, N7248, N7247, N7246, N7245, N7244, N7243, N7242, N7241, N7240, N7239, N7238, N7237, N7236, N7235, N7234, N7233, N7232, N7231, N7230, N7229, N7228, N7227, N7226, N7225, N7224, N7223, N7222, N7221, N7220, N7219, N7218, N7217, N7216, N7215, N7214, N7213, N7212, N7211, N7210, N7209, N7208, N7207, N7206, N7205, N7204, N7203, N7202, N7201, N7200, N7199, N7198, N7197, N7196, N7195, N7194, N7193, N7192, N7191, N7190, N7189, N7188, N7187, N7186, N7185, N7184, N7183, N7182, N7181, N7180, N7179, N7178, N7177, N7176, N7175, N7174, N7173, N7172, N7171, N7170, N7169, N7168, N7167, N7166, N7165, N7164, N7163, N7162, N7161, N7160, N7159, N7158, N7157, N7156, N7155, N7154, N7153, N7152, N7151, N7150, N7149, N7148, N7147, N7146, N7145, N7144, N7143, N7142, N7141, N7140, N7139, N7138, N7137, N7136, N7135, N7134, N7133, N7132, N7131, N7130, N7129, N7128, N7127, N7126, N7125, N7124, N7123, N7122, N7121, N7120, N7119, N7118, N7117, N7116, N7115, N7114, N7113, N7112, N7111, N7110, N7109, N7108, N7107, N7106, N7105, N7104, N7103, N7102, N7101, N7100, N7099, N7098, N7097, N7096, N7095, N7094, N7093, N7092, N7091, N7090, N7089, N7088, N7087, N7086, N7085, N7084, N7083, N7082, N7081, N7080, N7079, N7078, N7077, N7076, N7075, N7074, N7073, N7072, N7071, N7070, N7069, N7068, N7067, N7066, N7065, N7064, N7063, N7062, N7061, N7060, N7059, N7058, N7057, N7056, N7055, N7054, N7053, N7052, N7051, N7050, N7049, N7048, N7047, N7046, N7045, N7044, N7043, N7042, N7041, N7040, N7039, N7038, N7037, N7036, N7035, N7034, N7033, N7032, N7031, N7030, N7029, N7028, N7027, N7026, N7025, N7024, N7023, N7022, N7021, N7020, N7019, N7018, N7017, N7016, N7015, N7014, N7013, N7012, N7011, N7010, N7009, N7008, N7007, N7006, N7005, N7004, N7003, N7002, N7001, N7000, N6999, N6998, N6997, N6996, N6995, N6994, N6993, N6992, N6991, N6990, N6989, N6988, N6987, N6986, N6985, N6984, N6983, N6982, N6981, N6980, N6979, N6978, N6977, N6976, N6975, N6974, N6973, N6972, N6971, N6970, N6969, N6968, N6967, N6966, N6965, N6964, N6963, N6962, N6961, N6960, N6959, N6958, N6957, N6956, N6955, N6954, N6953, N6952, N6951, N6950, N6949, N6948, N6947, N6946, N6945, N6944, N6943, N6942, N6941, N6940, N6939, N6938, N6937, N6936, N6935, N6934, N6933, N6932, N6931, N6930, N6929, N6928, N6927, N6926, N6925, N6924, N6923, N6922, N6921, N6920, N6919, N6918, N6917, N6916, N6915, N6914, N6913, N6912, N6911, N6910, N6909, N6908, N6907, N6906, N6905, N6904, N6903, N6902, N6901, N6900, N6899, N6898, N6897, N6896, N6895, N6894, N6893, N6892, N6891, N6890, N6889, N6888, N6887, N6886, N6885, N6884, N6883, N6882, N6881, N6880, N6879, N6878, N6877, N6876, N6875, N6874, N6873, N6872, N6871, N6870, N6869, N6868, N6867, N6866, N6865, N6864, N6863, N6862, N6861, N6860, N6859, N6858, N6857, N6856, N6855, N6854, N6853, N6852, N6851, N6850, N6849, N6848, N6847, N6846, N6845, N6844, N6843, N6842, N6841, N6840, N6839, N6838, N6837, N6836, N6835, N6834, N6833, N6832, N6831, N6830, N6829, N6828, N6827, N6826, N6825, N6824, N6823, N6822, N6821, N6820, N6819, N6818, N6817, N6816, N6815, N6814, N6813, N6812, N6811, N6810, N6809, N6808, N6807, N6806, N6805, N6804, N6803, N6802, N6801, N6800, N6799, N6798, N6797, N6796, N6795, N6794, N6793, N6792, N6791, N6790, N6789, N6788, N6787, N6786, N6785, N6784, N6783, N6782, N6781, N6780, N6779, N6778, N6777, N6776, N6775, N6774, N6773, N6772, N6771, N6770, N6769, N6768, N6767, N6766, N6765, N6764, N6763, N6762, N6761, N6760, N6759, N6758, N6757, N6756, N6755, N6754, N6753, N6752, N6751, N6750, N6749, N6748, N6747, N6746, N6745, N6744, N6743, N6742, N6741, N6740, N6739, N6738, N6737, N6736, N6735, N6734, N6733, N6732, N6731, N6730, N6729, N6728, N6727, N6726, N6725, N6724, N6723, N6722, N6721, N6720, N6719, N6718, N6717, N6716, N6715, N6714, N6713, N6712, N6711, N6710, N6709, N6708, N6707, N6706, N6705, N6704, N6703, N6702, N6701, N6700, N6699, N6698, N6697, N6696, N6695, N6694, N6693, N6692, N6691, N6690, N6689, N6688, N6687, N6686, N6685, N6684, N6683, N6682, N6681, N6680, N6679, N6678, N6677, N6676, N6675, N6674, N6673, N6672, N6671, N6670, N6669, N6668, N6667, N6666, N6665, N6664, N6663, N6662, N6661, N6660, N6659, N6658, N6657, N6656, N6655, N6654, N6653, N6652, N6651, N6650, N6649, N6648, N6647, N6646, N6645, N6644, N6643, N6642, N6641, N6640, N6639, N6638, N6637, N6636, N6635, N6634, N6633, N6632, N6631, N6630, N6629, N6628, N6627, N6626, N6625, N6624, N6623, N6622, N6621, N6620, N6619, N6618, N6617, N6616, N6615, N6614, N6613, N6612, N6611, N6610, N6609, N6608, N6607, N6606, N6605, N6604, N6603, N6602, N6601, N6600, N6599, N6598, N6597, N6596, N6595, N6594, N6593, N6592, N6591, N6590, N6589, N6588, N6587, N6586, N6585, N6584, N6583, N6582, N6581, N6580, N6579, N6578, N6577, N6576, N6575, N6574, N6573, N6572, N6571, N6570, N6569, N6568, N6567, N6566, N6565, N6564, N6563, N6562, N6561, N6560, N6559, N6558, N6557, N6556, N6555, N6554, N6553, N6552, N6551, N6550, N6549, N6548, N6547, N6546, N6545, N6544, N6543, N6542, N6541, N6540, N6539, N6538, N6537, N6536, N6535, N6534, N6533, N6532, N6531, N6530, N6529, N6528, N6527, N6526, N6525, N6524, N6523, N6522, N6521, N6520, N6519, N6518, N6517, N6516, N6515, N6514, N6513, N6512, N6511, N6510, N6509, N6508, N6507, N6506, N6505, N6504, N6503, N6502, N6501, N6500, N6499, N6498, N6497, N6496, N6495, N6494, N6493, N6492, N6491, N6490, N6489, N6488, N6487, N6486, N6485, N6484, N6483, N6482, N6481, N6480, N6479, N6478, N6477, N6476, N6475, N6474, N6473, N6472, N6471, N6470, N6469, N6468, N6467, N6466, N6465, N6464, N6463, N6462, N6461, N6460, N6459, N6458, N6457, N6456, N6455, N6454, N6453, N6452, N6451, N6450, N6449, N6448, N6447, N6446, N6445, N6444, N6443, N6442, N6441, N6440, N6439, N6438, N6437, N6436, N6435, N6434, N6433, N6432, N6431, N6430, N6429, N6428, N6427, N6426, N6425, N6424, N6423, N6422, N6421, N6420, N6419, N6418, N6417, N6416, N6415, N6414, N6413, N6412, N6411, N6410, N6409, N6408, N6407, N6406, N6405, N6404, N6403, N6402, N6401, N6400, N6399, N6398, N6397, N6396, N6395, N6394, N6393, N6392, N6391, N6390, N6389, N6388, N6387, N6386, N6385, N6384, N6383, N6382, N6381, N6380, N6379, N6378, N6377 } = (N96)? { N6376, N6247, N6127, N6007, N5927, N5847, N5782, N5717, N5652, N5587, N5522, N5457, N5392, N5288, N5223, N5126, N5061, N4996, N4917, N4852, N4787, N4722, N4657, N4592, N4527, N4423, N4310, N4197, N4084, N4005, N3940, N3875, N3810, N3745, N3680, N3615, N3550, N3446, N3381, N3316, N3213, N3148, N3083, N3018, N2953, N2888, N2823, N2758, N2693, N2589, N2524, N2395, N2275, N2155, N2082, N2017, N1952, N1887, N1822, N1757, N1692, N1627, N1562, N1458, N1393, N1296, N1231, N1166, N1101, N1036, N965, N900, N835, N770, N705, N601, N488, N423, N358, N293, N6375, N6246, N6126, N6006, N5926, N5846, N5781, N5716, N5651, N5586, N5521, N5456, N5391, N5287, N5222, N5125, N5060, N4995, N4916, N4851, N4786, N4721, N4656, N4591, N4526, N4422, N4309, N4196, N4083, N4004, N3939, N3874, N3809, N3744, N3679, N3614, N3549, N3445, N3380, N3315, N3212, N3147, N3082, N3017, N2952, N2887, N2822, N2757, N2692, N2588, N2523, N2394, N2274, N2154, N2081, N2016, N1951, N1886, N1821, N1756, N1691, N1626, N1561, N1457, N1392, N1295, N1230, N1165, N1100, N1035, N964, N899, N834, N769, N704, N600, N487, N422, N357, N292, N6374, N6245, N6125, N6005, N5925, N5845, N5780, N5715, N5650, N5585, N5520, N5455, N5390, N5286, N5221, N5124, N5059, N4994, N4915, N4850, N4785, N4720, N4655, N4590, N4525, N4421, N4308, N4195, N4082, N4003, N3938, N3873, N3808, N3743, N3678, N3613, N3548, N3444, N3379, N3314, N3211, N3146, N3081, N3016, N2951, N2886, N2821, N2756, N2691, N2587, N2522, N2393, N2273, N2153, N2080, N2015, N1950, N1885, N1820, N1755, N1690, N1625, N1560, N1456, N1391, N1294, N1229, N1164, N1099, N1034, N963, N898, N833, N768, N703, N599, N486, N421, N356, N291, N6373, N6244, N6124, N6004, N5924, N5844, N5779, N5714, N5649, N5584, N5519, N5454, N5389, N5285, N5220, N5123, N5058, N4993, N4914, N4849, N4784, N4719, N4654, N4589, N4524, N4420, N4307, N4194, N4081, N4002, N3937, N3872, N3807, N3742, N3677, N3612, N3547, N3443, N3378, N3313, N3210, N3145, N3080, N3015, N2950, N2885, N2820, N2755, N2690, N2586, N2521, N2392, N2272, N2152, N2079, N2014, N1949, N1884, N1819, N1754, N1689, N1624, N1559, N1455, N1390, N1293, N1228, N1163, N1098, N1033, N962, N897, N832, N767, N702, N598, N485, N420, N355, N290, N6372, N6243, N6123, N6003, N5923, N5843, N5778, N5713, N5648, N5583, N5518, N5453, N5388, N5284, N5219, N5122, N5057, N4992, N4913, N4848, N4783, N4718, N4653, N4588, N4523, N4419, N4306, N4193, N4080, N4001, N3936, N3871, N3806, N3741, N3676, N3611, N3546, N3442, N3377, N3312, N3209, N3144, N3079, N3014, N2949, N2884, N2819, N2754, N2689, N2585, N2520, N2391, N2271, N2151, N2078, N2013, N1948, N1883, N1818, N1753, N1688, N1623, N1558, N1454, N1389, N1292, N1227, N1162, N1097, N1032, N961, N896, N831, N766, N701, N597, N484, N419, N354, N289, N6371, N6242, N6122, N6002, N5922, N5842, N5777, N5712, N5647, N5582, N5517, N5452, N5387, N5283, N5218, N5121, N5056, N4991, N4912, N4847, N4782, N4717, N4652, N4587, N4522, N4418, N4305, N4192, N4079, N4000, N3935, N3870, N3805, N3740, N3675, N3610, N3545, N3441, N3376, N3311, N3208, N3143, N3078, N3013, N2948, N2883, N2818, N2753, N2688, N2584, N2519, N2390, N2270, N2150, N2077, N2012, N1947, N1882, N1817, N1752, N1687, N1622, N1557, N1453, N1388, N1291, N1226, N1161, N1096, N1031, N960, N895, N830, N765, N700, N596, N483, N418, N353, N288, N6370, N6241, N6121, N6001, N5921, N5841, N5776, N5711, N5646, N5581, N5516, N5451, N5386, N5282, N5217, N5120, N5055, N4990, N4911, N4846, N4781, N4716, N4651, N4586, N4521, N4417, N4304, N4191, N4078, N3999, N3934, N3869, N3804, N3739, N3674, N3609, N3544, N3440, N3375, N3310, N3207, N3142, N3077, N3012, N2947, N2882, N2817, N2752, N2687, N2583, N2518, N2389, N2269, N2149, N2076, N2011, N1946, N1881, N1816, N1751, N1686, N1621, N1556, N1452, N1387, N1290, N1225, N1160, N1095, N1030, N959, N894, N829, N764, N699, N595, N482, N417, N352, N287, N6369, N6240, N6120, N6000, N5920, N5840, N5775, N5710, N5645, N5580, N5515, N5450, N5385, N5281, N5216, N5119, N5054, N4989, N4910, N4845, N4780, N4715, N4650, N4585, N4520, N4416, N4303, N4190, N4077, N3998, N3933, N3868, N3803, N3738, N3673, N3608, N3543, N3439, N3374, N3309, N3206, N3141, N3076, N3011, N2946, N2881, N2816, N2751, N2686, N2582, N2517, N2388, N2268, N2148, N2075, N2010, N1945, N1880, N1815, N1750, N1685, N1620, N1555, N1451, N1386, N1289, N1224, N1159, N1094, N1029, N958, N893, N828, N763, N698, N594, N481, N416, N351, N286, N6368, N6239, N6119, N5999, N5919, N5839, N5774, N5709, N5644, N5579, N5514, N5449, N5384, N5280, N5215, N5118, N5053, N4988, N4909, N4844, N4779, N4714, N4649, N4584, N4519, N4415, N4302, N4189, N4076, N3997, N3932, N3867, N3802, N3737, N3672, N3607, N3542, N3438, N3373, N3308, N3205, N3140, N3075, N3010, N2945, N2880, N2815, N2750, N2685, N2581, N2516, N2387, N2267, N2147, N2074, N2009, N1944, N1879, N1814, N1749, N1684, N1619, N1554, N1450, N1385, N1288, N1223, N1158, N1093, N1028, N957, N892, N827, N762, N697, N593, N480, N415, N350, N285, N6367, N6238, N6118, N5998, N5918, N5838, N5773, N5708, N5643, N5578, N5513, N5448, N5383, N5279, N5214, N5117, N5052, N4987, N4908, N4843, N4778, N4713, N4648, N4583, N4518, N4414, N4301, N4188, N4075, N3996, N3931, N3866, N3801, N3736, N3671, N3606, N3541, N3437, N3372, N3307, N3204, N3139, N3074, N3009, N2944, N2879, N2814, N2749, N2684, N2580, N2515, N2386, N2266, N2146, N2073, N2008, N1943, N1878, N1813, N1748, N1683, N1618, N1553, N1449, N1384, N1287, N1222, N1157, N1092, N1027, N956, N891, N826, N761, N696, N592, N479, N414, N349, N284, N6366, N6237, N6117, N5997, N5917, N5837, N5772, N5707, N5642, N5577, N5512, N5447, N5382, N5278, N5213, N5116, N5051, N4986, N4907, N4842, N4777, N4712, N4647, N4582, N4517, N4413, N4300, N4187, N4074, N3995, N3930, N3865, N3800, N3735, N3670, N3605, N3540, N3436, N3371, N3306, N3203, N3138, N3073, N3008, N2943, N2878, N2813, N2748, N2683, N2579, N2514, N2385, N2265, N2145, N2072, N2007, N1942, N1877, N1812, N1747, N1682, N1617, N1552, N1448, N1383, N1286, N1221, N1156, N1091, N1026, N955, N890, N825, N760, N695, N591, N478, N413, N348, N283, N6365, N6236, N6116, N5996, N5916, N5836, N5771, N5706, N5641, N5576, N5511, N5446, N5381, N5277, N5212, N5115, N5050, N4985, N4906, N4841, N4776, N4711, N4646, N4581, N4516, N4412, N4299, N4186, N4073, N3994, N3929, N3864, N3799, N3734, N3669, N3604, N3539, N3435, N3370, N3305, N3202, N3137, N3072, N3007, N2942, N2877, N2812, N2747, N2682, N2578, N2513, N2384, N2264, N2144, N2071, N2006, N1941, N1876, N1811, N1746, N1681, N1616, N1551, N1447, N1382, N1285, N1220, N1155, N1090, N1025, N954, N889, N824, N759, N694, N590, N477, N412, N347, N282, N6364, N6235, N6115, N5995, N5915, N5835, N5770, N5705, N5640, N5575, N5510, N5445, N5380, N5276, N5211, N5114, N5049, N4984, N4905, N4840, N4775, N4710, N4645, N4580, N4515, N4411, N4298, N4185, N4072, N3993, N3928, N3863, N3798, N3733, N3668, N3603, N3538, N3434, N3369, N3304, N3201, N3136, N3071, N3006, N2941, N2876, N2811, N2746, N2681, N2577, N2512, N2383, N2263, N2143, N2070, N2005, N1940, N1875, N1810, N1745, N1680, N1615, N1550, N1446, N1381, N1284, N1219, N1154, N1089, N1024, N953, N888, N823, N758, N693, N589, N476, N411, N346, N281, N6363, N6234, N6114, N5994, N5914, N5834, N5769, N5704, N5639, N5574, N5509, N5444, N5379, N5275, N5210, N5113, N5048, N4983, N4904, N4839, N4774, N4709, N4644, N4579, N4514, N4410, N4297, N4184, N4071, N3992, N3927, N3862, N3797, N3732, N3667, N3602, N3537, N3433, N3368, N3303, N3200, N3135, N3070, N3005, N2940, N2875, N2810, N2745, N2680, N2576, N2511, N2382, N2262, N2142, N2069, N2004, N1939, N1874, N1809, N1744, N1679, N1614, N1549, N1445, N1380, N1283, N1218, N1153, N1088, N1023, N952, N887, N822, N757, N692, N588, N475, N410, N345, N280, N6362, N6233, N6113, N5993, N5913, N5833, N5768, N5703, N5638, N5573, N5508, N5443, N5378, N5274, N5209, N5112, N5047, N4982, N4903, N4838, N4773, N4708, N4643, N4578, N4513, N4409, N4296, N4183, N4070, N3991, N3926, N3861, N3796, N3731, N3666, N3601, N3536, N3432, N3367, N3302, N3199, N3134, N3069, N3004, N2939, N2874, N2809, N2744, N2679, N2575, N2510, N2381, N2261, N2141, N2068, N2003, N1938, N1873, N1808, N1743, N1678, N1613, N1548, N1444, N1379, N1282, N1217, N1152, N1087, N1022, N951, N886, N821, N756, N691, N587, N474, N409, N344, N279, N6361, N6232, N6112, N5992, N5912, N5832, N5767, N5702, N5637, N5572, N5507, N5442, N5377, N5273, N5208, N5111, N5046, N4981, N4902, N4837, N4772, N4707, N4642, N4577, N4512, N4408, N4295, N4182, N4069, N3990, N3925, N3860, N3795, N3730, N3665, N3600, N3535, N3431, N3366, N3301, N3198, N3133, N3068, N3003, N2938, N2873, N2808, N2743, N2678, N2574, N2509, N2380, N2260, N2140, N2067, N2002, N1937, N1872, N1807, N1742, N1677, N1612, N1547, N1443, N1378, N1281, N1216, N1151, N1086, N1021, N950, N885, N820, N755, N690, N586, N473, N408, N343, N278, N6360, N6231, N6111, N5991, N5911, N5831, N5766, N5701, N5636, N5571, N5506, N5441, N5376, N5272, N5207, N5110, N5045, N4980, N4901, N4836, N4771, N4706, N4641, N4576, N4511, N4407, N4294, N4181, N4068, N3989, N3924, N3859, N3794, N3729, N3664, N3599, N3534, N3430, N3365, N3300, N3197, N3132, N3067, N3002, N2937, N2872, N2807, N2742, N2677, N2573, N2508, N2379, N2259, N2139, N2066, N2001, N1936, N1871, N1806, N1741, N1676, N1611, N1546, N1442, N1377, N1280, N1215, N1150, N1085, N1020, N949, N884, N819, N754, N689, N585, N472, N407, N342, N277, N6359, N6230, N6110, N5990, N5910, N5830, N5765, N5700, N5635, N5570, N5505, N5440, N5375, N5271, N5206, N5109, N5044, N4979, N4900, N4835, N4770, N4705, N4640, N4575, N4510, N4406, N4293, N4180, N4067, N3988, N3923, N3858, N3793, N3728, N3663, N3598, N3533, N3429, N3364, N3299, N3196, N3131, N3066, N3001, N2936, N2871, N2806, N2741, N2676, N2572, N2507, N2378, N2258, N2138, N2065, N2000, N1935, N1870, N1805, N1740, N1675, N1610, N1545, N1441, N1376, N1279, N1214, N1149, N1084, N1019, N948, N883, N818, N753, N688, N584, N471, N406, N341, N276, N6358, N6229, N6109, N5989, N5909, N5829, N5764, N5699, N5634, N5569, N5504, N5439, N5374, N5270, N5205, N5108, N5043, N4978, N4899, N4834, N4769, N4704, N4639, N4574, N4509, N4405, N4292, N4179, N4066, N3987, N3922, N3857, N3792, N3727, N3662, N3597, N3532, N3428, N3363, N3298, N3195, N3130, N3065, N3000, N2935, N2870, N2805, N2740, N2675, N2571, N2506, N2377, N2257, N2137, N2064, N1999, N1934, N1869, N1804, N1739, N1674, N1609, N1544, N1440, N1375, N1278, N1213, N1148, N1083, N1018, N947, N882, N817, N752, N687, N583, N470, N405, N340, N275, N6357, N6228, N6108, N5988, N5908, N5828, N5763, N5698, N5633, N5568, N5503, N5438, N5373, N5269, N5204, N5107, N5042, N4977, N4898, N4833, N4768, N4703, N4638, N4573, N4508, N4404, N4291, N4178, N4065, N3986, N3921, N3856, N3791, N3726, N3661, N3596, N3531, N3427, N3362, N3297, N3194, N3129, N3064, N2999, N2934, N2869, N2804, N2739, N2674, N2570, N2505, N2376, N2256, N2136, N2063, N1998, N1933, N1868, N1803, N1738, N1673, N1608, N1543, N1439, N1374, N1277, N1212, N1147, N1082, N1017, N946, N881, N816, N751, N686, N582, N469, N404, N339, N274, N6356, N6227, N6107, N5987, N5907, N5827, N5762, N5697, N5632, N5567, N5502, N5437, N5372, N5268, N5203, N5106, N5041, N4976, N4897, N4832, N4767, N4702, N4637, N4572, N4507, N4403, N4290, N4177, N4064, N3985, N3920, N3855, N3790, N3725, N3660, N3595, N3530, N3426, N3361, N3296, N3193, N3128, N3063, N2998, N2933, N2868, N2803, N2738, N2673, N2569, N2504, N2375, N2255, N2135, N2062, N1997, N1932, N1867, N1802, N1737, N1672, N1607, N1542, N1438, N1373, N1276, N1211, N1146, N1081, N1016, N945, N880, N815, N750, N685, N581, N468, N403, N338, N273, N6355, N6226, N6106, N5986, N5906, N5826, N5761, N5696, N5631, N5566, N5501, N5436, N5371, N5267, N5202, N5105, N5040, N4975, N4896, N4831, N4766, N4701, N4636, N4571, N4506, N4402, N4289, N4176, N4063, N3984, N3919, N3854, N3789, N3724, N3659, N3594, N3529, N3425, N3360, N3295, N3192, N3127, N3062, N2997, N2932, N2867, N2802, N2737, N2672, N2568, N2503, N2374, N2254, N2134, N2061, N1996, N1931, N1866, N1801, N1736, N1671, N1606, N1541, N1437, N1372, N1275, N1210, N1145, N1080, N1015, N944, N879, N814, N749, N684, N580, N467, N402, N337, N272, N6354, N6225, N6105, N5985, N5905, N5825, N5760, N5695, N5630, N5565, N5500, N5435, N5370, N5266, N5201, N5104, N5039, N4974, N4895, N4830, N4765, N4700, N4635, N4570, N4505, N4401, N4288, N4175, N4062, N3983, N3918, N3853, N3788, N3723, N3658, N3593, N3528, N3424, N3359, N3294, N3191, N3126, N3061, N2996, N2931, N2866, N2801, N2736, N2671, N2567, N2502, N2373, N2253, N2133, N2060, N1995, N1930, N1865, N1800, N1735, N1670, N1605, N1540, N1436, N1371, N1274, N1209, N1144, N1079, N1014, N943, N878, N813, N748, N683, N579, N466, N401, N336, N271, N6353, N6224, N6104, N5984, N5904, N5824, N5759, N5694, N5629, N5564, N5499, N5434, N5369, N5265, N5200, N5103, N5038, N4973, N4894, N4829, N4764, N4699, N4634, N4569, N4504, N4400, N4287, N4174, N4061, N3982, N3917, N3852, N3787, N3722, N3657, N3592, N3527, N3423, N3358, N3293, N3190, N3125, N3060, N2995, N2930, N2865, N2800, N2735, N2670, N2566, N2501, N2372, N2252, N2132, N2059, N1994, N1929, N1864, N1799, N1734, N1669, N1604, N1539, N1435, N1370, N1273, N1208, N1143, N1078, N1013, N942, N877, N812, N747, N682, N578, N465, N400, N335, N270, N6352, N6223, N6103, N5983, N5903, N5823, N5758, N5693, N5628, N5563, N5498, N5433, N5368, N5264, N5199, N5102, N5037, N4972, N4893, N4828, N4763, N4698, N4633, N4568, N4503, N4399, N4286, N4173, N4060, N3981, N3916, N3851, N3786, N3721, N3656, N3591, N3526, N3422, N3357, N3292, N3189, N3124, N3059, N2994, N2929, N2864, N2799, N2734, N2669, N2565, N2500, N2371, N2251, N2131, N2058, N1993, N1928, N1863, N1798, N1733, N1668, N1603, N1538, N1434, N1369, N1272, N1207, N1142, N1077, N1012, N941, N876, N811, N746, N681, N577, N464, N399, N334, N269, N6351, N6222, N6102, N5982, N5902, N5822, N5757, N5692, N5627, N5562, N5497, N5432, N5367, N5263, N5198, N5101, N5036, N4971, N4892, N4827, N4762, N4697, N4632, N4567, N4502, N4398, N4285, N4172, N4059, N3980, N3915, N3850, N3785, N3720, N3655, N3590, N3525, N3421, N3356, N3291, N3188, N3123, N3058, N2993, N2928, N2863, N2798, N2733, N2668, N2564, N2499, N2370, N2250, N2130, N2057, N1992, N1927, N1862, N1797, N1732, N1667, N1602, N1537, N1433, N1368, N1271, N1206, N1141, N1076, N1011, N940, N875, N810, N745, N680, N576, N463, N398, N333, N268, N6350, N6221, N6101, N5981, N5901, N5821, N5756, N5691, N5626, N5561, N5496, N5431, N5366, N5262, N5197, N5100, N5035, N4970, N4891, N4826, N4761, N4696, N4631, N4566, N4501, N4397, N4284, N4171, N4058, N3979, N3914, N3849, N3784, N3719, N3654, N3589, N3524, N3420, N3355, N3290, N3187, N3122, N3057, N2992, N2927, N2862, N2797, N2732, N2667, N2563, N2498, N2369, N2249, N2129, N2056, N1991, N1926, N1861, N1796, N1731, N1666, N1601, N1536, N1432, N1367, N1270, N1205, N1140, N1075, N1010, N939, N874, N809, N744, N679, N575, N462, N397, N332, N267, N6349, N6220, N6100, N5980, N5900, N5820, N5755, N5690, N5625, N5560, N5495, N5430, N5365, N5261, N5196, N5099, N5034, N4969, N4890, N4825, N4760, N4695, N4630, N4565, N4500, N4396, N4283, N4170, N4057, N3978, N3913, N3848, N3783, N3718, N3653, N3588, N3523, N3419, N3354, N3289, N3186, N3121, N3056, N2991, N2926, N2861, N2796, N2731, N2666, N2562, N2497, N2368, N2248, N2128, N2055, N1990, N1925, N1860, N1795, N1730, N1665, N1600, N1535, N1431, N1366, N1269, N1204, N1139, N1074, N1009, N938, N873, N808, N743, N678, N574, N461, N396, N331, N266, N6348, N6219, N6099, N5979, N5899, N5819, N5754, N5689, N5624, N5559, N5494, N5429, N5364, N5260, N5195, N5098, N5033, N4968, N4889, N4824, N4759, N4694, N4629, N4564, N4499, N4395, N4282, N4169, N4056, N3977, N3912, N3847, N3782, N3717, N3652, N3587, N3522, N3418, N3353, N3288, N3185, N3120, N3055, N2990, N2925, N2860, N2795, N2730, N2665, N2561, N2496, N2367, N2247, N2127, N2054, N1989, N1924, N1859, N1794, N1729, N1664, N1599, N1534, N1430, N1365, N1268, N1203, N1138, N1073, N1008, N937, N872, N807, N742, N677, N573, N460, N395, N330, N265, N6347, N6218, N6098, N5978, N5898, N5818, N5753, N5688, N5623, N5558, N5493, N5428, N5363, N5259, N5194, N5097, N5032, N4967, N4888, N4823, N4758, N4693, N4628, N4563, N4498, N4394, N4281, N4168, N4055, N3976, N3911, N3846, N3781, N3716, N3651, N3586, N3521, N3417, N3352, N3287, N3184, N3119, N3054, N2989, N2924, N2859, N2794, N2729, N2664, N2560, N2495, N2366, N2246, N2126, N2053, N1988, N1923, N1858, N1793, N1728, N1663, N1598, N1533, N1429, N1364, N1267, N1202, N1137, N1072, N1007, N936, N871, N806, N741, N676, N572, N459, N394, N329, N264, N6346, N6217, N6097, N5977, N5897, N5817, N5752, N5687, N5622, N5557, N5492, N5427, N5362, N5258, N5193, N5096, N5031, N4966, N4887, N4822, N4757, N4692, N4627, N4562, N4497, N4393, N4280, N4167, N4054, N3975, N3910, N3845, N3780, N3715, N3650, N3585, N3520, N3416, N3351, N3286, N3183, N3118, N3053, N2988, N2923, N2858, N2793, N2728, N2663, N2559, N2494, N2365, N2245, N2125, N2052, N1987, N1922, N1857, N1792, N1727, N1662, N1597, N1532, N1428, N1363, N1266, N1201, N1136, N1071, N1006, N935, N870, N805, N740, N675, N571, N458, N393, N328, N263, N6345, N6216, N6096, N5976, N5896, N5816, N5751, N5686, N5621, N5556, N5491, N5426, N5361, N5257, N5192, N5095, N5030, N4965, N4886, N4821, N4756, N4691, N4626, N4561, N4496, N4392, N4279, N4166, N4053, N3974, N3909, N3844, N3779, N3714, N3649, N3584, N3519, N3415, N3350, N3285, N3182, N3117, N3052, N2987, N2922, N2857, N2792, N2727, N2662, N2558, N2493, N2364, N2244, N2124, N2051, N1986, N1921, N1856, N1791, N1726, N1661, N1596, N1531, N1427, N1362, N1265, N1200, N1135, N1070, N1005, N934, N869, N804, N739, N674, N570, N457, N392, N327, N262, N6344, N6215, N6095, N5975, N5895, N5815, N5750, N5685, N5620, N5555, N5490, N5425, N5360, N5256, N5191, N5094, N5029, N4964, N4885, N4820, N4755, N4690, N4625, N4560, N4495, N4391, N4278, N4165, N4052, N3973, N3908, N3843, N3778, N3713, N3648, N3583, N3518, N3414, N3349, N3284, N3181, N3116, N3051, N2986, N2921, N2856, N2791, N2726, N2661, N2557, N2492, N2363, N2243, N2123, N2050, N1985, N1920, N1855, N1790, N1725, N1660, N1595, N1530, N1426, N1361, N1264, N1199, N1134, N1069, N1004, N933, N868, N803, N738, N673, N569, N456, N391, N326, N261, N6343, N6214, N6094, N5974, N5894, N5814, N5749, N5684, N5619, N5554, N5489, N5424, N5359, N5255, N5190, N5093, N5028, N4963, N4884, N4819, N4754, N4689, N4624, N4559, N4494, N4390, N4277, N4164, N4051, N3972, N3907, N3842, N3777, N3712, N3647, N3582, N3517, N3413, N3348, N3283, N3180, N3115, N3050, N2985, N2920, N2855, N2790, N2725, N2660, N2556, N2491, N2362, N2242, N2122, N2049, N1984, N1919, N1854, N1789, N1724, N1659, N1594, N1529, N1425, N1360, N1263, N1198, N1133, N1068, N1003, N932, N867, N802, N737, N672, N568, N455, N390, N325, N260, N6342, N6213, N6093, N5973, N5893, N5813, N5748, N5683, N5618, N5553, N5488, N5423, N5358, N5254, N5189, N5092, N5027, N4962, N4883, N4818, N4753, N4688, N4623, N4558, N4493, N4389, N4276, N4163, N4050, N3971, N3906, N3841, N3776, N3711, N3646, N3581, N3516, N3412, N3347, N3282, N3179, N3114, N3049, N2984, N2919, N2854, N2789, N2724, N2659, N2555, N2490, N2361, N2241, N2121, N2048, N1983, N1918, N1853, N1788, N1723, N1658, N1593, N1528, N1424, N1359, N1262, N1197, N1132, N1067, N1002, N931, N866, N801, N736, N671, N567, N454, N389, N324, N259, N6341, N6212, N6092, N5972, N5892, N5812, N5747, N5682, N5617, N5552, N5487, N5422, N5357, N5253, N5188, N5091, N5026, N4961, N4882, N4817, N4752, N4687, N4622, N4557, N4492, N4388, N4275, N4162, N4049, N3970, N3905, N3840, N3775, N3710, N3645, N3580, N3515, N3411, N3346, N3281, N3178, N3113, N3048, N2983, N2918, N2853, N2788, N2723, N2658, N2554, N2489, N2360, N2240, N2120, N2047, N1982, N1917, N1852, N1787, N1722, N1657, N1592, N1527, N1423, N1358, N1261, N1196, N1131, N1066, N1001, N930, N865, N800, N735, N670, N566, N453, N388, N323, N258, N6340, N6211, N6091, N5971, N5891, N5811, N5746, N5681, N5616, N5551, N5486, N5421, N5356, N5252, N5187, N5090, N5025, N4960, N4881, N4816, N4751, N4686, N4621, N4556, N4491, N4387, N4274, N4161, N4048, N3969, N3904, N3839, N3774, N3709, N3644, N3579, N3514, N3410, N3345, N3280, N3177, N3112, N3047, N2982, N2917, N2852, N2787, N2722, N2657, N2553, N2488, N2359, N2239, N2119, N2046, N1981, N1916, N1851, N1786, N1721, N1656, N1591, N1526, N1422, N1357, N1260, N1195, N1130, N1065, N1000, N929, N864, N799, N734, N669, N565, N452, N387, N322, N257, N6339, N6210, N6090, N5970, N5890, N5810, N5745, N5680, N5615, N5550, N5485, N5420, N5355, N5251, N5186, N5089, N5024, N4959, N4880, N4815, N4750, N4685, N4620, N4555, N4490, N4386, N4273, N4160, N4047, N3968, N3903, N3838, N3773, N3708, N3643, N3578, N3513, N3409, N3344, N3279, N3176, N3111, N3046, N2981, N2916, N2851, N2786, N2721, N2656, N2552, N2487, N2358, N2238, N2118, N2045, N1980, N1915, N1850, N1785, N1720, N1655, N1590, N1525, N1421, N1356, N1259, N1194, N1129, N1064, N999, N928, N863, N798, N733, N668, N564, N451, N386, N321, N256, N6338, N6209, N6089, N5969, N5889, N5809, N5744, N5679, N5614, N5549, N5484, N5419, N5354, N5250, N5185, N5088, N5023, N4958, N4879, N4814, N4749, N4684, N4619, N4554, N4489, N4385, N4272, N4159, N4046, N3967, N3902, N3837, N3772, N3707, N3642, N3577, N3512, N3408, N3343, N3278, N3175, N3110, N3045, N2980, N2915, N2850, N2785, N2720, N2655, N2551, N2486, N2357, N2237, N2117, N2044, N1979, N1914, N1849, N1784, N1719, N1654, N1589, N1524, N1420, N1355, N1258, N1193, N1128, N1063, N998, N927, N862, N797, N732, N667, N563, N450, N385, N320, N255, N6337, N6208, N6088, N5968, N5888, N5808, N5743, N5678, N5613, N5548, N5483, N5418, N5353, N5249, N5184, N5087, N5022, N4957, N4878, N4813, N4748, N4683, N4618, N4553, N4488, N4384, N4271, N4158, N4045, N3966, N3901, N3836, N3771, N3706, N3641, N3576, N3511, N3407, N3342, N3277, N3174, N3109, N3044, N2979, N2914, N2849, N2784, N2719, N2654, N2550, N2485, N2356, N2236, N2116, N2043, N1978, N1913, N1848, N1783, N1718, N1653, N1588, N1523, N1419, N1354, N1257, N1192, N1127, N1062, N997, N926, N861, N796, N731, N666, N562, N449, N384, N319, N254, N6336, N6207, N6087, N5967, N5887, N5807, N5742, N5677, N5612, N5547, N5482, N5417, N5352, N5248, N5183, N5086, N5021, N4956, N4877, N4812, N4747, N4682, N4617, N4552, N4487, N4383, N4270, N4157, N4044, N3965, N3900, N3835, N3770, N3705, N3640, N3575, N3510, N3406, N3341, N3276, N3173, N3108, N3043, N2978, N2913, N2848, N2783, N2718, N2653, N2549, N2484, N2355, N2235, N2115, N2042, N1977, N1912, N1847, N1782, N1717, N1652, N1587, N1522, N1418, N1353, N1256, N1191, N1126, N1061, N996, N925, N860, N795, N730, N665, N561, N448, N383, N318, N253, N6335, N6206, N6086, N5966, N5886, N5806, N5741, N5676, N5611, N5546, N5481, N5416, N5351, N5247, N5182, N5085, N5020, N4955, N4876, N4811, N4746, N4681, N4616, N4551, N4486, N4382, N4269, N4156, N4043, N3964, N3899, N3834, N3769, N3704, N3639, N3574, N3509, N3405, N3340, N3275, N3172, N3107, N3042, N2977, N2912, N2847, N2782, N2717, N2652, N2548, N2483, N2354, N2234, N2114, N2041, N1976, N1911, N1846, N1781, N1716, N1651, N1586, N1521, N1417, N1352, N1255, N1190, N1125, N1060, N995, N924, N859, N794, N729, N664, N560, N447, N382, N317, N252, N6334, N6205, N6085, N5965, N5885, N5805, N5740, N5675, N5610, N5545, N5480, N5415, N5350, N5246, N5181, N5084, N5019, N4954, N4875, N4810, N4745, N4680, N4615, N4550, N4485, N4381, N4268, N4155, N4042, N3963, N3898, N3833, N3768, N3703, N3638, N3573, N3508, N3404, N3339, N3274, N3171, N3106, N3041, N2976, N2911, N2846, N2781, N2716, N2651, N2547, N2482, N2353, N2233, N2113, N2040, N1975, N1910, N1845, N1780, N1715, N1650, N1585, N1520, N1416, N1351, N1254, N1189, N1124, N1059, N994, N923, N858, N793, N728, N663, N559, N446, N381, N316, N251, N6333, N6204, N6084, N5964, N5884, N5804, N5739, N5674, N5609, N5544, N5479, N5414, N5349, N5245, N5180, N5083, N5018, N4953, N4874, N4809, N4744, N4679, N4614, N4549, N4484, N4380, N4267, N4154, N4041, N3962, N3897, N3832, N3767, N3702, N3637, N3572, N3507, N3403, N3338, N3273, N3170, N3105, N3040, N2975, N2910, N2845, N2780, N2715, N2650, N2546, N2481, N2352, N2232, N2112, N2039, N1974, N1909, N1844, N1779, N1714, N1649, N1584, N1519, N1415, N1350, N1253, N1188, N1123, N1058, N993, N922, N857, N792, N727, N662, N558, N445, N380, N315, N250, N6332, N6203, N6083, N5963, N5883, N5803, N5738, N5673, N5608, N5543, N5478, N5413, N5348, N5244, N5179, N5082, N5017, N4952, N4873, N4808, N4743, N4678, N4613, N4548, N4483, N4379, N4266, N4153, N4040, N3961, N3896, N3831, N3766, N3701, N3636, N3571, N3506, N3402, N3337, N3272, N3169, N3104, N3039, N2974, N2909, N2844, N2779, N2714, N2649, N2545, N2480, N2351, N2231, N2111, N2038, N1973, N1908, N1843, N1778, N1713, N1648, N1583, N1518, N1414, N1349, N1252, N1187, N1122, N1057, N992, N921, N856, N791, N726, N661, N557, N444, N379, N314, N249, N6331, N6202, N6082, N5962, N5882, N5802, N5737, N5672, N5607, N5542, N5477, N5412, N5347, N5243, N5178, N5081, N5016, N4951, N4872, N4807, N4742, N4677, N4612, N4547, N4482, N4378, N4265, N4152, N4039, N3960, N3895, N3830, N3765, N3700, N3635, N3570, N3505, N3401, N3336, N3271, N3168, N3103, N3038, N2973, N2908, N2843, N2778, N2713, N2648, N2544, N2479, N2350, N2230, N2110, N2037, N1972, N1907, N1842, N1777, N1712, N1647, N1582, N1517, N1413, N1348, N1251, N1186, N1121, N1056, N991, N920, N855, N790, N725, N660, N556, N443, N378, N313, N248, N6330, N6201, N6081, N5961, N5881, N5801, N5736, N5671, N5606, N5541, N5476, N5411, N5346, N5242, N5177, N5080, N5015, N4950, N4871, N4806, N4741, N4676, N4611, N4546, N4481, N4377, N4264, N4151, N4038, N3959, N3894, N3829, N3764, N3699, N3634, N3569, N3504, N3400, N3335, N3270, N3167, N3102, N3037, N2972, N2907, N2842, N2777, N2712, N2647, N2543, N2478, N2349, N2229, N2109, N2036, N1971, N1906, N1841, N1776, N1711, N1646, N1581, N1516, N1412, N1347, N1250, N1185, N1120, N1055, N990, N919, N854, N789, N724, N659, N555, N442, N377, N312, N247, N6329, N6200, N6080, N5960, N5880, N5800, N5735, N5670, N5605, N5540, N5475, N5410, N5345, N5241, N5176, N5079, N5014, N4949, N4870, N4805, N4740, N4675, N4610, N4545, N4480, N4376, N4263, N4150, N4037, N3958, N3893, N3828, N3763, N3698, N3633, N3568, N3503, N3399, N3334, N3269, N3166, N3101, N3036, N2971, N2906, N2841, N2776, N2711, N2646, N2542, N2477, N2348, N2228, N2108, N2035, N1970, N1905, N1840, N1775, N1710, N1645, N1580, N1515, N1411, N1346, N1249, N1184, N1119, N1054, N989, N918, N853, N788, N723, N658, N554, N441, N376, N311, N246, N6328, N6199, N6079, N5959, N5879, N5799, N5734, N5669, N5604, N5539, N5474, N5409, N5344, N5240, N5175, N5078, N5013, N4948, N4869, N4804, N4739, N4674, N4609, N4544, N4479, N4375, N4262, N4149, N4036, N3957, N3892, N3827, N3762, N3697, N3632, N3567, N3502, N3398, N3333, N3268, N3165, N3100, N3035, N2970, N2905, N2840, N2775, N2710, N2645, N2541, N2476, N2347, N2227, N2107, N2034, N1969, N1904, N1839, N1774, N1709, N1644, N1579, N1514, N1410, N1345, N1248, N1183, N1118, N1053, N988, N917, N852, N787, N722, N657, N553, N440, N375, N310, N245, N6327, N6198, N6078, N5958, N5878, N5798, N5733, N5668, N5603, N5538, N5473, N5408, N5343, N5239, N5174, N5077, N5012, N4947, N4868, N4803, N4738, N4673, N4608, N4543, N4478, N4374, N4261, N4148, N4035, N3956, N3891, N3826, N3761, N3696, N3631, N3566, N3501, N3397, N3332, N3267, N3164, N3099, N3034, N2969, N2904, N2839, N2774, N2709, N2644, N2540, N2475, N2346, N2226, N2106, N2033, N1968, N1903, N1838, N1773, N1708, N1643, N1578, N1513, N1409, N1344, N1247, N1182, N1117, N1052, N987, N916, N851, N786, N721, N656, N552, N439, N374, N309, N244, N6326, N6197, N6077, N5957, N5877, N5797, N5732, N5667, N5602, N5537, N5472, N5407, N5342, N5238, N5173, N5076, N5011, N4946, N4867, N4802, N4737, N4672, N4607, N4542, N4477, N4373, N4260, N4147, N4034, N3955, N3890, N3825, N3760, N3695, N3630, N3565, N3500, N3396, N3331, N3266, N3163, N3098, N3033, N2968, N2903, N2838, N2773, N2708, N2643, N2539, N2474, N2345, N2225, N2105, N2032, N1967, N1902, N1837, N1772, N1707, N1642, N1577, N1512, N1408, N1343, N1246, N1181, N1116, N1051, N986, N915, N850, N785, N720, N655, N551, N438, N373, N308, N243, N6325, N6196, N6076, N5956, N5876, N5796, N5731, N5666, N5601, N5536, N5471, N5406, N5341, N5237, N5172, N5075, N5010, N4945, N4866, N4801, N4736, N4671, N4606, N4541, N4476, N4372, N4259, N4146, N4033, N3954, N3889, N3824, N3759, N3694, N3629, N3564, N3499, N3395, N3330, N3265, N3162, N3097, N3032, N2967, N2902, N2837, N2772, N2707, N2642, N2538, N2473, N2344, N2224, N2104, N2031, N1966, N1901, N1836, N1771, N1706, N1641, N1576, N1511, N1407, N1342, N1245, N1180, N1115, N1050, N985, N914, N849, N784, N719, N654, N550, N437, N372, N307, N242, N6324, N6195, N6075, N5955, N5875, N5795, N5730, N5665, N5600, N5535, N5470, N5405, N5340, N5236, N5171, N5074, N5009, N4944, N4865, N4800, N4735, N4670, N4605, N4540, N4475, N4371, N4258, N4145, N4032, N3953, N3888, N3823, N3758, N3693, N3628, N3563, N3498, N3394, N3329, N3264, N3161, N3096, N3031, N2966, N2901, N2836, N2771, N2706, N2641, N2537, N2472, N2343, N2223, N2103, N2030, N1965, N1900, N1835, N1770, N1705, N1640, N1575, N1510, N1406, N1341, N1244, N1179, N1114, N1049, N984, N913, N848, N783, N718, N653, N549, N436, N371, N306, N241, N6323, N6194, N6074, N5954, N5874, N5794, N5729, N5664, N5599, N5534, N5469, N5404, N5339, N5235, N5170, N5073, N5008, N4943, N4864, N4799, N4734, N4669, N4604, N4539, N4474, N4370, N4257, N4144, N4031, N3952, N3887, N3822, N3757, N3692, N3627, N3562, N3497, N3393, N3328, N3263, N3160, N3095, N3030, N2965, N2900, N2835, N2770, N2705, N2640, N2536, N2471, N2342, N2222, N2102, N2029, N1964, N1899, N1834, N1769, N1704, N1639, N1574, N1509, N1405, N1340, N1243, N1178, N1113, N1048, N983, N912, N847, N782, N717, N652, N548, N435, N370, N305, N240, N6322, N6193, N6073, N5953, N5873, N5793, N5728, N5663, N5598, N5533, N5468, N5403, N5338, N5234, N5169, N5072, N5007, N4942, N4863, N4798, N4733, N4668, N4603, N4538, N4473, N4369, N4256, N4143, N4030, N3951, N3886, N3821, N3756, N3691, N3626, N3561, N3496, N3392, N3327, N3262, N3159, N3094, N3029, N2964, N2899, N2834, N2769, N2704, N2639, N2535, N2470, N2341, N2221, N2101, N2028, N1963, N1898, N1833, N1768, N1703, N1638, N1573, N1508, N1404, N1339, N1242, N1177, N1112, N1047, N982, N911, N846, N781, N716, N651, N547, N434, N369, N304, N239, N6321, N6192, N6072, N5952, N5872, N5792, N5727, N5662, N5597, N5532, N5467, N5402, N5337, N5233, N5168, N5071, N5006, N4941, N4862, N4797, N4732, N4667, N4602, N4537, N4472, N4368, N4255, N4142, N4029, N3950, N3885, N3820, N3755, N3690, N3625, N3560, N3495, N3391, N3326, N3261, N3158, N3093, N3028, N2963, N2898, N2833, N2768, N2703, N2638, N2534, N2469, N2340, N2220, N2100, N2027, N1962, N1897, N1832, N1767, N1702, N1637, N1572, N1507, N1403, N1338, N1241, N1176, N1111, N1046, N981, N910, N845, N780, N715, N650, N546, N433, N368, N303, N238, N6320, N6191, N6071, N5951, N5871, N5791, N5726, N5661, N5596, N5531, N5466, N5401, N5336, N5232, N5167, N5070, N5005, N4940, N4861, N4796, N4731, N4666, N4601, N4536, N4471, N4367, N4254, N4141, N4028, N3949, N3884, N3819, N3754, N3689, N3624, N3559, N3494, N3390, N3325, N3260, N3157, N3092, N3027, N2962, N2897, N2832, N2767, N2702, N2637, N2533, N2468, N2339, N2219, N2099, N2026, N1961, N1896, N1831, N1766, N1701, N1636, N1571, N1506, N1402, N1337, N1240, N1175, N1110, N1045, N980, N909, N844, N779, N714, N649, N545, N432, N367, N302, N237, N6319, N6190, N6070, N5950, N5870, N5790, N5725, N5660, N5595, N5530, N5465, N5400, N5335, N5231, N5166, N5069, N5004, N4939, N4860, N4795, N4730, N4665, N4600, N4535, N4470, N4366, N4253, N4140, N4027, N3948, N3883, N3818, N3753, N3688, N3623, N3558, N3493, N3389, N3324, N3259, N3156, N3091, N3026, N2961, N2896, N2831, N2766, N2701, N2636, N2532, N2467, N2338, N2218, N2098, N2025, N1960, N1895, N1830, N1765, N1700, N1635, N1570, N1505, N1401, N1336, N1239, N1174, N1109, N1044, N979, N908, N843, N778, N713, N648, N544, N431, N366, N301, N236, N6318, N6189, N6069, N5949, N5869, N5789, N5724, N5659, N5594, N5529, N5464, N5399, N5334, N5230, N5165, N5068, N5003, N4938, N4859, N4794, N4729, N4664, N4599, N4534, N4469, N4365, N4252, N4139, N4026, N3947, N3882, N3817, N3752, N3687, N3622, N3557, N3492, N3388, N3323, N3258, N3155, N3090, N3025, N2960, N2895, N2830, N2765, N2700, N2635, N2531, N2466, N2337, N2217, N2097, N2024, N1959, N1894, N1829, N1764, N1699, N1634, N1569, N1504, N1400, N1335, N1238, N1173, N1108, N1043, N978, N907, N842, N777, N712, N647, N543, N430, N365, N300, N235, N6317, N6188, N6068, N5948, N5868, N5788, N5723, N5658, N5593, N5528, N5463, N5398, N5333, N5229, N5164, N5067, N5002, N4937, N4858, N4793, N4728, N4663, N4598, N4533, N4468, N4364, N4251, N4138, N4025, N3946, N3881, N3816, N3751, N3686, N3621, N3556, N3491, N3387, N3322, N3257, N3154, N3089, N3024, N2959, N2894, N2829, N2764, N2699, N2634, N2530, N2465, N2336, N2216, N2096, N2023, N1958, N1893, N1828, N1763, N1698, N1633, N1568, N1503, N1399, N1334, N1237, N1172, N1107, N1042, N977, N906, N841, N776, N711, N646, N542, N429, N364, N299, N234, N6316, N6187, N6067, N5947, N5867, N5787, N5722, N5657, N5592, N5527, N5462, N5397, N5332, N5228, N5163, N5066, N5001, N4936, N4857, N4792, N4727, N4662, N4597, N4532, N4467, N4363, N4250, N4137, N4024, N3945, N3880, N3815, N3750, N3685, N3620, N3555, N3490, N3386, N3321, N3256, N3153, N3088, N3023, N2958, N2893, N2828, N2763, N2698, N2633, N2529, N2464, N2335, N2215, N2095, N2022, N1957, N1892, N1827, N1762, N1697, N1632, N1567, N1502, N1398, N1333, N1236, N1171, N1106, N1041, N976, N905, N840, N775, N710, N645, N541, N428, N363, N298, N233, N6315, N6186, N6066, N5946, N5866, N5786, N5721, N5656, N5591, N5526, N5461, N5396, N5331, N5227, N5162, N5065, N5000, N4935, N4856, N4791, N4726, N4661, N4596, N4531, N4466, N4362, N4249, N4136, N4023, N3944, N3879, N3814, N3749, N3684, N3619, N3554, N3489, N3385, N3320, N3255, N3152, N3087, N3022, N2957, N2892, N2827, N2762, N2697, N2632, N2528, N2463, N2334, N2214, N2094, N2021, N1956, N1891, N1826, N1761, N1696, N1631, N1566, N1501, N1397, N1332, N1235, N1170, N1105, N1040, N975, N904, N839, N774, N709, N644, N540, N427, N362, N297, N232, N6314, N6185, N6065, N5945, N5865, N5785, N5720, N5655, N5590, N5525, N5460, N5395, N5330, N5226, N5161, N5064, N4999, N4934, N4855, N4790, N4725, N4660, N4595, N4530, N4465, N4361, N4248, N4135, N4022, N3943, N3878, N3813, N3748, N3683, N3618, N3553, N3488, N3384, N3319, N3254, N3151, N3086, N3021, N2956, N2891, N2826, N2761, N2696, N2631, N2527, N2462, N2333, N2213, N2093, N2020, N1955, N1890, N1825, N1760, N1695, N1630, N1565, N1500, N1396, N1331, N1234, N1169, N1104, N1039, N974, N903, N838, N773, N708, N643, N539, N426, N361, N296, N231, N6313, N6184, N6064, N5944, N5864, N5784, N5719, N5654, N5589, N5524, N5459, N5394, N5329, N5225, N5160, N5063, N4998, N4933, N4854, N4789, N4724, N4659, N4594, N4529, N4464, N4360, N4247, N4134, N4021, N3942, N3877, N3812, N3747, N3682, N3617, N3552, N3487, N3383, N3318, N3253, N3150, N3085, N3020, N2955, N2890, N2825, N2760, N2695, N2630, N2526, N2461, N2332, N2212, N2092, N2019, N1954, N1889, N1824, N1759, N1694, N1629, N1564, N1499, N1395, N1330, N1233, N1168, N1103, N1038, N973, N902, N837, N772, N707, N642, N538, N425, N360, N295, N230 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       (N228)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N96 = N227;
  assign read_en = v_i & N11659;
  assign N11659 = ~w_i;
  assign N97 = ~addr_r[0];
  assign N98 = ~addr_r[1];
  assign N99 = N97 & N98;
  assign N100 = N97 & addr_r[1];
  assign N101 = addr_r[0] & N98;
  assign N102 = addr_r[0] & addr_r[1];
  assign N103 = ~addr_r[2];
  assign N104 = N99 & N103;
  assign N105 = N99 & addr_r[2];
  assign N106 = N101 & N103;
  assign N107 = N101 & addr_r[2];
  assign N108 = N100 & N103;
  assign N109 = N100 & addr_r[2];
  assign N110 = N102 & N103;
  assign N111 = N102 & addr_r[2];
  assign N112 = ~addr_r[3];
  assign N113 = N104 & N112;
  assign N114 = N104 & addr_r[3];
  assign N115 = N106 & N112;
  assign N116 = N106 & addr_r[3];
  assign N117 = N108 & N112;
  assign N118 = N108 & addr_r[3];
  assign N119 = N110 & N112;
  assign N120 = N110 & addr_r[3];
  assign N121 = N105 & N112;
  assign N122 = N105 & addr_r[3];
  assign N123 = N107 & N112;
  assign N124 = N107 & addr_r[3];
  assign N125 = N109 & N112;
  assign N126 = N109 & addr_r[3];
  assign N127 = N111 & N112;
  assign N128 = N111 & addr_r[3];
  assign N129 = ~addr_r[4];
  assign N130 = N113 & N129;
  assign N131 = N113 & addr_r[4];
  assign N132 = N115 & N129;
  assign N133 = N115 & addr_r[4];
  assign N134 = N117 & N129;
  assign N135 = N117 & addr_r[4];
  assign N136 = N119 & N129;
  assign N137 = N119 & addr_r[4];
  assign N138 = N121 & N129;
  assign N139 = N121 & addr_r[4];
  assign N140 = N123 & N129;
  assign N141 = N123 & addr_r[4];
  assign N142 = N125 & N129;
  assign N143 = N125 & addr_r[4];
  assign N144 = N127 & N129;
  assign N145 = N127 & addr_r[4];
  assign N146 = N114 & N129;
  assign N147 = N114 & addr_r[4];
  assign N148 = N116 & N129;
  assign N149 = N116 & addr_r[4];
  assign N150 = N118 & N129;
  assign N151 = N118 & addr_r[4];
  assign N152 = N120 & N129;
  assign N153 = N120 & addr_r[4];
  assign N154 = N122 & N129;
  assign N155 = N122 & addr_r[4];
  assign N156 = N124 & N129;
  assign N157 = N124 & addr_r[4];
  assign N158 = N126 & N129;
  assign N159 = N126 & addr_r[4];
  assign N160 = N128 & N129;
  assign N161 = N128 & addr_r[4];
  assign N162 = ~addr_r[5];
  assign N163 = N130 & N162;
  assign N164 = N130 & addr_r[5];
  assign N165 = N132 & N162;
  assign N166 = N132 & addr_r[5];
  assign N167 = N134 & N162;
  assign N168 = N134 & addr_r[5];
  assign N169 = N136 & N162;
  assign N170 = N136 & addr_r[5];
  assign N171 = N138 & N162;
  assign N172 = N138 & addr_r[5];
  assign N173 = N140 & N162;
  assign N174 = N140 & addr_r[5];
  assign N175 = N142 & N162;
  assign N176 = N142 & addr_r[5];
  assign N177 = N144 & N162;
  assign N178 = N144 & addr_r[5];
  assign N179 = N146 & N162;
  assign N180 = N146 & addr_r[5];
  assign N181 = N148 & N162;
  assign N182 = N148 & addr_r[5];
  assign N183 = N150 & N162;
  assign N184 = N150 & addr_r[5];
  assign N185 = N152 & N162;
  assign N186 = N152 & addr_r[5];
  assign N187 = N154 & N162;
  assign N188 = N154 & addr_r[5];
  assign N189 = N156 & N162;
  assign N190 = N156 & addr_r[5];
  assign N191 = N158 & N162;
  assign N192 = N158 & addr_r[5];
  assign N193 = N160 & N162;
  assign N194 = N160 & addr_r[5];
  assign N195 = N131 & N162;
  assign N196 = N131 & addr_r[5];
  assign N197 = N133 & N162;
  assign N198 = N133 & addr_r[5];
  assign N199 = N135 & N162;
  assign N200 = N135 & addr_r[5];
  assign N201 = N137 & N162;
  assign N202 = N137 & addr_r[5];
  assign N203 = N139 & N162;
  assign N204 = N139 & addr_r[5];
  assign N205 = N141 & N162;
  assign N206 = N141 & addr_r[5];
  assign N207 = N143 & N162;
  assign N208 = N143 & addr_r[5];
  assign N209 = N145 & N162;
  assign N210 = N145 & addr_r[5];
  assign N211 = N147 & N162;
  assign N212 = N147 & addr_r[5];
  assign N213 = N149 & N162;
  assign N214 = N149 & addr_r[5];
  assign N215 = N151 & N162;
  assign N216 = N151 & addr_r[5];
  assign N217 = N153 & N162;
  assign N218 = N153 & addr_r[5];
  assign N219 = N155 & N162;
  assign N220 = N155 & addr_r[5];
  assign N221 = N157 & N162;
  assign N222 = N157 & addr_r[5];
  assign N223 = N159 & N162;
  assign N224 = N159 & addr_r[5];
  assign N225 = N161 & N162;
  assign N226 = N161 & addr_r[5];
  assign N227 = v_i & w_i;
  assign N228 = ~N227;
  assign N229 = ~w_mask_i[0];
  assign N294 = ~w_mask_i[1];
  assign N359 = ~w_mask_i[2];
  assign N424 = ~w_mask_i[3];
  assign N489 = ~w_mask_i[4];
  assign N602 = ~w_mask_i[5];
  assign N706 = ~w_mask_i[6];
  assign N771 = ~w_mask_i[7];
  assign N836 = ~w_mask_i[8];
  assign N901 = ~w_mask_i[9];
  assign N966 = ~w_mask_i[10];
  assign N1037 = ~w_mask_i[11];
  assign N1102 = ~w_mask_i[12];
  assign N1167 = ~w_mask_i[13];
  assign N1232 = ~w_mask_i[14];
  assign N1297 = ~w_mask_i[15];
  assign N1394 = ~w_mask_i[16];
  assign N1459 = ~w_mask_i[17];
  assign N1563 = ~w_mask_i[18];
  assign N1628 = ~w_mask_i[19];
  assign N1693 = ~w_mask_i[20];
  assign N1758 = ~w_mask_i[21];
  assign N1823 = ~w_mask_i[22];
  assign N1888 = ~w_mask_i[23];
  assign N1953 = ~w_mask_i[24];
  assign N2018 = ~w_mask_i[25];
  assign N2083 = ~w_mask_i[26];
  assign N2156 = ~w_mask_i[27];
  assign N2276 = ~w_mask_i[28];
  assign N2396 = ~w_mask_i[29];
  assign N2525 = ~w_mask_i[30];
  assign N2590 = ~w_mask_i[31];
  assign N2694 = ~w_mask_i[32];
  assign N2759 = ~w_mask_i[33];
  assign N2824 = ~w_mask_i[34];
  assign N2889 = ~w_mask_i[35];
  assign N2954 = ~w_mask_i[36];
  assign N3019 = ~w_mask_i[37];
  assign N3084 = ~w_mask_i[38];
  assign N3149 = ~w_mask_i[39];
  assign N3214 = ~w_mask_i[40];
  assign N3317 = ~w_mask_i[41];
  assign N3382 = ~w_mask_i[42];
  assign N3447 = ~w_mask_i[43];
  assign N3551 = ~w_mask_i[44];
  assign N3616 = ~w_mask_i[45];
  assign N3681 = ~w_mask_i[46];
  assign N3746 = ~w_mask_i[47];
  assign N3811 = ~w_mask_i[48];
  assign N3876 = ~w_mask_i[49];
  assign N3941 = ~w_mask_i[50];
  assign N4006 = ~w_mask_i[51];
  assign N4085 = ~w_mask_i[52];
  assign N4198 = ~w_mask_i[53];
  assign N4311 = ~w_mask_i[54];
  assign N4424 = ~w_mask_i[55];
  assign N4528 = ~w_mask_i[56];
  assign N4593 = ~w_mask_i[57];
  assign N4658 = ~w_mask_i[58];
  assign N4723 = ~w_mask_i[59];
  assign N4788 = ~w_mask_i[60];
  assign N4853 = ~w_mask_i[61];
  assign N4918 = ~w_mask_i[62];
  assign N4997 = ~w_mask_i[63];
  assign N5062 = ~w_mask_i[64];
  assign N5127 = ~w_mask_i[65];
  assign N5224 = ~w_mask_i[66];
  assign N5289 = ~w_mask_i[67];
  assign N5393 = ~w_mask_i[68];
  assign N5458 = ~w_mask_i[69];
  assign N5523 = ~w_mask_i[70];
  assign N5588 = ~w_mask_i[71];
  assign N5653 = ~w_mask_i[72];
  assign N5718 = ~w_mask_i[73];
  assign N5783 = ~w_mask_i[74];
  assign N5848 = ~w_mask_i[75];
  assign N5928 = ~w_mask_i[76];
  assign N6008 = ~w_mask_i[77];
  assign N6128 = ~w_mask_i[78];
  assign N6248 = ~w_mask_i[79];

  always @(posedge clk_i) begin
    if(1'b1) begin
      { addr_r[5:0] } <= { addr_i[5:0] };
    end 
    if(N11496) begin
      { mem[5119:5119] } <= { data_i[79:79] };
    end 
    if(N11495) begin
      { mem[5118:5118] } <= { data_i[78:78] };
    end 
    if(N11494) begin
      { mem[5117:5117] } <= { data_i[77:77] };
    end 
    if(N11493) begin
      { mem[5116:5116] } <= { data_i[76:76] };
    end 
    if(N11492) begin
      { mem[5115:5115] } <= { data_i[75:75] };
    end 
    if(N11491) begin
      { mem[5114:5114] } <= { data_i[74:74] };
    end 
    if(N11490) begin
      { mem[5113:5113] } <= { data_i[73:73] };
    end 
    if(N11489) begin
      { mem[5112:5112] } <= { data_i[72:72] };
    end 
    if(N11488) begin
      { mem[5111:5111] } <= { data_i[71:71] };
    end 
    if(N11487) begin
      { mem[5110:5110] } <= { data_i[70:70] };
    end 
    if(N11486) begin
      { mem[5109:5109] } <= { data_i[69:69] };
    end 
    if(N11485) begin
      { mem[5108:5108] } <= { data_i[68:68] };
    end 
    if(N11484) begin
      { mem[5107:5107] } <= { data_i[67:67] };
    end 
    if(N11483) begin
      { mem[5106:5106] } <= { data_i[66:66] };
    end 
    if(N11482) begin
      { mem[5105:5105] } <= { data_i[65:65] };
    end 
    if(N11481) begin
      { mem[5104:5104] } <= { data_i[64:64] };
    end 
    if(N11480) begin
      { mem[5103:5103] } <= { data_i[63:63] };
    end 
    if(N11479) begin
      { mem[5102:5102] } <= { data_i[62:62] };
    end 
    if(N11478) begin
      { mem[5101:5101] } <= { data_i[61:61] };
    end 
    if(N11477) begin
      { mem[5100:5100] } <= { data_i[60:60] };
    end 
    if(N11476) begin
      { mem[5099:5099] } <= { data_i[59:59] };
    end 
    if(N11475) begin
      { mem[5098:5098] } <= { data_i[58:58] };
    end 
    if(N11474) begin
      { mem[5097:5097] } <= { data_i[57:57] };
    end 
    if(N11473) begin
      { mem[5096:5096] } <= { data_i[56:56] };
    end 
    if(N11472) begin
      { mem[5095:5095] } <= { data_i[55:55] };
    end 
    if(N11471) begin
      { mem[5094:5094] } <= { data_i[54:54] };
    end 
    if(N11470) begin
      { mem[5093:5093] } <= { data_i[53:53] };
    end 
    if(N11469) begin
      { mem[5092:5092] } <= { data_i[52:52] };
    end 
    if(N11468) begin
      { mem[5091:5091] } <= { data_i[51:51] };
    end 
    if(N11467) begin
      { mem[5090:5090] } <= { data_i[50:50] };
    end 
    if(N11466) begin
      { mem[5089:5089] } <= { data_i[49:49] };
    end 
    if(N11465) begin
      { mem[5088:5088] } <= { data_i[48:48] };
    end 
    if(N11464) begin
      { mem[5087:5087] } <= { data_i[47:47] };
    end 
    if(N11463) begin
      { mem[5086:5086] } <= { data_i[46:46] };
    end 
    if(N11462) begin
      { mem[5085:5085] } <= { data_i[45:45] };
    end 
    if(N11461) begin
      { mem[5084:5084] } <= { data_i[44:44] };
    end 
    if(N11460) begin
      { mem[5083:5083] } <= { data_i[43:43] };
    end 
    if(N11459) begin
      { mem[5082:5082] } <= { data_i[42:42] };
    end 
    if(N11458) begin
      { mem[5081:5081] } <= { data_i[41:41] };
    end 
    if(N11457) begin
      { mem[5080:5080] } <= { data_i[40:40] };
    end 
    if(N11456) begin
      { mem[5079:5079] } <= { data_i[39:39] };
    end 
    if(N11455) begin
      { mem[5078:5078] } <= { data_i[38:38] };
    end 
    if(N11454) begin
      { mem[5077:5077] } <= { data_i[37:37] };
    end 
    if(N11453) begin
      { mem[5076:5076] } <= { data_i[36:36] };
    end 
    if(N11452) begin
      { mem[5075:5075] } <= { data_i[35:35] };
    end 
    if(N11451) begin
      { mem[5074:5074] } <= { data_i[34:34] };
    end 
    if(N11450) begin
      { mem[5073:5073] } <= { data_i[33:33] };
    end 
    if(N11449) begin
      { mem[5072:5072] } <= { data_i[32:32] };
    end 
    if(N11448) begin
      { mem[5071:5071] } <= { data_i[31:31] };
    end 
    if(N11447) begin
      { mem[5070:5070] } <= { data_i[30:30] };
    end 
    if(N11446) begin
      { mem[5069:5069] } <= { data_i[29:29] };
    end 
    if(N11445) begin
      { mem[5068:5068] } <= { data_i[28:28] };
    end 
    if(N11444) begin
      { mem[5067:5067] } <= { data_i[27:27] };
    end 
    if(N11443) begin
      { mem[5066:5066] } <= { data_i[26:26] };
    end 
    if(N11442) begin
      { mem[5065:5065] } <= { data_i[25:25] };
    end 
    if(N11441) begin
      { mem[5064:5064] } <= { data_i[24:24] };
    end 
    if(N11440) begin
      { mem[5063:5063] } <= { data_i[23:23] };
    end 
    if(N11439) begin
      { mem[5062:5062] } <= { data_i[22:22] };
    end 
    if(N11438) begin
      { mem[5061:5061] } <= { data_i[21:21] };
    end 
    if(N11437) begin
      { mem[5060:5060] } <= { data_i[20:20] };
    end 
    if(N11436) begin
      { mem[5059:5059] } <= { data_i[19:19] };
    end 
    if(N11435) begin
      { mem[5058:5058] } <= { data_i[18:18] };
    end 
    if(N11434) begin
      { mem[5057:5057] } <= { data_i[17:17] };
    end 
    if(N11433) begin
      { mem[5056:5056] } <= { data_i[16:16] };
    end 
    if(N11432) begin
      { mem[5055:5055] } <= { data_i[15:15] };
    end 
    if(N11431) begin
      { mem[5054:5054] } <= { data_i[14:14] };
    end 
    if(N11430) begin
      { mem[5053:5053] } <= { data_i[13:13] };
    end 
    if(N11429) begin
      { mem[5052:5052] } <= { data_i[12:12] };
    end 
    if(N11428) begin
      { mem[5051:5051] } <= { data_i[11:11] };
    end 
    if(N11427) begin
      { mem[5050:5050] } <= { data_i[10:10] };
    end 
    if(N11426) begin
      { mem[5049:5049] } <= { data_i[9:9] };
    end 
    if(N11425) begin
      { mem[5048:5048] } <= { data_i[8:8] };
    end 
    if(N11424) begin
      { mem[5047:5047] } <= { data_i[7:7] };
    end 
    if(N11423) begin
      { mem[5046:5046] } <= { data_i[6:6] };
    end 
    if(N11422) begin
      { mem[5045:5045] } <= { data_i[5:5] };
    end 
    if(N11421) begin
      { mem[5044:5044] } <= { data_i[4:4] };
    end 
    if(N11420) begin
      { mem[5043:5043] } <= { data_i[3:3] };
    end 
    if(N11419) begin
      { mem[5042:5042] } <= { data_i[2:2] };
    end 
    if(N11418) begin
      { mem[5041:5041] } <= { data_i[1:1] };
    end 
    if(N11417) begin
      { mem[5040:5040] } <= { data_i[0:0] };
    end 
    if(N11416) begin
      { mem[5039:5039] } <= { data_i[79:79] };
    end 
    if(N11415) begin
      { mem[5038:5038] } <= { data_i[78:78] };
    end 
    if(N11414) begin
      { mem[5037:5037] } <= { data_i[77:77] };
    end 
    if(N11413) begin
      { mem[5036:5036] } <= { data_i[76:76] };
    end 
    if(N11412) begin
      { mem[5035:5035] } <= { data_i[75:75] };
    end 
    if(N11411) begin
      { mem[5034:5034] } <= { data_i[74:74] };
    end 
    if(N11410) begin
      { mem[5033:5033] } <= { data_i[73:73] };
    end 
    if(N11409) begin
      { mem[5032:5032] } <= { data_i[72:72] };
    end 
    if(N11408) begin
      { mem[5031:5031] } <= { data_i[71:71] };
    end 
    if(N11407) begin
      { mem[5030:5030] } <= { data_i[70:70] };
    end 
    if(N11406) begin
      { mem[5029:5029] } <= { data_i[69:69] };
    end 
    if(N11405) begin
      { mem[5028:5028] } <= { data_i[68:68] };
    end 
    if(N11404) begin
      { mem[5027:5027] } <= { data_i[67:67] };
    end 
    if(N11403) begin
      { mem[5026:5026] } <= { data_i[66:66] };
    end 
    if(N11402) begin
      { mem[5025:5025] } <= { data_i[65:65] };
    end 
    if(N11401) begin
      { mem[5024:5024] } <= { data_i[64:64] };
    end 
    if(N11400) begin
      { mem[5023:5023] } <= { data_i[63:63] };
    end 
    if(N11399) begin
      { mem[5022:5022] } <= { data_i[62:62] };
    end 
    if(N11398) begin
      { mem[5021:5021] } <= { data_i[61:61] };
    end 
    if(N11397) begin
      { mem[5020:5020] } <= { data_i[60:60] };
    end 
    if(N11396) begin
      { mem[5019:5019] } <= { data_i[59:59] };
    end 
    if(N11395) begin
      { mem[5018:5018] } <= { data_i[58:58] };
    end 
    if(N11394) begin
      { mem[5017:5017] } <= { data_i[57:57] };
    end 
    if(N11393) begin
      { mem[5016:5016] } <= { data_i[56:56] };
    end 
    if(N11392) begin
      { mem[5015:5015] } <= { data_i[55:55] };
    end 
    if(N11391) begin
      { mem[5014:5014] } <= { data_i[54:54] };
    end 
    if(N11390) begin
      { mem[5013:5013] } <= { data_i[53:53] };
    end 
    if(N11389) begin
      { mem[5012:5012] } <= { data_i[52:52] };
    end 
    if(N11388) begin
      { mem[5011:5011] } <= { data_i[51:51] };
    end 
    if(N11387) begin
      { mem[5010:5010] } <= { data_i[50:50] };
    end 
    if(N11386) begin
      { mem[5009:5009] } <= { data_i[49:49] };
    end 
    if(N11385) begin
      { mem[5008:5008] } <= { data_i[48:48] };
    end 
    if(N11384) begin
      { mem[5007:5007] } <= { data_i[47:47] };
    end 
    if(N11383) begin
      { mem[5006:5006] } <= { data_i[46:46] };
    end 
    if(N11382) begin
      { mem[5005:5005] } <= { data_i[45:45] };
    end 
    if(N11381) begin
      { mem[5004:5004] } <= { data_i[44:44] };
    end 
    if(N11380) begin
      { mem[5003:5003] } <= { data_i[43:43] };
    end 
    if(N11379) begin
      { mem[5002:5002] } <= { data_i[42:42] };
    end 
    if(N11378) begin
      { mem[5001:5001] } <= { data_i[41:41] };
    end 
    if(N11377) begin
      { mem[5000:5000] } <= { data_i[40:40] };
    end 
    if(N11376) begin
      { mem[4999:4999] } <= { data_i[39:39] };
    end 
    if(N11375) begin
      { mem[4998:4998] } <= { data_i[38:38] };
    end 
    if(N11374) begin
      { mem[4997:4997] } <= { data_i[37:37] };
    end 
    if(N11373) begin
      { mem[4996:4996] } <= { data_i[36:36] };
    end 
    if(N11372) begin
      { mem[4995:4995] } <= { data_i[35:35] };
    end 
    if(N11371) begin
      { mem[4994:4994] } <= { data_i[34:34] };
    end 
    if(N11370) begin
      { mem[4993:4993] } <= { data_i[33:33] };
    end 
    if(N11369) begin
      { mem[4992:4992] } <= { data_i[32:32] };
    end 
    if(N11368) begin
      { mem[4991:4991] } <= { data_i[31:31] };
    end 
    if(N11367) begin
      { mem[4990:4990] } <= { data_i[30:30] };
    end 
    if(N11366) begin
      { mem[4989:4989] } <= { data_i[29:29] };
    end 
    if(N11365) begin
      { mem[4988:4988] } <= { data_i[28:28] };
    end 
    if(N11364) begin
      { mem[4987:4987] } <= { data_i[27:27] };
    end 
    if(N11363) begin
      { mem[4986:4986] } <= { data_i[26:26] };
    end 
    if(N11362) begin
      { mem[4985:4985] } <= { data_i[25:25] };
    end 
    if(N11361) begin
      { mem[4984:4984] } <= { data_i[24:24] };
    end 
    if(N11360) begin
      { mem[4983:4983] } <= { data_i[23:23] };
    end 
    if(N11359) begin
      { mem[4982:4982] } <= { data_i[22:22] };
    end 
    if(N11358) begin
      { mem[4981:4981] } <= { data_i[21:21] };
    end 
    if(N11357) begin
      { mem[4980:4980] } <= { data_i[20:20] };
    end 
    if(N11356) begin
      { mem[4979:4979] } <= { data_i[19:19] };
    end 
    if(N11355) begin
      { mem[4978:4978] } <= { data_i[18:18] };
    end 
    if(N11354) begin
      { mem[4977:4977] } <= { data_i[17:17] };
    end 
    if(N11353) begin
      { mem[4976:4976] } <= { data_i[16:16] };
    end 
    if(N11352) begin
      { mem[4975:4975] } <= { data_i[15:15] };
    end 
    if(N11351) begin
      { mem[4974:4974] } <= { data_i[14:14] };
    end 
    if(N11350) begin
      { mem[4973:4973] } <= { data_i[13:13] };
    end 
    if(N11349) begin
      { mem[4972:4972] } <= { data_i[12:12] };
    end 
    if(N11348) begin
      { mem[4971:4971] } <= { data_i[11:11] };
    end 
    if(N11347) begin
      { mem[4970:4970] } <= { data_i[10:10] };
    end 
    if(N11346) begin
      { mem[4969:4969] } <= { data_i[9:9] };
    end 
    if(N11345) begin
      { mem[4968:4968] } <= { data_i[8:8] };
    end 
    if(N11344) begin
      { mem[4967:4967] } <= { data_i[7:7] };
    end 
    if(N11343) begin
      { mem[4966:4966] } <= { data_i[6:6] };
    end 
    if(N11342) begin
      { mem[4965:4965] } <= { data_i[5:5] };
    end 
    if(N11341) begin
      { mem[4964:4964] } <= { data_i[4:4] };
    end 
    if(N11340) begin
      { mem[4963:4963] } <= { data_i[3:3] };
    end 
    if(N11339) begin
      { mem[4962:4962] } <= { data_i[2:2] };
    end 
    if(N11338) begin
      { mem[4961:4961] } <= { data_i[1:1] };
    end 
    if(N11337) begin
      { mem[4960:4960] } <= { data_i[0:0] };
    end 
    if(N11336) begin
      { mem[4959:4959] } <= { data_i[79:79] };
    end 
    if(N11335) begin
      { mem[4958:4958] } <= { data_i[78:78] };
    end 
    if(N11334) begin
      { mem[4957:4957] } <= { data_i[77:77] };
    end 
    if(N11333) begin
      { mem[4956:4956] } <= { data_i[76:76] };
    end 
    if(N11332) begin
      { mem[4955:4955] } <= { data_i[75:75] };
    end 
    if(N11331) begin
      { mem[4954:4954] } <= { data_i[74:74] };
    end 
    if(N11330) begin
      { mem[4953:4953] } <= { data_i[73:73] };
    end 
    if(N11329) begin
      { mem[4952:4952] } <= { data_i[72:72] };
    end 
    if(N11328) begin
      { mem[4951:4951] } <= { data_i[71:71] };
    end 
    if(N11327) begin
      { mem[4950:4950] } <= { data_i[70:70] };
    end 
    if(N11326) begin
      { mem[4949:4949] } <= { data_i[69:69] };
    end 
    if(N11325) begin
      { mem[4948:4948] } <= { data_i[68:68] };
    end 
    if(N11324) begin
      { mem[4947:4947] } <= { data_i[67:67] };
    end 
    if(N11323) begin
      { mem[4946:4946] } <= { data_i[66:66] };
    end 
    if(N11322) begin
      { mem[4945:4945] } <= { data_i[65:65] };
    end 
    if(N11321) begin
      { mem[4944:4944] } <= { data_i[64:64] };
    end 
    if(N11320) begin
      { mem[4943:4943] } <= { data_i[63:63] };
    end 
    if(N11319) begin
      { mem[4942:4942] } <= { data_i[62:62] };
    end 
    if(N11318) begin
      { mem[4941:4941] } <= { data_i[61:61] };
    end 
    if(N11317) begin
      { mem[4940:4940] } <= { data_i[60:60] };
    end 
    if(N11316) begin
      { mem[4939:4939] } <= { data_i[59:59] };
    end 
    if(N11315) begin
      { mem[4938:4938] } <= { data_i[58:58] };
    end 
    if(N11314) begin
      { mem[4937:4937] } <= { data_i[57:57] };
    end 
    if(N11313) begin
      { mem[4936:4936] } <= { data_i[56:56] };
    end 
    if(N11312) begin
      { mem[4935:4935] } <= { data_i[55:55] };
    end 
    if(N11311) begin
      { mem[4934:4934] } <= { data_i[54:54] };
    end 
    if(N11310) begin
      { mem[4933:4933] } <= { data_i[53:53] };
    end 
    if(N11309) begin
      { mem[4932:4932] } <= { data_i[52:52] };
    end 
    if(N11308) begin
      { mem[4931:4931] } <= { data_i[51:51] };
    end 
    if(N11307) begin
      { mem[4930:4930] } <= { data_i[50:50] };
    end 
    if(N11306) begin
      { mem[4929:4929] } <= { data_i[49:49] };
    end 
    if(N11305) begin
      { mem[4928:4928] } <= { data_i[48:48] };
    end 
    if(N11304) begin
      { mem[4927:4927] } <= { data_i[47:47] };
    end 
    if(N11303) begin
      { mem[4926:4926] } <= { data_i[46:46] };
    end 
    if(N11302) begin
      { mem[4925:4925] } <= { data_i[45:45] };
    end 
    if(N11301) begin
      { mem[4924:4924] } <= { data_i[44:44] };
    end 
    if(N11300) begin
      { mem[4923:4923] } <= { data_i[43:43] };
    end 
    if(N11299) begin
      { mem[4922:4922] } <= { data_i[42:42] };
    end 
    if(N11298) begin
      { mem[4921:4921] } <= { data_i[41:41] };
    end 
    if(N11297) begin
      { mem[4920:4920] } <= { data_i[40:40] };
    end 
    if(N11296) begin
      { mem[4919:4919] } <= { data_i[39:39] };
    end 
    if(N11295) begin
      { mem[4918:4918] } <= { data_i[38:38] };
    end 
    if(N11294) begin
      { mem[4917:4917] } <= { data_i[37:37] };
    end 
    if(N11293) begin
      { mem[4916:4916] } <= { data_i[36:36] };
    end 
    if(N11292) begin
      { mem[4915:4915] } <= { data_i[35:35] };
    end 
    if(N11291) begin
      { mem[4914:4914] } <= { data_i[34:34] };
    end 
    if(N11290) begin
      { mem[4913:4913] } <= { data_i[33:33] };
    end 
    if(N11289) begin
      { mem[4912:4912] } <= { data_i[32:32] };
    end 
    if(N11288) begin
      { mem[4911:4911] } <= { data_i[31:31] };
    end 
    if(N11287) begin
      { mem[4910:4910] } <= { data_i[30:30] };
    end 
    if(N11286) begin
      { mem[4909:4909] } <= { data_i[29:29] };
    end 
    if(N11285) begin
      { mem[4908:4908] } <= { data_i[28:28] };
    end 
    if(N11284) begin
      { mem[4907:4907] } <= { data_i[27:27] };
    end 
    if(N11283) begin
      { mem[4906:4906] } <= { data_i[26:26] };
    end 
    if(N11282) begin
      { mem[4905:4905] } <= { data_i[25:25] };
    end 
    if(N11281) begin
      { mem[4904:4904] } <= { data_i[24:24] };
    end 
    if(N11280) begin
      { mem[4903:4903] } <= { data_i[23:23] };
    end 
    if(N11279) begin
      { mem[4902:4902] } <= { data_i[22:22] };
    end 
    if(N11278) begin
      { mem[4901:4901] } <= { data_i[21:21] };
    end 
    if(N11277) begin
      { mem[4900:4900] } <= { data_i[20:20] };
    end 
    if(N11276) begin
      { mem[4899:4899] } <= { data_i[19:19] };
    end 
    if(N11275) begin
      { mem[4898:4898] } <= { data_i[18:18] };
    end 
    if(N11274) begin
      { mem[4897:4897] } <= { data_i[17:17] };
    end 
    if(N11273) begin
      { mem[4896:4896] } <= { data_i[16:16] };
    end 
    if(N11272) begin
      { mem[4895:4895] } <= { data_i[15:15] };
    end 
    if(N11271) begin
      { mem[4894:4894] } <= { data_i[14:14] };
    end 
    if(N11270) begin
      { mem[4893:4893] } <= { data_i[13:13] };
    end 
    if(N11269) begin
      { mem[4892:4892] } <= { data_i[12:12] };
    end 
    if(N11268) begin
      { mem[4891:4891] } <= { data_i[11:11] };
    end 
    if(N11267) begin
      { mem[4890:4890] } <= { data_i[10:10] };
    end 
    if(N11266) begin
      { mem[4889:4889] } <= { data_i[9:9] };
    end 
    if(N11265) begin
      { mem[4888:4888] } <= { data_i[8:8] };
    end 
    if(N11264) begin
      { mem[4887:4887] } <= { data_i[7:7] };
    end 
    if(N11263) begin
      { mem[4886:4886] } <= { data_i[6:6] };
    end 
    if(N11262) begin
      { mem[4885:4885] } <= { data_i[5:5] };
    end 
    if(N11261) begin
      { mem[4884:4884] } <= { data_i[4:4] };
    end 
    if(N11260) begin
      { mem[4883:4883] } <= { data_i[3:3] };
    end 
    if(N11259) begin
      { mem[4882:4882] } <= { data_i[2:2] };
    end 
    if(N11258) begin
      { mem[4881:4881] } <= { data_i[1:1] };
    end 
    if(N11257) begin
      { mem[4880:4880] } <= { data_i[0:0] };
    end 
    if(N11256) begin
      { mem[4879:4879] } <= { data_i[79:79] };
    end 
    if(N11255) begin
      { mem[4878:4878] } <= { data_i[78:78] };
    end 
    if(N11254) begin
      { mem[4877:4877] } <= { data_i[77:77] };
    end 
    if(N11253) begin
      { mem[4876:4876] } <= { data_i[76:76] };
    end 
    if(N11252) begin
      { mem[4875:4875] } <= { data_i[75:75] };
    end 
    if(N11251) begin
      { mem[4874:4874] } <= { data_i[74:74] };
    end 
    if(N11250) begin
      { mem[4873:4873] } <= { data_i[73:73] };
    end 
    if(N11249) begin
      { mem[4872:4872] } <= { data_i[72:72] };
    end 
    if(N11248) begin
      { mem[4871:4871] } <= { data_i[71:71] };
    end 
    if(N11247) begin
      { mem[4870:4870] } <= { data_i[70:70] };
    end 
    if(N11246) begin
      { mem[4869:4869] } <= { data_i[69:69] };
    end 
    if(N11245) begin
      { mem[4868:4868] } <= { data_i[68:68] };
    end 
    if(N11244) begin
      { mem[4867:4867] } <= { data_i[67:67] };
    end 
    if(N11243) begin
      { mem[4866:4866] } <= { data_i[66:66] };
    end 
    if(N11242) begin
      { mem[4865:4865] } <= { data_i[65:65] };
    end 
    if(N11241) begin
      { mem[4864:4864] } <= { data_i[64:64] };
    end 
    if(N11240) begin
      { mem[4863:4863] } <= { data_i[63:63] };
    end 
    if(N11239) begin
      { mem[4862:4862] } <= { data_i[62:62] };
    end 
    if(N11238) begin
      { mem[4861:4861] } <= { data_i[61:61] };
    end 
    if(N11237) begin
      { mem[4860:4860] } <= { data_i[60:60] };
    end 
    if(N11236) begin
      { mem[4859:4859] } <= { data_i[59:59] };
    end 
    if(N11235) begin
      { mem[4858:4858] } <= { data_i[58:58] };
    end 
    if(N11234) begin
      { mem[4857:4857] } <= { data_i[57:57] };
    end 
    if(N11233) begin
      { mem[4856:4856] } <= { data_i[56:56] };
    end 
    if(N11232) begin
      { mem[4855:4855] } <= { data_i[55:55] };
    end 
    if(N11231) begin
      { mem[4854:4854] } <= { data_i[54:54] };
    end 
    if(N11230) begin
      { mem[4853:4853] } <= { data_i[53:53] };
    end 
    if(N11229) begin
      { mem[4852:4852] } <= { data_i[52:52] };
    end 
    if(N11228) begin
      { mem[4851:4851] } <= { data_i[51:51] };
    end 
    if(N11227) begin
      { mem[4850:4850] } <= { data_i[50:50] };
    end 
    if(N11226) begin
      { mem[4849:4849] } <= { data_i[49:49] };
    end 
    if(N11225) begin
      { mem[4848:4848] } <= { data_i[48:48] };
    end 
    if(N11224) begin
      { mem[4847:4847] } <= { data_i[47:47] };
    end 
    if(N11223) begin
      { mem[4846:4846] } <= { data_i[46:46] };
    end 
    if(N11222) begin
      { mem[4845:4845] } <= { data_i[45:45] };
    end 
    if(N11221) begin
      { mem[4844:4844] } <= { data_i[44:44] };
    end 
    if(N11220) begin
      { mem[4843:4843] } <= { data_i[43:43] };
    end 
    if(N11219) begin
      { mem[4842:4842] } <= { data_i[42:42] };
    end 
    if(N11218) begin
      { mem[4841:4841] } <= { data_i[41:41] };
    end 
    if(N11217) begin
      { mem[4840:4840] } <= { data_i[40:40] };
    end 
    if(N11216) begin
      { mem[4839:4839] } <= { data_i[39:39] };
    end 
    if(N11215) begin
      { mem[4838:4838] } <= { data_i[38:38] };
    end 
    if(N11214) begin
      { mem[4837:4837] } <= { data_i[37:37] };
    end 
    if(N11213) begin
      { mem[4836:4836] } <= { data_i[36:36] };
    end 
    if(N11212) begin
      { mem[4835:4835] } <= { data_i[35:35] };
    end 
    if(N11211) begin
      { mem[4834:4834] } <= { data_i[34:34] };
    end 
    if(N11210) begin
      { mem[4833:4833] } <= { data_i[33:33] };
    end 
    if(N11209) begin
      { mem[4832:4832] } <= { data_i[32:32] };
    end 
    if(N11208) begin
      { mem[4831:4831] } <= { data_i[31:31] };
    end 
    if(N11207) begin
      { mem[4830:4830] } <= { data_i[30:30] };
    end 
    if(N11206) begin
      { mem[4829:4829] } <= { data_i[29:29] };
    end 
    if(N11205) begin
      { mem[4828:4828] } <= { data_i[28:28] };
    end 
    if(N11204) begin
      { mem[4827:4827] } <= { data_i[27:27] };
    end 
    if(N11203) begin
      { mem[4826:4826] } <= { data_i[26:26] };
    end 
    if(N11202) begin
      { mem[4825:4825] } <= { data_i[25:25] };
    end 
    if(N11201) begin
      { mem[4824:4824] } <= { data_i[24:24] };
    end 
    if(N11200) begin
      { mem[4823:4823] } <= { data_i[23:23] };
    end 
    if(N11199) begin
      { mem[4822:4822] } <= { data_i[22:22] };
    end 
    if(N11198) begin
      { mem[4821:4821] } <= { data_i[21:21] };
    end 
    if(N11197) begin
      { mem[4820:4820] } <= { data_i[20:20] };
    end 
    if(N11196) begin
      { mem[4819:4819] } <= { data_i[19:19] };
    end 
    if(N11195) begin
      { mem[4818:4818] } <= { data_i[18:18] };
    end 
    if(N11194) begin
      { mem[4817:4817] } <= { data_i[17:17] };
    end 
    if(N11193) begin
      { mem[4816:4816] } <= { data_i[16:16] };
    end 
    if(N11192) begin
      { mem[4815:4815] } <= { data_i[15:15] };
    end 
    if(N11191) begin
      { mem[4814:4814] } <= { data_i[14:14] };
    end 
    if(N11190) begin
      { mem[4813:4813] } <= { data_i[13:13] };
    end 
    if(N11189) begin
      { mem[4812:4812] } <= { data_i[12:12] };
    end 
    if(N11188) begin
      { mem[4811:4811] } <= { data_i[11:11] };
    end 
    if(N11187) begin
      { mem[4810:4810] } <= { data_i[10:10] };
    end 
    if(N11186) begin
      { mem[4809:4809] } <= { data_i[9:9] };
    end 
    if(N11185) begin
      { mem[4808:4808] } <= { data_i[8:8] };
    end 
    if(N11184) begin
      { mem[4807:4807] } <= { data_i[7:7] };
    end 
    if(N11183) begin
      { mem[4806:4806] } <= { data_i[6:6] };
    end 
    if(N11182) begin
      { mem[4805:4805] } <= { data_i[5:5] };
    end 
    if(N11181) begin
      { mem[4804:4804] } <= { data_i[4:4] };
    end 
    if(N11180) begin
      { mem[4803:4803] } <= { data_i[3:3] };
    end 
    if(N11179) begin
      { mem[4802:4802] } <= { data_i[2:2] };
    end 
    if(N11178) begin
      { mem[4801:4801] } <= { data_i[1:1] };
    end 
    if(N11177) begin
      { mem[4800:4800] } <= { data_i[0:0] };
    end 
    if(N11176) begin
      { mem[4799:4799] } <= { data_i[79:79] };
    end 
    if(N11175) begin
      { mem[4798:4798] } <= { data_i[78:78] };
    end 
    if(N11174) begin
      { mem[4797:4797] } <= { data_i[77:77] };
    end 
    if(N11173) begin
      { mem[4796:4796] } <= { data_i[76:76] };
    end 
    if(N11172) begin
      { mem[4795:4795] } <= { data_i[75:75] };
    end 
    if(N11171) begin
      { mem[4794:4794] } <= { data_i[74:74] };
    end 
    if(N11170) begin
      { mem[4793:4793] } <= { data_i[73:73] };
    end 
    if(N11169) begin
      { mem[4792:4792] } <= { data_i[72:72] };
    end 
    if(N11168) begin
      { mem[4791:4791] } <= { data_i[71:71] };
    end 
    if(N11167) begin
      { mem[4790:4790] } <= { data_i[70:70] };
    end 
    if(N11166) begin
      { mem[4789:4789] } <= { data_i[69:69] };
    end 
    if(N11165) begin
      { mem[4788:4788] } <= { data_i[68:68] };
    end 
    if(N11164) begin
      { mem[4787:4787] } <= { data_i[67:67] };
    end 
    if(N11163) begin
      { mem[4786:4786] } <= { data_i[66:66] };
    end 
    if(N11162) begin
      { mem[4785:4785] } <= { data_i[65:65] };
    end 
    if(N11161) begin
      { mem[4784:4784] } <= { data_i[64:64] };
    end 
    if(N11160) begin
      { mem[4783:4783] } <= { data_i[63:63] };
    end 
    if(N11159) begin
      { mem[4782:4782] } <= { data_i[62:62] };
    end 
    if(N11158) begin
      { mem[4781:4781] } <= { data_i[61:61] };
    end 
    if(N11157) begin
      { mem[4780:4780] } <= { data_i[60:60] };
    end 
    if(N11156) begin
      { mem[4779:4779] } <= { data_i[59:59] };
    end 
    if(N11155) begin
      { mem[4778:4778] } <= { data_i[58:58] };
    end 
    if(N11154) begin
      { mem[4777:4777] } <= { data_i[57:57] };
    end 
    if(N11153) begin
      { mem[4776:4776] } <= { data_i[56:56] };
    end 
    if(N11152) begin
      { mem[4775:4775] } <= { data_i[55:55] };
    end 
    if(N11151) begin
      { mem[4774:4774] } <= { data_i[54:54] };
    end 
    if(N11150) begin
      { mem[4773:4773] } <= { data_i[53:53] };
    end 
    if(N11149) begin
      { mem[4772:4772] } <= { data_i[52:52] };
    end 
    if(N11148) begin
      { mem[4771:4771] } <= { data_i[51:51] };
    end 
    if(N11147) begin
      { mem[4770:4770] } <= { data_i[50:50] };
    end 
    if(N11146) begin
      { mem[4769:4769] } <= { data_i[49:49] };
    end 
    if(N11145) begin
      { mem[4768:4768] } <= { data_i[48:48] };
    end 
    if(N11144) begin
      { mem[4767:4767] } <= { data_i[47:47] };
    end 
    if(N11143) begin
      { mem[4766:4766] } <= { data_i[46:46] };
    end 
    if(N11142) begin
      { mem[4765:4765] } <= { data_i[45:45] };
    end 
    if(N11141) begin
      { mem[4764:4764] } <= { data_i[44:44] };
    end 
    if(N11140) begin
      { mem[4763:4763] } <= { data_i[43:43] };
    end 
    if(N11139) begin
      { mem[4762:4762] } <= { data_i[42:42] };
    end 
    if(N11138) begin
      { mem[4761:4761] } <= { data_i[41:41] };
    end 
    if(N11137) begin
      { mem[4760:4760] } <= { data_i[40:40] };
    end 
    if(N11136) begin
      { mem[4759:4759] } <= { data_i[39:39] };
    end 
    if(N11135) begin
      { mem[4758:4758] } <= { data_i[38:38] };
    end 
    if(N11134) begin
      { mem[4757:4757] } <= { data_i[37:37] };
    end 
    if(N11133) begin
      { mem[4756:4756] } <= { data_i[36:36] };
    end 
    if(N11132) begin
      { mem[4755:4755] } <= { data_i[35:35] };
    end 
    if(N11131) begin
      { mem[4754:4754] } <= { data_i[34:34] };
    end 
    if(N11130) begin
      { mem[4753:4753] } <= { data_i[33:33] };
    end 
    if(N11129) begin
      { mem[4752:4752] } <= { data_i[32:32] };
    end 
    if(N11128) begin
      { mem[4751:4751] } <= { data_i[31:31] };
    end 
    if(N11127) begin
      { mem[4750:4750] } <= { data_i[30:30] };
    end 
    if(N11126) begin
      { mem[4749:4749] } <= { data_i[29:29] };
    end 
    if(N11125) begin
      { mem[4748:4748] } <= { data_i[28:28] };
    end 
    if(N11124) begin
      { mem[4747:4747] } <= { data_i[27:27] };
    end 
    if(N11123) begin
      { mem[4746:4746] } <= { data_i[26:26] };
    end 
    if(N11122) begin
      { mem[4745:4745] } <= { data_i[25:25] };
    end 
    if(N11121) begin
      { mem[4744:4744] } <= { data_i[24:24] };
    end 
    if(N11120) begin
      { mem[4743:4743] } <= { data_i[23:23] };
    end 
    if(N11119) begin
      { mem[4742:4742] } <= { data_i[22:22] };
    end 
    if(N11118) begin
      { mem[4741:4741] } <= { data_i[21:21] };
    end 
    if(N11117) begin
      { mem[4740:4740] } <= { data_i[20:20] };
    end 
    if(N11116) begin
      { mem[4739:4739] } <= { data_i[19:19] };
    end 
    if(N11115) begin
      { mem[4738:4738] } <= { data_i[18:18] };
    end 
    if(N11114) begin
      { mem[4737:4737] } <= { data_i[17:17] };
    end 
    if(N11113) begin
      { mem[4736:4736] } <= { data_i[16:16] };
    end 
    if(N11112) begin
      { mem[4735:4735] } <= { data_i[15:15] };
    end 
    if(N11111) begin
      { mem[4734:4734] } <= { data_i[14:14] };
    end 
    if(N11110) begin
      { mem[4733:4733] } <= { data_i[13:13] };
    end 
    if(N11109) begin
      { mem[4732:4732] } <= { data_i[12:12] };
    end 
    if(N11108) begin
      { mem[4731:4731] } <= { data_i[11:11] };
    end 
    if(N11107) begin
      { mem[4730:4730] } <= { data_i[10:10] };
    end 
    if(N11106) begin
      { mem[4729:4729] } <= { data_i[9:9] };
    end 
    if(N11105) begin
      { mem[4728:4728] } <= { data_i[8:8] };
    end 
    if(N11104) begin
      { mem[4727:4727] } <= { data_i[7:7] };
    end 
    if(N11103) begin
      { mem[4726:4726] } <= { data_i[6:6] };
    end 
    if(N11102) begin
      { mem[4725:4725] } <= { data_i[5:5] };
    end 
    if(N11101) begin
      { mem[4724:4724] } <= { data_i[4:4] };
    end 
    if(N11100) begin
      { mem[4723:4723] } <= { data_i[3:3] };
    end 
    if(N11099) begin
      { mem[4722:4722] } <= { data_i[2:2] };
    end 
    if(N11098) begin
      { mem[4721:4721] } <= { data_i[1:1] };
    end 
    if(N11097) begin
      { mem[4720:4720] } <= { data_i[0:0] };
    end 
    if(N11096) begin
      { mem[4719:4719] } <= { data_i[79:79] };
    end 
    if(N11095) begin
      { mem[4718:4718] } <= { data_i[78:78] };
    end 
    if(N11094) begin
      { mem[4717:4717] } <= { data_i[77:77] };
    end 
    if(N11093) begin
      { mem[4716:4716] } <= { data_i[76:76] };
    end 
    if(N11092) begin
      { mem[4715:4715] } <= { data_i[75:75] };
    end 
    if(N11091) begin
      { mem[4714:4714] } <= { data_i[74:74] };
    end 
    if(N11090) begin
      { mem[4713:4713] } <= { data_i[73:73] };
    end 
    if(N11089) begin
      { mem[4712:4712] } <= { data_i[72:72] };
    end 
    if(N11088) begin
      { mem[4711:4711] } <= { data_i[71:71] };
    end 
    if(N11087) begin
      { mem[4710:4710] } <= { data_i[70:70] };
    end 
    if(N11086) begin
      { mem[4709:4709] } <= { data_i[69:69] };
    end 
    if(N11085) begin
      { mem[4708:4708] } <= { data_i[68:68] };
    end 
    if(N11084) begin
      { mem[4707:4707] } <= { data_i[67:67] };
    end 
    if(N11083) begin
      { mem[4706:4706] } <= { data_i[66:66] };
    end 
    if(N11082) begin
      { mem[4705:4705] } <= { data_i[65:65] };
    end 
    if(N11081) begin
      { mem[4704:4704] } <= { data_i[64:64] };
    end 
    if(N11080) begin
      { mem[4703:4703] } <= { data_i[63:63] };
    end 
    if(N11079) begin
      { mem[4702:4702] } <= { data_i[62:62] };
    end 
    if(N11078) begin
      { mem[4701:4701] } <= { data_i[61:61] };
    end 
    if(N11077) begin
      { mem[4700:4700] } <= { data_i[60:60] };
    end 
    if(N11076) begin
      { mem[4699:4699] } <= { data_i[59:59] };
    end 
    if(N11075) begin
      { mem[4698:4698] } <= { data_i[58:58] };
    end 
    if(N11074) begin
      { mem[4697:4697] } <= { data_i[57:57] };
    end 
    if(N11073) begin
      { mem[4696:4696] } <= { data_i[56:56] };
    end 
    if(N11072) begin
      { mem[4695:4695] } <= { data_i[55:55] };
    end 
    if(N11071) begin
      { mem[4694:4694] } <= { data_i[54:54] };
    end 
    if(N11070) begin
      { mem[4693:4693] } <= { data_i[53:53] };
    end 
    if(N11069) begin
      { mem[4692:4692] } <= { data_i[52:52] };
    end 
    if(N11068) begin
      { mem[4691:4691] } <= { data_i[51:51] };
    end 
    if(N11067) begin
      { mem[4690:4690] } <= { data_i[50:50] };
    end 
    if(N11066) begin
      { mem[4689:4689] } <= { data_i[49:49] };
    end 
    if(N11065) begin
      { mem[4688:4688] } <= { data_i[48:48] };
    end 
    if(N11064) begin
      { mem[4687:4687] } <= { data_i[47:47] };
    end 
    if(N11063) begin
      { mem[4686:4686] } <= { data_i[46:46] };
    end 
    if(N11062) begin
      { mem[4685:4685] } <= { data_i[45:45] };
    end 
    if(N11061) begin
      { mem[4684:4684] } <= { data_i[44:44] };
    end 
    if(N11060) begin
      { mem[4683:4683] } <= { data_i[43:43] };
    end 
    if(N11059) begin
      { mem[4682:4682] } <= { data_i[42:42] };
    end 
    if(N11058) begin
      { mem[4681:4681] } <= { data_i[41:41] };
    end 
    if(N11057) begin
      { mem[4680:4680] } <= { data_i[40:40] };
    end 
    if(N11056) begin
      { mem[4679:4679] } <= { data_i[39:39] };
    end 
    if(N11055) begin
      { mem[4678:4678] } <= { data_i[38:38] };
    end 
    if(N11054) begin
      { mem[4677:4677] } <= { data_i[37:37] };
    end 
    if(N11053) begin
      { mem[4676:4676] } <= { data_i[36:36] };
    end 
    if(N11052) begin
      { mem[4675:4675] } <= { data_i[35:35] };
    end 
    if(N11051) begin
      { mem[4674:4674] } <= { data_i[34:34] };
    end 
    if(N11050) begin
      { mem[4673:4673] } <= { data_i[33:33] };
    end 
    if(N11049) begin
      { mem[4672:4672] } <= { data_i[32:32] };
    end 
    if(N11048) begin
      { mem[4671:4671] } <= { data_i[31:31] };
    end 
    if(N11047) begin
      { mem[4670:4670] } <= { data_i[30:30] };
    end 
    if(N11046) begin
      { mem[4669:4669] } <= { data_i[29:29] };
    end 
    if(N11045) begin
      { mem[4668:4668] } <= { data_i[28:28] };
    end 
    if(N11044) begin
      { mem[4667:4667] } <= { data_i[27:27] };
    end 
    if(N11043) begin
      { mem[4666:4666] } <= { data_i[26:26] };
    end 
    if(N11042) begin
      { mem[4665:4665] } <= { data_i[25:25] };
    end 
    if(N11041) begin
      { mem[4664:4664] } <= { data_i[24:24] };
    end 
    if(N11040) begin
      { mem[4663:4663] } <= { data_i[23:23] };
    end 
    if(N11039) begin
      { mem[4662:4662] } <= { data_i[22:22] };
    end 
    if(N11038) begin
      { mem[4661:4661] } <= { data_i[21:21] };
    end 
    if(N11037) begin
      { mem[4660:4660] } <= { data_i[20:20] };
    end 
    if(N11036) begin
      { mem[4659:4659] } <= { data_i[19:19] };
    end 
    if(N11035) begin
      { mem[4658:4658] } <= { data_i[18:18] };
    end 
    if(N11034) begin
      { mem[4657:4657] } <= { data_i[17:17] };
    end 
    if(N11033) begin
      { mem[4656:4656] } <= { data_i[16:16] };
    end 
    if(N11032) begin
      { mem[4655:4655] } <= { data_i[15:15] };
    end 
    if(N11031) begin
      { mem[4654:4654] } <= { data_i[14:14] };
    end 
    if(N11030) begin
      { mem[4653:4653] } <= { data_i[13:13] };
    end 
    if(N11029) begin
      { mem[4652:4652] } <= { data_i[12:12] };
    end 
    if(N11028) begin
      { mem[4651:4651] } <= { data_i[11:11] };
    end 
    if(N11027) begin
      { mem[4650:4650] } <= { data_i[10:10] };
    end 
    if(N11026) begin
      { mem[4649:4649] } <= { data_i[9:9] };
    end 
    if(N11025) begin
      { mem[4648:4648] } <= { data_i[8:8] };
    end 
    if(N11024) begin
      { mem[4647:4647] } <= { data_i[7:7] };
    end 
    if(N11023) begin
      { mem[4646:4646] } <= { data_i[6:6] };
    end 
    if(N11022) begin
      { mem[4645:4645] } <= { data_i[5:5] };
    end 
    if(N11021) begin
      { mem[4644:4644] } <= { data_i[4:4] };
    end 
    if(N11020) begin
      { mem[4643:4643] } <= { data_i[3:3] };
    end 
    if(N11019) begin
      { mem[4642:4642] } <= { data_i[2:2] };
    end 
    if(N11018) begin
      { mem[4641:4641] } <= { data_i[1:1] };
    end 
    if(N11017) begin
      { mem[4640:4640] } <= { data_i[0:0] };
    end 
    if(N11016) begin
      { mem[4639:4639] } <= { data_i[79:79] };
    end 
    if(N11015) begin
      { mem[4638:4638] } <= { data_i[78:78] };
    end 
    if(N11014) begin
      { mem[4637:4637] } <= { data_i[77:77] };
    end 
    if(N11013) begin
      { mem[4636:4636] } <= { data_i[76:76] };
    end 
    if(N11012) begin
      { mem[4635:4635] } <= { data_i[75:75] };
    end 
    if(N11011) begin
      { mem[4634:4634] } <= { data_i[74:74] };
    end 
    if(N11010) begin
      { mem[4633:4633] } <= { data_i[73:73] };
    end 
    if(N11009) begin
      { mem[4632:4632] } <= { data_i[72:72] };
    end 
    if(N11008) begin
      { mem[4631:4631] } <= { data_i[71:71] };
    end 
    if(N11007) begin
      { mem[4630:4630] } <= { data_i[70:70] };
    end 
    if(N11006) begin
      { mem[4629:4629] } <= { data_i[69:69] };
    end 
    if(N11005) begin
      { mem[4628:4628] } <= { data_i[68:68] };
    end 
    if(N11004) begin
      { mem[4627:4627] } <= { data_i[67:67] };
    end 
    if(N11003) begin
      { mem[4626:4626] } <= { data_i[66:66] };
    end 
    if(N11002) begin
      { mem[4625:4625] } <= { data_i[65:65] };
    end 
    if(N11001) begin
      { mem[4624:4624] } <= { data_i[64:64] };
    end 
    if(N11000) begin
      { mem[4623:4623] } <= { data_i[63:63] };
    end 
    if(N10999) begin
      { mem[4622:4622] } <= { data_i[62:62] };
    end 
    if(N10998) begin
      { mem[4621:4621] } <= { data_i[61:61] };
    end 
    if(N10997) begin
      { mem[4620:4620] } <= { data_i[60:60] };
    end 
    if(N10996) begin
      { mem[4619:4619] } <= { data_i[59:59] };
    end 
    if(N10995) begin
      { mem[4618:4618] } <= { data_i[58:58] };
    end 
    if(N10994) begin
      { mem[4617:4617] } <= { data_i[57:57] };
    end 
    if(N10993) begin
      { mem[4616:4616] } <= { data_i[56:56] };
    end 
    if(N10992) begin
      { mem[4615:4615] } <= { data_i[55:55] };
    end 
    if(N10991) begin
      { mem[4614:4614] } <= { data_i[54:54] };
    end 
    if(N10990) begin
      { mem[4613:4613] } <= { data_i[53:53] };
    end 
    if(N10989) begin
      { mem[4612:4612] } <= { data_i[52:52] };
    end 
    if(N10988) begin
      { mem[4611:4611] } <= { data_i[51:51] };
    end 
    if(N10987) begin
      { mem[4610:4610] } <= { data_i[50:50] };
    end 
    if(N10986) begin
      { mem[4609:4609] } <= { data_i[49:49] };
    end 
    if(N10985) begin
      { mem[4608:4608] } <= { data_i[48:48] };
    end 
    if(N10984) begin
      { mem[4607:4607] } <= { data_i[47:47] };
    end 
    if(N10983) begin
      { mem[4606:4606] } <= { data_i[46:46] };
    end 
    if(N10982) begin
      { mem[4605:4605] } <= { data_i[45:45] };
    end 
    if(N10981) begin
      { mem[4604:4604] } <= { data_i[44:44] };
    end 
    if(N10980) begin
      { mem[4603:4603] } <= { data_i[43:43] };
    end 
    if(N10979) begin
      { mem[4602:4602] } <= { data_i[42:42] };
    end 
    if(N10978) begin
      { mem[4601:4601] } <= { data_i[41:41] };
    end 
    if(N10977) begin
      { mem[4600:4600] } <= { data_i[40:40] };
    end 
    if(N10976) begin
      { mem[4599:4599] } <= { data_i[39:39] };
    end 
    if(N10975) begin
      { mem[4598:4598] } <= { data_i[38:38] };
    end 
    if(N10974) begin
      { mem[4597:4597] } <= { data_i[37:37] };
    end 
    if(N10973) begin
      { mem[4596:4596] } <= { data_i[36:36] };
    end 
    if(N10972) begin
      { mem[4595:4595] } <= { data_i[35:35] };
    end 
    if(N10971) begin
      { mem[4594:4594] } <= { data_i[34:34] };
    end 
    if(N10970) begin
      { mem[4593:4593] } <= { data_i[33:33] };
    end 
    if(N10969) begin
      { mem[4592:4592] } <= { data_i[32:32] };
    end 
    if(N10968) begin
      { mem[4591:4591] } <= { data_i[31:31] };
    end 
    if(N10967) begin
      { mem[4590:4590] } <= { data_i[30:30] };
    end 
    if(N10966) begin
      { mem[4589:4589] } <= { data_i[29:29] };
    end 
    if(N10965) begin
      { mem[4588:4588] } <= { data_i[28:28] };
    end 
    if(N10964) begin
      { mem[4587:4587] } <= { data_i[27:27] };
    end 
    if(N10963) begin
      { mem[4586:4586] } <= { data_i[26:26] };
    end 
    if(N10962) begin
      { mem[4585:4585] } <= { data_i[25:25] };
    end 
    if(N10961) begin
      { mem[4584:4584] } <= { data_i[24:24] };
    end 
    if(N10960) begin
      { mem[4583:4583] } <= { data_i[23:23] };
    end 
    if(N10959) begin
      { mem[4582:4582] } <= { data_i[22:22] };
    end 
    if(N10958) begin
      { mem[4581:4581] } <= { data_i[21:21] };
    end 
    if(N10957) begin
      { mem[4580:4580] } <= { data_i[20:20] };
    end 
    if(N10956) begin
      { mem[4579:4579] } <= { data_i[19:19] };
    end 
    if(N10955) begin
      { mem[4578:4578] } <= { data_i[18:18] };
    end 
    if(N10954) begin
      { mem[4577:4577] } <= { data_i[17:17] };
    end 
    if(N10953) begin
      { mem[4576:4576] } <= { data_i[16:16] };
    end 
    if(N10952) begin
      { mem[4575:4575] } <= { data_i[15:15] };
    end 
    if(N10951) begin
      { mem[4574:4574] } <= { data_i[14:14] };
    end 
    if(N10950) begin
      { mem[4573:4573] } <= { data_i[13:13] };
    end 
    if(N10949) begin
      { mem[4572:4572] } <= { data_i[12:12] };
    end 
    if(N10948) begin
      { mem[4571:4571] } <= { data_i[11:11] };
    end 
    if(N10947) begin
      { mem[4570:4570] } <= { data_i[10:10] };
    end 
    if(N10946) begin
      { mem[4569:4569] } <= { data_i[9:9] };
    end 
    if(N10945) begin
      { mem[4568:4568] } <= { data_i[8:8] };
    end 
    if(N10944) begin
      { mem[4567:4567] } <= { data_i[7:7] };
    end 
    if(N10943) begin
      { mem[4566:4566] } <= { data_i[6:6] };
    end 
    if(N10942) begin
      { mem[4565:4565] } <= { data_i[5:5] };
    end 
    if(N10941) begin
      { mem[4564:4564] } <= { data_i[4:4] };
    end 
    if(N10940) begin
      { mem[4563:4563] } <= { data_i[3:3] };
    end 
    if(N10939) begin
      { mem[4562:4562] } <= { data_i[2:2] };
    end 
    if(N10938) begin
      { mem[4561:4561] } <= { data_i[1:1] };
    end 
    if(N10937) begin
      { mem[4560:4560] } <= { data_i[0:0] };
    end 
    if(N10936) begin
      { mem[4559:4559] } <= { data_i[79:79] };
    end 
    if(N10935) begin
      { mem[4558:4558] } <= { data_i[78:78] };
    end 
    if(N10934) begin
      { mem[4557:4557] } <= { data_i[77:77] };
    end 
    if(N10933) begin
      { mem[4556:4556] } <= { data_i[76:76] };
    end 
    if(N10932) begin
      { mem[4555:4555] } <= { data_i[75:75] };
    end 
    if(N10931) begin
      { mem[4554:4554] } <= { data_i[74:74] };
    end 
    if(N10930) begin
      { mem[4553:4553] } <= { data_i[73:73] };
    end 
    if(N10929) begin
      { mem[4552:4552] } <= { data_i[72:72] };
    end 
    if(N10928) begin
      { mem[4551:4551] } <= { data_i[71:71] };
    end 
    if(N10927) begin
      { mem[4550:4550] } <= { data_i[70:70] };
    end 
    if(N10926) begin
      { mem[4549:4549] } <= { data_i[69:69] };
    end 
    if(N10925) begin
      { mem[4548:4548] } <= { data_i[68:68] };
    end 
    if(N10924) begin
      { mem[4547:4547] } <= { data_i[67:67] };
    end 
    if(N10923) begin
      { mem[4546:4546] } <= { data_i[66:66] };
    end 
    if(N10922) begin
      { mem[4545:4545] } <= { data_i[65:65] };
    end 
    if(N10921) begin
      { mem[4544:4544] } <= { data_i[64:64] };
    end 
    if(N10920) begin
      { mem[4543:4543] } <= { data_i[63:63] };
    end 
    if(N10919) begin
      { mem[4542:4542] } <= { data_i[62:62] };
    end 
    if(N10918) begin
      { mem[4541:4541] } <= { data_i[61:61] };
    end 
    if(N10917) begin
      { mem[4540:4540] } <= { data_i[60:60] };
    end 
    if(N10916) begin
      { mem[4539:4539] } <= { data_i[59:59] };
    end 
    if(N10915) begin
      { mem[4538:4538] } <= { data_i[58:58] };
    end 
    if(N10914) begin
      { mem[4537:4537] } <= { data_i[57:57] };
    end 
    if(N10913) begin
      { mem[4536:4536] } <= { data_i[56:56] };
    end 
    if(N10912) begin
      { mem[4535:4535] } <= { data_i[55:55] };
    end 
    if(N10911) begin
      { mem[4534:4534] } <= { data_i[54:54] };
    end 
    if(N10910) begin
      { mem[4533:4533] } <= { data_i[53:53] };
    end 
    if(N10909) begin
      { mem[4532:4532] } <= { data_i[52:52] };
    end 
    if(N10908) begin
      { mem[4531:4531] } <= { data_i[51:51] };
    end 
    if(N10907) begin
      { mem[4530:4530] } <= { data_i[50:50] };
    end 
    if(N10906) begin
      { mem[4529:4529] } <= { data_i[49:49] };
    end 
    if(N10905) begin
      { mem[4528:4528] } <= { data_i[48:48] };
    end 
    if(N10904) begin
      { mem[4527:4527] } <= { data_i[47:47] };
    end 
    if(N10903) begin
      { mem[4526:4526] } <= { data_i[46:46] };
    end 
    if(N10902) begin
      { mem[4525:4525] } <= { data_i[45:45] };
    end 
    if(N10901) begin
      { mem[4524:4524] } <= { data_i[44:44] };
    end 
    if(N10900) begin
      { mem[4523:4523] } <= { data_i[43:43] };
    end 
    if(N10899) begin
      { mem[4522:4522] } <= { data_i[42:42] };
    end 
    if(N10898) begin
      { mem[4521:4521] } <= { data_i[41:41] };
    end 
    if(N10897) begin
      { mem[4520:4520] } <= { data_i[40:40] };
    end 
    if(N10896) begin
      { mem[4519:4519] } <= { data_i[39:39] };
    end 
    if(N10895) begin
      { mem[4518:4518] } <= { data_i[38:38] };
    end 
    if(N10894) begin
      { mem[4517:4517] } <= { data_i[37:37] };
    end 
    if(N10893) begin
      { mem[4516:4516] } <= { data_i[36:36] };
    end 
    if(N10892) begin
      { mem[4515:4515] } <= { data_i[35:35] };
    end 
    if(N10891) begin
      { mem[4514:4514] } <= { data_i[34:34] };
    end 
    if(N10890) begin
      { mem[4513:4513] } <= { data_i[33:33] };
    end 
    if(N10889) begin
      { mem[4512:4512] } <= { data_i[32:32] };
    end 
    if(N10888) begin
      { mem[4511:4511] } <= { data_i[31:31] };
    end 
    if(N10887) begin
      { mem[4510:4510] } <= { data_i[30:30] };
    end 
    if(N10886) begin
      { mem[4509:4509] } <= { data_i[29:29] };
    end 
    if(N10885) begin
      { mem[4508:4508] } <= { data_i[28:28] };
    end 
    if(N10884) begin
      { mem[4507:4507] } <= { data_i[27:27] };
    end 
    if(N10883) begin
      { mem[4506:4506] } <= { data_i[26:26] };
    end 
    if(N10882) begin
      { mem[4505:4505] } <= { data_i[25:25] };
    end 
    if(N10881) begin
      { mem[4504:4504] } <= { data_i[24:24] };
    end 
    if(N10880) begin
      { mem[4503:4503] } <= { data_i[23:23] };
    end 
    if(N10879) begin
      { mem[4502:4502] } <= { data_i[22:22] };
    end 
    if(N10878) begin
      { mem[4501:4501] } <= { data_i[21:21] };
    end 
    if(N10877) begin
      { mem[4500:4500] } <= { data_i[20:20] };
    end 
    if(N10876) begin
      { mem[4499:4499] } <= { data_i[19:19] };
    end 
    if(N10875) begin
      { mem[4498:4498] } <= { data_i[18:18] };
    end 
    if(N10874) begin
      { mem[4497:4497] } <= { data_i[17:17] };
    end 
    if(N10873) begin
      { mem[4496:4496] } <= { data_i[16:16] };
    end 
    if(N10872) begin
      { mem[4495:4495] } <= { data_i[15:15] };
    end 
    if(N10871) begin
      { mem[4494:4494] } <= { data_i[14:14] };
    end 
    if(N10870) begin
      { mem[4493:4493] } <= { data_i[13:13] };
    end 
    if(N10869) begin
      { mem[4492:4492] } <= { data_i[12:12] };
    end 
    if(N10868) begin
      { mem[4491:4491] } <= { data_i[11:11] };
    end 
    if(N10867) begin
      { mem[4490:4490] } <= { data_i[10:10] };
    end 
    if(N10866) begin
      { mem[4489:4489] } <= { data_i[9:9] };
    end 
    if(N10865) begin
      { mem[4488:4488] } <= { data_i[8:8] };
    end 
    if(N10864) begin
      { mem[4487:4487] } <= { data_i[7:7] };
    end 
    if(N10863) begin
      { mem[4486:4486] } <= { data_i[6:6] };
    end 
    if(N10862) begin
      { mem[4485:4485] } <= { data_i[5:5] };
    end 
    if(N10861) begin
      { mem[4484:4484] } <= { data_i[4:4] };
    end 
    if(N10860) begin
      { mem[4483:4483] } <= { data_i[3:3] };
    end 
    if(N10859) begin
      { mem[4482:4482] } <= { data_i[2:2] };
    end 
    if(N10858) begin
      { mem[4481:4481] } <= { data_i[1:1] };
    end 
    if(N10857) begin
      { mem[4480:4480] } <= { data_i[0:0] };
    end 
    if(N10856) begin
      { mem[4479:4479] } <= { data_i[79:79] };
    end 
    if(N10855) begin
      { mem[4478:4478] } <= { data_i[78:78] };
    end 
    if(N10854) begin
      { mem[4477:4477] } <= { data_i[77:77] };
    end 
    if(N10853) begin
      { mem[4476:4476] } <= { data_i[76:76] };
    end 
    if(N10852) begin
      { mem[4475:4475] } <= { data_i[75:75] };
    end 
    if(N10851) begin
      { mem[4474:4474] } <= { data_i[74:74] };
    end 
    if(N10850) begin
      { mem[4473:4473] } <= { data_i[73:73] };
    end 
    if(N10849) begin
      { mem[4472:4472] } <= { data_i[72:72] };
    end 
    if(N10848) begin
      { mem[4471:4471] } <= { data_i[71:71] };
    end 
    if(N10847) begin
      { mem[4470:4470] } <= { data_i[70:70] };
    end 
    if(N10846) begin
      { mem[4469:4469] } <= { data_i[69:69] };
    end 
    if(N10845) begin
      { mem[4468:4468] } <= { data_i[68:68] };
    end 
    if(N10844) begin
      { mem[4467:4467] } <= { data_i[67:67] };
    end 
    if(N10843) begin
      { mem[4466:4466] } <= { data_i[66:66] };
    end 
    if(N10842) begin
      { mem[4465:4465] } <= { data_i[65:65] };
    end 
    if(N10841) begin
      { mem[4464:4464] } <= { data_i[64:64] };
    end 
    if(N10840) begin
      { mem[4463:4463] } <= { data_i[63:63] };
    end 
    if(N10839) begin
      { mem[4462:4462] } <= { data_i[62:62] };
    end 
    if(N10838) begin
      { mem[4461:4461] } <= { data_i[61:61] };
    end 
    if(N10837) begin
      { mem[4460:4460] } <= { data_i[60:60] };
    end 
    if(N10836) begin
      { mem[4459:4459] } <= { data_i[59:59] };
    end 
    if(N10835) begin
      { mem[4458:4458] } <= { data_i[58:58] };
    end 
    if(N10834) begin
      { mem[4457:4457] } <= { data_i[57:57] };
    end 
    if(N10833) begin
      { mem[4456:4456] } <= { data_i[56:56] };
    end 
    if(N10832) begin
      { mem[4455:4455] } <= { data_i[55:55] };
    end 
    if(N10831) begin
      { mem[4454:4454] } <= { data_i[54:54] };
    end 
    if(N10830) begin
      { mem[4453:4453] } <= { data_i[53:53] };
    end 
    if(N10829) begin
      { mem[4452:4452] } <= { data_i[52:52] };
    end 
    if(N10828) begin
      { mem[4451:4451] } <= { data_i[51:51] };
    end 
    if(N10827) begin
      { mem[4450:4450] } <= { data_i[50:50] };
    end 
    if(N10826) begin
      { mem[4449:4449] } <= { data_i[49:49] };
    end 
    if(N10825) begin
      { mem[4448:4448] } <= { data_i[48:48] };
    end 
    if(N10824) begin
      { mem[4447:4447] } <= { data_i[47:47] };
    end 
    if(N10823) begin
      { mem[4446:4446] } <= { data_i[46:46] };
    end 
    if(N10822) begin
      { mem[4445:4445] } <= { data_i[45:45] };
    end 
    if(N10821) begin
      { mem[4444:4444] } <= { data_i[44:44] };
    end 
    if(N10820) begin
      { mem[4443:4443] } <= { data_i[43:43] };
    end 
    if(N10819) begin
      { mem[4442:4442] } <= { data_i[42:42] };
    end 
    if(N10818) begin
      { mem[4441:4441] } <= { data_i[41:41] };
    end 
    if(N10817) begin
      { mem[4440:4440] } <= { data_i[40:40] };
    end 
    if(N10816) begin
      { mem[4439:4439] } <= { data_i[39:39] };
    end 
    if(N10815) begin
      { mem[4438:4438] } <= { data_i[38:38] };
    end 
    if(N10814) begin
      { mem[4437:4437] } <= { data_i[37:37] };
    end 
    if(N10813) begin
      { mem[4436:4436] } <= { data_i[36:36] };
    end 
    if(N10812) begin
      { mem[4435:4435] } <= { data_i[35:35] };
    end 
    if(N10811) begin
      { mem[4434:4434] } <= { data_i[34:34] };
    end 
    if(N10810) begin
      { mem[4433:4433] } <= { data_i[33:33] };
    end 
    if(N10809) begin
      { mem[4432:4432] } <= { data_i[32:32] };
    end 
    if(N10808) begin
      { mem[4431:4431] } <= { data_i[31:31] };
    end 
    if(N10807) begin
      { mem[4430:4430] } <= { data_i[30:30] };
    end 
    if(N10806) begin
      { mem[4429:4429] } <= { data_i[29:29] };
    end 
    if(N10805) begin
      { mem[4428:4428] } <= { data_i[28:28] };
    end 
    if(N10804) begin
      { mem[4427:4427] } <= { data_i[27:27] };
    end 
    if(N10803) begin
      { mem[4426:4426] } <= { data_i[26:26] };
    end 
    if(N10802) begin
      { mem[4425:4425] } <= { data_i[25:25] };
    end 
    if(N10801) begin
      { mem[4424:4424] } <= { data_i[24:24] };
    end 
    if(N10800) begin
      { mem[4423:4423] } <= { data_i[23:23] };
    end 
    if(N10799) begin
      { mem[4422:4422] } <= { data_i[22:22] };
    end 
    if(N10798) begin
      { mem[4421:4421] } <= { data_i[21:21] };
    end 
    if(N10797) begin
      { mem[4420:4420] } <= { data_i[20:20] };
    end 
    if(N10796) begin
      { mem[4419:4419] } <= { data_i[19:19] };
    end 
    if(N10795) begin
      { mem[4418:4418] } <= { data_i[18:18] };
    end 
    if(N10794) begin
      { mem[4417:4417] } <= { data_i[17:17] };
    end 
    if(N10793) begin
      { mem[4416:4416] } <= { data_i[16:16] };
    end 
    if(N10792) begin
      { mem[4415:4415] } <= { data_i[15:15] };
    end 
    if(N10791) begin
      { mem[4414:4414] } <= { data_i[14:14] };
    end 
    if(N10790) begin
      { mem[4413:4413] } <= { data_i[13:13] };
    end 
    if(N10789) begin
      { mem[4412:4412] } <= { data_i[12:12] };
    end 
    if(N10788) begin
      { mem[4411:4411] } <= { data_i[11:11] };
    end 
    if(N10787) begin
      { mem[4410:4410] } <= { data_i[10:10] };
    end 
    if(N10786) begin
      { mem[4409:4409] } <= { data_i[9:9] };
    end 
    if(N10785) begin
      { mem[4408:4408] } <= { data_i[8:8] };
    end 
    if(N10784) begin
      { mem[4407:4407] } <= { data_i[7:7] };
    end 
    if(N10783) begin
      { mem[4406:4406] } <= { data_i[6:6] };
    end 
    if(N10782) begin
      { mem[4405:4405] } <= { data_i[5:5] };
    end 
    if(N10781) begin
      { mem[4404:4404] } <= { data_i[4:4] };
    end 
    if(N10780) begin
      { mem[4403:4403] } <= { data_i[3:3] };
    end 
    if(N10779) begin
      { mem[4402:4402] } <= { data_i[2:2] };
    end 
    if(N10778) begin
      { mem[4401:4401] } <= { data_i[1:1] };
    end 
    if(N10777) begin
      { mem[4400:4400] } <= { data_i[0:0] };
    end 
    if(N10776) begin
      { mem[4399:4399] } <= { data_i[79:79] };
    end 
    if(N10775) begin
      { mem[4398:4398] } <= { data_i[78:78] };
    end 
    if(N10774) begin
      { mem[4397:4397] } <= { data_i[77:77] };
    end 
    if(N10773) begin
      { mem[4396:4396] } <= { data_i[76:76] };
    end 
    if(N10772) begin
      { mem[4395:4395] } <= { data_i[75:75] };
    end 
    if(N10771) begin
      { mem[4394:4394] } <= { data_i[74:74] };
    end 
    if(N10770) begin
      { mem[4393:4393] } <= { data_i[73:73] };
    end 
    if(N10769) begin
      { mem[4392:4392] } <= { data_i[72:72] };
    end 
    if(N10768) begin
      { mem[4391:4391] } <= { data_i[71:71] };
    end 
    if(N10767) begin
      { mem[4390:4390] } <= { data_i[70:70] };
    end 
    if(N10766) begin
      { mem[4389:4389] } <= { data_i[69:69] };
    end 
    if(N10765) begin
      { mem[4388:4388] } <= { data_i[68:68] };
    end 
    if(N10764) begin
      { mem[4387:4387] } <= { data_i[67:67] };
    end 
    if(N10763) begin
      { mem[4386:4386] } <= { data_i[66:66] };
    end 
    if(N10762) begin
      { mem[4385:4385] } <= { data_i[65:65] };
    end 
    if(N10761) begin
      { mem[4384:4384] } <= { data_i[64:64] };
    end 
    if(N10760) begin
      { mem[4383:4383] } <= { data_i[63:63] };
    end 
    if(N10759) begin
      { mem[4382:4382] } <= { data_i[62:62] };
    end 
    if(N10758) begin
      { mem[4381:4381] } <= { data_i[61:61] };
    end 
    if(N10757) begin
      { mem[4380:4380] } <= { data_i[60:60] };
    end 
    if(N10756) begin
      { mem[4379:4379] } <= { data_i[59:59] };
    end 
    if(N10755) begin
      { mem[4378:4378] } <= { data_i[58:58] };
    end 
    if(N10754) begin
      { mem[4377:4377] } <= { data_i[57:57] };
    end 
    if(N10753) begin
      { mem[4376:4376] } <= { data_i[56:56] };
    end 
    if(N10752) begin
      { mem[4375:4375] } <= { data_i[55:55] };
    end 
    if(N10751) begin
      { mem[4374:4374] } <= { data_i[54:54] };
    end 
    if(N10750) begin
      { mem[4373:4373] } <= { data_i[53:53] };
    end 
    if(N10749) begin
      { mem[4372:4372] } <= { data_i[52:52] };
    end 
    if(N10748) begin
      { mem[4371:4371] } <= { data_i[51:51] };
    end 
    if(N10747) begin
      { mem[4370:4370] } <= { data_i[50:50] };
    end 
    if(N10746) begin
      { mem[4369:4369] } <= { data_i[49:49] };
    end 
    if(N10745) begin
      { mem[4368:4368] } <= { data_i[48:48] };
    end 
    if(N10744) begin
      { mem[4367:4367] } <= { data_i[47:47] };
    end 
    if(N10743) begin
      { mem[4366:4366] } <= { data_i[46:46] };
    end 
    if(N10742) begin
      { mem[4365:4365] } <= { data_i[45:45] };
    end 
    if(N10741) begin
      { mem[4364:4364] } <= { data_i[44:44] };
    end 
    if(N10740) begin
      { mem[4363:4363] } <= { data_i[43:43] };
    end 
    if(N10739) begin
      { mem[4362:4362] } <= { data_i[42:42] };
    end 
    if(N10738) begin
      { mem[4361:4361] } <= { data_i[41:41] };
    end 
    if(N10737) begin
      { mem[4360:4360] } <= { data_i[40:40] };
    end 
    if(N10736) begin
      { mem[4359:4359] } <= { data_i[39:39] };
    end 
    if(N10735) begin
      { mem[4358:4358] } <= { data_i[38:38] };
    end 
    if(N10734) begin
      { mem[4357:4357] } <= { data_i[37:37] };
    end 
    if(N10733) begin
      { mem[4356:4356] } <= { data_i[36:36] };
    end 
    if(N10732) begin
      { mem[4355:4355] } <= { data_i[35:35] };
    end 
    if(N10731) begin
      { mem[4354:4354] } <= { data_i[34:34] };
    end 
    if(N10730) begin
      { mem[4353:4353] } <= { data_i[33:33] };
    end 
    if(N10729) begin
      { mem[4352:4352] } <= { data_i[32:32] };
    end 
    if(N10728) begin
      { mem[4351:4351] } <= { data_i[31:31] };
    end 
    if(N10727) begin
      { mem[4350:4350] } <= { data_i[30:30] };
    end 
    if(N10726) begin
      { mem[4349:4349] } <= { data_i[29:29] };
    end 
    if(N10725) begin
      { mem[4348:4348] } <= { data_i[28:28] };
    end 
    if(N10724) begin
      { mem[4347:4347] } <= { data_i[27:27] };
    end 
    if(N10723) begin
      { mem[4346:4346] } <= { data_i[26:26] };
    end 
    if(N10722) begin
      { mem[4345:4345] } <= { data_i[25:25] };
    end 
    if(N10721) begin
      { mem[4344:4344] } <= { data_i[24:24] };
    end 
    if(N10720) begin
      { mem[4343:4343] } <= { data_i[23:23] };
    end 
    if(N10719) begin
      { mem[4342:4342] } <= { data_i[22:22] };
    end 
    if(N10718) begin
      { mem[4341:4341] } <= { data_i[21:21] };
    end 
    if(N10717) begin
      { mem[4340:4340] } <= { data_i[20:20] };
    end 
    if(N10716) begin
      { mem[4339:4339] } <= { data_i[19:19] };
    end 
    if(N10715) begin
      { mem[4338:4338] } <= { data_i[18:18] };
    end 
    if(N10714) begin
      { mem[4337:4337] } <= { data_i[17:17] };
    end 
    if(N10713) begin
      { mem[4336:4336] } <= { data_i[16:16] };
    end 
    if(N10712) begin
      { mem[4335:4335] } <= { data_i[15:15] };
    end 
    if(N10711) begin
      { mem[4334:4334] } <= { data_i[14:14] };
    end 
    if(N10710) begin
      { mem[4333:4333] } <= { data_i[13:13] };
    end 
    if(N10709) begin
      { mem[4332:4332] } <= { data_i[12:12] };
    end 
    if(N10708) begin
      { mem[4331:4331] } <= { data_i[11:11] };
    end 
    if(N10707) begin
      { mem[4330:4330] } <= { data_i[10:10] };
    end 
    if(N10706) begin
      { mem[4329:4329] } <= { data_i[9:9] };
    end 
    if(N10705) begin
      { mem[4328:4328] } <= { data_i[8:8] };
    end 
    if(N10704) begin
      { mem[4327:4327] } <= { data_i[7:7] };
    end 
    if(N10703) begin
      { mem[4326:4326] } <= { data_i[6:6] };
    end 
    if(N10702) begin
      { mem[4325:4325] } <= { data_i[5:5] };
    end 
    if(N10701) begin
      { mem[4324:4324] } <= { data_i[4:4] };
    end 
    if(N10700) begin
      { mem[4323:4323] } <= { data_i[3:3] };
    end 
    if(N10699) begin
      { mem[4322:4322] } <= { data_i[2:2] };
    end 
    if(N10698) begin
      { mem[4321:4321] } <= { data_i[1:1] };
    end 
    if(N10697) begin
      { mem[4320:4320] } <= { data_i[0:0] };
    end 
    if(N10696) begin
      { mem[4319:4319] } <= { data_i[79:79] };
    end 
    if(N10695) begin
      { mem[4318:4318] } <= { data_i[78:78] };
    end 
    if(N10694) begin
      { mem[4317:4317] } <= { data_i[77:77] };
    end 
    if(N10693) begin
      { mem[4316:4316] } <= { data_i[76:76] };
    end 
    if(N10692) begin
      { mem[4315:4315] } <= { data_i[75:75] };
    end 
    if(N10691) begin
      { mem[4314:4314] } <= { data_i[74:74] };
    end 
    if(N10690) begin
      { mem[4313:4313] } <= { data_i[73:73] };
    end 
    if(N10689) begin
      { mem[4312:4312] } <= { data_i[72:72] };
    end 
    if(N10688) begin
      { mem[4311:4311] } <= { data_i[71:71] };
    end 
    if(N10687) begin
      { mem[4310:4310] } <= { data_i[70:70] };
    end 
    if(N10686) begin
      { mem[4309:4309] } <= { data_i[69:69] };
    end 
    if(N10685) begin
      { mem[4308:4308] } <= { data_i[68:68] };
    end 
    if(N10684) begin
      { mem[4307:4307] } <= { data_i[67:67] };
    end 
    if(N10683) begin
      { mem[4306:4306] } <= { data_i[66:66] };
    end 
    if(N10682) begin
      { mem[4305:4305] } <= { data_i[65:65] };
    end 
    if(N10681) begin
      { mem[4304:4304] } <= { data_i[64:64] };
    end 
    if(N10680) begin
      { mem[4303:4303] } <= { data_i[63:63] };
    end 
    if(N10679) begin
      { mem[4302:4302] } <= { data_i[62:62] };
    end 
    if(N10678) begin
      { mem[4301:4301] } <= { data_i[61:61] };
    end 
    if(N10677) begin
      { mem[4300:4300] } <= { data_i[60:60] };
    end 
    if(N10676) begin
      { mem[4299:4299] } <= { data_i[59:59] };
    end 
    if(N10675) begin
      { mem[4298:4298] } <= { data_i[58:58] };
    end 
    if(N10674) begin
      { mem[4297:4297] } <= { data_i[57:57] };
    end 
    if(N10673) begin
      { mem[4296:4296] } <= { data_i[56:56] };
    end 
    if(N10672) begin
      { mem[4295:4295] } <= { data_i[55:55] };
    end 
    if(N10671) begin
      { mem[4294:4294] } <= { data_i[54:54] };
    end 
    if(N10670) begin
      { mem[4293:4293] } <= { data_i[53:53] };
    end 
    if(N10669) begin
      { mem[4292:4292] } <= { data_i[52:52] };
    end 
    if(N10668) begin
      { mem[4291:4291] } <= { data_i[51:51] };
    end 
    if(N10667) begin
      { mem[4290:4290] } <= { data_i[50:50] };
    end 
    if(N10666) begin
      { mem[4289:4289] } <= { data_i[49:49] };
    end 
    if(N10665) begin
      { mem[4288:4288] } <= { data_i[48:48] };
    end 
    if(N10664) begin
      { mem[4287:4287] } <= { data_i[47:47] };
    end 
    if(N10663) begin
      { mem[4286:4286] } <= { data_i[46:46] };
    end 
    if(N10662) begin
      { mem[4285:4285] } <= { data_i[45:45] };
    end 
    if(N10661) begin
      { mem[4284:4284] } <= { data_i[44:44] };
    end 
    if(N10660) begin
      { mem[4283:4283] } <= { data_i[43:43] };
    end 
    if(N10659) begin
      { mem[4282:4282] } <= { data_i[42:42] };
    end 
    if(N10658) begin
      { mem[4281:4281] } <= { data_i[41:41] };
    end 
    if(N10657) begin
      { mem[4280:4280] } <= { data_i[40:40] };
    end 
    if(N10656) begin
      { mem[4279:4279] } <= { data_i[39:39] };
    end 
    if(N10655) begin
      { mem[4278:4278] } <= { data_i[38:38] };
    end 
    if(N10654) begin
      { mem[4277:4277] } <= { data_i[37:37] };
    end 
    if(N10653) begin
      { mem[4276:4276] } <= { data_i[36:36] };
    end 
    if(N10652) begin
      { mem[4275:4275] } <= { data_i[35:35] };
    end 
    if(N10651) begin
      { mem[4274:4274] } <= { data_i[34:34] };
    end 
    if(N10650) begin
      { mem[4273:4273] } <= { data_i[33:33] };
    end 
    if(N10649) begin
      { mem[4272:4272] } <= { data_i[32:32] };
    end 
    if(N10648) begin
      { mem[4271:4271] } <= { data_i[31:31] };
    end 
    if(N10647) begin
      { mem[4270:4270] } <= { data_i[30:30] };
    end 
    if(N10646) begin
      { mem[4269:4269] } <= { data_i[29:29] };
    end 
    if(N10645) begin
      { mem[4268:4268] } <= { data_i[28:28] };
    end 
    if(N10644) begin
      { mem[4267:4267] } <= { data_i[27:27] };
    end 
    if(N10643) begin
      { mem[4266:4266] } <= { data_i[26:26] };
    end 
    if(N10642) begin
      { mem[4265:4265] } <= { data_i[25:25] };
    end 
    if(N10641) begin
      { mem[4264:4264] } <= { data_i[24:24] };
    end 
    if(N10640) begin
      { mem[4263:4263] } <= { data_i[23:23] };
    end 
    if(N10639) begin
      { mem[4262:4262] } <= { data_i[22:22] };
    end 
    if(N10638) begin
      { mem[4261:4261] } <= { data_i[21:21] };
    end 
    if(N10637) begin
      { mem[4260:4260] } <= { data_i[20:20] };
    end 
    if(N10636) begin
      { mem[4259:4259] } <= { data_i[19:19] };
    end 
    if(N10635) begin
      { mem[4258:4258] } <= { data_i[18:18] };
    end 
    if(N10634) begin
      { mem[4257:4257] } <= { data_i[17:17] };
    end 
    if(N10633) begin
      { mem[4256:4256] } <= { data_i[16:16] };
    end 
    if(N10632) begin
      { mem[4255:4255] } <= { data_i[15:15] };
    end 
    if(N10631) begin
      { mem[4254:4254] } <= { data_i[14:14] };
    end 
    if(N10630) begin
      { mem[4253:4253] } <= { data_i[13:13] };
    end 
    if(N10629) begin
      { mem[4252:4252] } <= { data_i[12:12] };
    end 
    if(N10628) begin
      { mem[4251:4251] } <= { data_i[11:11] };
    end 
    if(N10627) begin
      { mem[4250:4250] } <= { data_i[10:10] };
    end 
    if(N10626) begin
      { mem[4249:4249] } <= { data_i[9:9] };
    end 
    if(N10625) begin
      { mem[4248:4248] } <= { data_i[8:8] };
    end 
    if(N10624) begin
      { mem[4247:4247] } <= { data_i[7:7] };
    end 
    if(N10623) begin
      { mem[4246:4246] } <= { data_i[6:6] };
    end 
    if(N10622) begin
      { mem[4245:4245] } <= { data_i[5:5] };
    end 
    if(N10621) begin
      { mem[4244:4244] } <= { data_i[4:4] };
    end 
    if(N10620) begin
      { mem[4243:4243] } <= { data_i[3:3] };
    end 
    if(N10619) begin
      { mem[4242:4242] } <= { data_i[2:2] };
    end 
    if(N10618) begin
      { mem[4241:4241] } <= { data_i[1:1] };
    end 
    if(N10617) begin
      { mem[4240:4240] } <= { data_i[0:0] };
    end 
    if(N10616) begin
      { mem[4239:4239] } <= { data_i[79:79] };
    end 
    if(N10615) begin
      { mem[4238:4238] } <= { data_i[78:78] };
    end 
    if(N10614) begin
      { mem[4237:4237] } <= { data_i[77:77] };
    end 
    if(N10613) begin
      { mem[4236:4236] } <= { data_i[76:76] };
    end 
    if(N10612) begin
      { mem[4235:4235] } <= { data_i[75:75] };
    end 
    if(N10611) begin
      { mem[4234:4234] } <= { data_i[74:74] };
    end 
    if(N10610) begin
      { mem[4233:4233] } <= { data_i[73:73] };
    end 
    if(N10609) begin
      { mem[4232:4232] } <= { data_i[72:72] };
    end 
    if(N10608) begin
      { mem[4231:4231] } <= { data_i[71:71] };
    end 
    if(N10607) begin
      { mem[4230:4230] } <= { data_i[70:70] };
    end 
    if(N10606) begin
      { mem[4229:4229] } <= { data_i[69:69] };
    end 
    if(N10605) begin
      { mem[4228:4228] } <= { data_i[68:68] };
    end 
    if(N10604) begin
      { mem[4227:4227] } <= { data_i[67:67] };
    end 
    if(N10603) begin
      { mem[4226:4226] } <= { data_i[66:66] };
    end 
    if(N10602) begin
      { mem[4225:4225] } <= { data_i[65:65] };
    end 
    if(N10601) begin
      { mem[4224:4224] } <= { data_i[64:64] };
    end 
    if(N10600) begin
      { mem[4223:4223] } <= { data_i[63:63] };
    end 
    if(N10599) begin
      { mem[4222:4222] } <= { data_i[62:62] };
    end 
    if(N10598) begin
      { mem[4221:4221] } <= { data_i[61:61] };
    end 
    if(N10597) begin
      { mem[4220:4220] } <= { data_i[60:60] };
    end 
    if(N10596) begin
      { mem[4219:4219] } <= { data_i[59:59] };
    end 
    if(N10595) begin
      { mem[4218:4218] } <= { data_i[58:58] };
    end 
    if(N10594) begin
      { mem[4217:4217] } <= { data_i[57:57] };
    end 
    if(N10593) begin
      { mem[4216:4216] } <= { data_i[56:56] };
    end 
    if(N10592) begin
      { mem[4215:4215] } <= { data_i[55:55] };
    end 
    if(N10591) begin
      { mem[4214:4214] } <= { data_i[54:54] };
    end 
    if(N10590) begin
      { mem[4213:4213] } <= { data_i[53:53] };
    end 
    if(N10589) begin
      { mem[4212:4212] } <= { data_i[52:52] };
    end 
    if(N10588) begin
      { mem[4211:4211] } <= { data_i[51:51] };
    end 
    if(N10587) begin
      { mem[4210:4210] } <= { data_i[50:50] };
    end 
    if(N10586) begin
      { mem[4209:4209] } <= { data_i[49:49] };
    end 
    if(N10585) begin
      { mem[4208:4208] } <= { data_i[48:48] };
    end 
    if(N10584) begin
      { mem[4207:4207] } <= { data_i[47:47] };
    end 
    if(N10583) begin
      { mem[4206:4206] } <= { data_i[46:46] };
    end 
    if(N10582) begin
      { mem[4205:4205] } <= { data_i[45:45] };
    end 
    if(N10581) begin
      { mem[4204:4204] } <= { data_i[44:44] };
    end 
    if(N10580) begin
      { mem[4203:4203] } <= { data_i[43:43] };
    end 
    if(N10579) begin
      { mem[4202:4202] } <= { data_i[42:42] };
    end 
    if(N10578) begin
      { mem[4201:4201] } <= { data_i[41:41] };
    end 
    if(N10577) begin
      { mem[4200:4200] } <= { data_i[40:40] };
    end 
    if(N10576) begin
      { mem[4199:4199] } <= { data_i[39:39] };
    end 
    if(N10575) begin
      { mem[4198:4198] } <= { data_i[38:38] };
    end 
    if(N10574) begin
      { mem[4197:4197] } <= { data_i[37:37] };
    end 
    if(N10573) begin
      { mem[4196:4196] } <= { data_i[36:36] };
    end 
    if(N10572) begin
      { mem[4195:4195] } <= { data_i[35:35] };
    end 
    if(N10571) begin
      { mem[4194:4194] } <= { data_i[34:34] };
    end 
    if(N10570) begin
      { mem[4193:4193] } <= { data_i[33:33] };
    end 
    if(N10569) begin
      { mem[4192:4192] } <= { data_i[32:32] };
    end 
    if(N10568) begin
      { mem[4191:4191] } <= { data_i[31:31] };
    end 
    if(N10567) begin
      { mem[4190:4190] } <= { data_i[30:30] };
    end 
    if(N10566) begin
      { mem[4189:4189] } <= { data_i[29:29] };
    end 
    if(N10565) begin
      { mem[4188:4188] } <= { data_i[28:28] };
    end 
    if(N10564) begin
      { mem[4187:4187] } <= { data_i[27:27] };
    end 
    if(N10563) begin
      { mem[4186:4186] } <= { data_i[26:26] };
    end 
    if(N10562) begin
      { mem[4185:4185] } <= { data_i[25:25] };
    end 
    if(N10561) begin
      { mem[4184:4184] } <= { data_i[24:24] };
    end 
    if(N10560) begin
      { mem[4183:4183] } <= { data_i[23:23] };
    end 
    if(N10559) begin
      { mem[4182:4182] } <= { data_i[22:22] };
    end 
    if(N10558) begin
      { mem[4181:4181] } <= { data_i[21:21] };
    end 
    if(N10557) begin
      { mem[4180:4180] } <= { data_i[20:20] };
    end 
    if(N10556) begin
      { mem[4179:4179] } <= { data_i[19:19] };
    end 
    if(N10555) begin
      { mem[4178:4178] } <= { data_i[18:18] };
    end 
    if(N10554) begin
      { mem[4177:4177] } <= { data_i[17:17] };
    end 
    if(N10553) begin
      { mem[4176:4176] } <= { data_i[16:16] };
    end 
    if(N10552) begin
      { mem[4175:4175] } <= { data_i[15:15] };
    end 
    if(N10551) begin
      { mem[4174:4174] } <= { data_i[14:14] };
    end 
    if(N10550) begin
      { mem[4173:4173] } <= { data_i[13:13] };
    end 
    if(N10549) begin
      { mem[4172:4172] } <= { data_i[12:12] };
    end 
    if(N10548) begin
      { mem[4171:4171] } <= { data_i[11:11] };
    end 
    if(N10547) begin
      { mem[4170:4170] } <= { data_i[10:10] };
    end 
    if(N10546) begin
      { mem[4169:4169] } <= { data_i[9:9] };
    end 
    if(N10545) begin
      { mem[4168:4168] } <= { data_i[8:8] };
    end 
    if(N10544) begin
      { mem[4167:4167] } <= { data_i[7:7] };
    end 
    if(N10543) begin
      { mem[4166:4166] } <= { data_i[6:6] };
    end 
    if(N10542) begin
      { mem[4165:4165] } <= { data_i[5:5] };
    end 
    if(N10541) begin
      { mem[4164:4164] } <= { data_i[4:4] };
    end 
    if(N10540) begin
      { mem[4163:4163] } <= { data_i[3:3] };
    end 
    if(N10539) begin
      { mem[4162:4162] } <= { data_i[2:2] };
    end 
    if(N10538) begin
      { mem[4161:4161] } <= { data_i[1:1] };
    end 
    if(N10537) begin
      { mem[4160:4160] } <= { data_i[0:0] };
    end 
    if(N10536) begin
      { mem[4159:4159] } <= { data_i[79:79] };
    end 
    if(N10535) begin
      { mem[4158:4158] } <= { data_i[78:78] };
    end 
    if(N10534) begin
      { mem[4157:4157] } <= { data_i[77:77] };
    end 
    if(N10533) begin
      { mem[4156:4156] } <= { data_i[76:76] };
    end 
    if(N10532) begin
      { mem[4155:4155] } <= { data_i[75:75] };
    end 
    if(N10531) begin
      { mem[4154:4154] } <= { data_i[74:74] };
    end 
    if(N10530) begin
      { mem[4153:4153] } <= { data_i[73:73] };
    end 
    if(N10529) begin
      { mem[4152:4152] } <= { data_i[72:72] };
    end 
    if(N10528) begin
      { mem[4151:4151] } <= { data_i[71:71] };
    end 
    if(N10527) begin
      { mem[4150:4150] } <= { data_i[70:70] };
    end 
    if(N10526) begin
      { mem[4149:4149] } <= { data_i[69:69] };
    end 
    if(N10525) begin
      { mem[4148:4148] } <= { data_i[68:68] };
    end 
    if(N10524) begin
      { mem[4147:4147] } <= { data_i[67:67] };
    end 
    if(N10523) begin
      { mem[4146:4146] } <= { data_i[66:66] };
    end 
    if(N10522) begin
      { mem[4145:4145] } <= { data_i[65:65] };
    end 
    if(N10521) begin
      { mem[4144:4144] } <= { data_i[64:64] };
    end 
    if(N10520) begin
      { mem[4143:4143] } <= { data_i[63:63] };
    end 
    if(N10519) begin
      { mem[4142:4142] } <= { data_i[62:62] };
    end 
    if(N10518) begin
      { mem[4141:4141] } <= { data_i[61:61] };
    end 
    if(N10517) begin
      { mem[4140:4140] } <= { data_i[60:60] };
    end 
    if(N10516) begin
      { mem[4139:4139] } <= { data_i[59:59] };
    end 
    if(N10515) begin
      { mem[4138:4138] } <= { data_i[58:58] };
    end 
    if(N10514) begin
      { mem[4137:4137] } <= { data_i[57:57] };
    end 
    if(N10513) begin
      { mem[4136:4136] } <= { data_i[56:56] };
    end 
    if(N10512) begin
      { mem[4135:4135] } <= { data_i[55:55] };
    end 
    if(N10511) begin
      { mem[4134:4134] } <= { data_i[54:54] };
    end 
    if(N10510) begin
      { mem[4133:4133] } <= { data_i[53:53] };
    end 
    if(N10509) begin
      { mem[4132:4132] } <= { data_i[52:52] };
    end 
    if(N10508) begin
      { mem[4131:4131] } <= { data_i[51:51] };
    end 
    if(N10507) begin
      { mem[4130:4130] } <= { data_i[50:50] };
    end 
    if(N10506) begin
      { mem[4129:4129] } <= { data_i[49:49] };
    end 
    if(N10505) begin
      { mem[4128:4128] } <= { data_i[48:48] };
    end 
    if(N10504) begin
      { mem[4127:4127] } <= { data_i[47:47] };
    end 
    if(N10503) begin
      { mem[4126:4126] } <= { data_i[46:46] };
    end 
    if(N10502) begin
      { mem[4125:4125] } <= { data_i[45:45] };
    end 
    if(N10501) begin
      { mem[4124:4124] } <= { data_i[44:44] };
    end 
    if(N10500) begin
      { mem[4123:4123] } <= { data_i[43:43] };
    end 
    if(N10499) begin
      { mem[4122:4122] } <= { data_i[42:42] };
    end 
    if(N10498) begin
      { mem[4121:4121] } <= { data_i[41:41] };
    end 
    if(N10497) begin
      { mem[4120:4120] } <= { data_i[40:40] };
    end 
    if(N10496) begin
      { mem[4119:4119] } <= { data_i[39:39] };
    end 
    if(N10495) begin
      { mem[4118:4118] } <= { data_i[38:38] };
    end 
    if(N10494) begin
      { mem[4117:4117] } <= { data_i[37:37] };
    end 
    if(N10493) begin
      { mem[4116:4116] } <= { data_i[36:36] };
    end 
    if(N10492) begin
      { mem[4115:4115] } <= { data_i[35:35] };
    end 
    if(N10491) begin
      { mem[4114:4114] } <= { data_i[34:34] };
    end 
    if(N10490) begin
      { mem[4113:4113] } <= { data_i[33:33] };
    end 
    if(N10489) begin
      { mem[4112:4112] } <= { data_i[32:32] };
    end 
    if(N10488) begin
      { mem[4111:4111] } <= { data_i[31:31] };
    end 
    if(N10487) begin
      { mem[4110:4110] } <= { data_i[30:30] };
    end 
    if(N10486) begin
      { mem[4109:4109] } <= { data_i[29:29] };
    end 
    if(N10485) begin
      { mem[4108:4108] } <= { data_i[28:28] };
    end 
    if(N10484) begin
      { mem[4107:4107] } <= { data_i[27:27] };
    end 
    if(N10483) begin
      { mem[4106:4106] } <= { data_i[26:26] };
    end 
    if(N10482) begin
      { mem[4105:4105] } <= { data_i[25:25] };
    end 
    if(N10481) begin
      { mem[4104:4104] } <= { data_i[24:24] };
    end 
    if(N10480) begin
      { mem[4103:4103] } <= { data_i[23:23] };
    end 
    if(N10479) begin
      { mem[4102:4102] } <= { data_i[22:22] };
    end 
    if(N10478) begin
      { mem[4101:4101] } <= { data_i[21:21] };
    end 
    if(N10477) begin
      { mem[4100:4100] } <= { data_i[20:20] };
    end 
    if(N10476) begin
      { mem[4099:4099] } <= { data_i[19:19] };
    end 
    if(N10475) begin
      { mem[4098:4098] } <= { data_i[18:18] };
    end 
    if(N10474) begin
      { mem[4097:4097] } <= { data_i[17:17] };
    end 
    if(N10473) begin
      { mem[4096:4096] } <= { data_i[16:16] };
    end 
    if(N10472) begin
      { mem[4095:4095] } <= { data_i[15:15] };
    end 
    if(N10471) begin
      { mem[4094:4094] } <= { data_i[14:14] };
    end 
    if(N10470) begin
      { mem[4093:4093] } <= { data_i[13:13] };
    end 
    if(N10469) begin
      { mem[4092:4092] } <= { data_i[12:12] };
    end 
    if(N10468) begin
      { mem[4091:4091] } <= { data_i[11:11] };
    end 
    if(N10467) begin
      { mem[4090:4090] } <= { data_i[10:10] };
    end 
    if(N10466) begin
      { mem[4089:4089] } <= { data_i[9:9] };
    end 
    if(N10465) begin
      { mem[4088:4088] } <= { data_i[8:8] };
    end 
    if(N10464) begin
      { mem[4087:4087] } <= { data_i[7:7] };
    end 
    if(N10463) begin
      { mem[4086:4086] } <= { data_i[6:6] };
    end 
    if(N10462) begin
      { mem[4085:4085] } <= { data_i[5:5] };
    end 
    if(N10461) begin
      { mem[4084:4084] } <= { data_i[4:4] };
    end 
    if(N10460) begin
      { mem[4083:4083] } <= { data_i[3:3] };
    end 
    if(N10459) begin
      { mem[4082:4082] } <= { data_i[2:2] };
    end 
    if(N10458) begin
      { mem[4081:4081] } <= { data_i[1:1] };
    end 
    if(N10457) begin
      { mem[4080:4080] } <= { data_i[0:0] };
    end 
    if(N10456) begin
      { mem[4079:4079] } <= { data_i[79:79] };
    end 
    if(N10455) begin
      { mem[4078:4078] } <= { data_i[78:78] };
    end 
    if(N10454) begin
      { mem[4077:4077] } <= { data_i[77:77] };
    end 
    if(N10453) begin
      { mem[4076:4076] } <= { data_i[76:76] };
    end 
    if(N10452) begin
      { mem[4075:4075] } <= { data_i[75:75] };
    end 
    if(N10451) begin
      { mem[4074:4074] } <= { data_i[74:74] };
    end 
    if(N10450) begin
      { mem[4073:4073] } <= { data_i[73:73] };
    end 
    if(N10449) begin
      { mem[4072:4072] } <= { data_i[72:72] };
    end 
    if(N10448) begin
      { mem[4071:4071] } <= { data_i[71:71] };
    end 
    if(N10447) begin
      { mem[4070:4070] } <= { data_i[70:70] };
    end 
    if(N10446) begin
      { mem[4069:4069] } <= { data_i[69:69] };
    end 
    if(N10445) begin
      { mem[4068:4068] } <= { data_i[68:68] };
    end 
    if(N10444) begin
      { mem[4067:4067] } <= { data_i[67:67] };
    end 
    if(N10443) begin
      { mem[4066:4066] } <= { data_i[66:66] };
    end 
    if(N10442) begin
      { mem[4065:4065] } <= { data_i[65:65] };
    end 
    if(N10441) begin
      { mem[4064:4064] } <= { data_i[64:64] };
    end 
    if(N10440) begin
      { mem[4063:4063] } <= { data_i[63:63] };
    end 
    if(N10439) begin
      { mem[4062:4062] } <= { data_i[62:62] };
    end 
    if(N10438) begin
      { mem[4061:4061] } <= { data_i[61:61] };
    end 
    if(N10437) begin
      { mem[4060:4060] } <= { data_i[60:60] };
    end 
    if(N10436) begin
      { mem[4059:4059] } <= { data_i[59:59] };
    end 
    if(N10435) begin
      { mem[4058:4058] } <= { data_i[58:58] };
    end 
    if(N10434) begin
      { mem[4057:4057] } <= { data_i[57:57] };
    end 
    if(N10433) begin
      { mem[4056:4056] } <= { data_i[56:56] };
    end 
    if(N10432) begin
      { mem[4055:4055] } <= { data_i[55:55] };
    end 
    if(N10431) begin
      { mem[4054:4054] } <= { data_i[54:54] };
    end 
    if(N10430) begin
      { mem[4053:4053] } <= { data_i[53:53] };
    end 
    if(N10429) begin
      { mem[4052:4052] } <= { data_i[52:52] };
    end 
    if(N10428) begin
      { mem[4051:4051] } <= { data_i[51:51] };
    end 
    if(N10427) begin
      { mem[4050:4050] } <= { data_i[50:50] };
    end 
    if(N10426) begin
      { mem[4049:4049] } <= { data_i[49:49] };
    end 
    if(N10425) begin
      { mem[4048:4048] } <= { data_i[48:48] };
    end 
    if(N10424) begin
      { mem[4047:4047] } <= { data_i[47:47] };
    end 
    if(N10423) begin
      { mem[4046:4046] } <= { data_i[46:46] };
    end 
    if(N10422) begin
      { mem[4045:4045] } <= { data_i[45:45] };
    end 
    if(N10421) begin
      { mem[4044:4044] } <= { data_i[44:44] };
    end 
    if(N10420) begin
      { mem[4043:4043] } <= { data_i[43:43] };
    end 
    if(N10419) begin
      { mem[4042:4042] } <= { data_i[42:42] };
    end 
    if(N10418) begin
      { mem[4041:4041] } <= { data_i[41:41] };
    end 
    if(N10417) begin
      { mem[4040:4040] } <= { data_i[40:40] };
    end 
    if(N10416) begin
      { mem[4039:4039] } <= { data_i[39:39] };
    end 
    if(N10415) begin
      { mem[4038:4038] } <= { data_i[38:38] };
    end 
    if(N10414) begin
      { mem[4037:4037] } <= { data_i[37:37] };
    end 
    if(N10413) begin
      { mem[4036:4036] } <= { data_i[36:36] };
    end 
    if(N10412) begin
      { mem[4035:4035] } <= { data_i[35:35] };
    end 
    if(N10411) begin
      { mem[4034:4034] } <= { data_i[34:34] };
    end 
    if(N10410) begin
      { mem[4033:4033] } <= { data_i[33:33] };
    end 
    if(N10409) begin
      { mem[4032:4032] } <= { data_i[32:32] };
    end 
    if(N10408) begin
      { mem[4031:4031] } <= { data_i[31:31] };
    end 
    if(N10407) begin
      { mem[4030:4030] } <= { data_i[30:30] };
    end 
    if(N10406) begin
      { mem[4029:4029] } <= { data_i[29:29] };
    end 
    if(N10405) begin
      { mem[4028:4028] } <= { data_i[28:28] };
    end 
    if(N10404) begin
      { mem[4027:4027] } <= { data_i[27:27] };
    end 
    if(N10403) begin
      { mem[4026:4026] } <= { data_i[26:26] };
    end 
    if(N10402) begin
      { mem[4025:4025] } <= { data_i[25:25] };
    end 
    if(N10401) begin
      { mem[4024:4024] } <= { data_i[24:24] };
    end 
    if(N10400) begin
      { mem[4023:4023] } <= { data_i[23:23] };
    end 
    if(N10399) begin
      { mem[4022:4022] } <= { data_i[22:22] };
    end 
    if(N10398) begin
      { mem[4021:4021] } <= { data_i[21:21] };
    end 
    if(N10397) begin
      { mem[4020:4020] } <= { data_i[20:20] };
    end 
    if(N10396) begin
      { mem[4019:4019] } <= { data_i[19:19] };
    end 
    if(N10395) begin
      { mem[4018:4018] } <= { data_i[18:18] };
    end 
    if(N10394) begin
      { mem[4017:4017] } <= { data_i[17:17] };
    end 
    if(N10393) begin
      { mem[4016:4016] } <= { data_i[16:16] };
    end 
    if(N10392) begin
      { mem[4015:4015] } <= { data_i[15:15] };
    end 
    if(N10391) begin
      { mem[4014:4014] } <= { data_i[14:14] };
    end 
    if(N10390) begin
      { mem[4013:4013] } <= { data_i[13:13] };
    end 
    if(N10389) begin
      { mem[4012:4012] } <= { data_i[12:12] };
    end 
    if(N10388) begin
      { mem[4011:4011] } <= { data_i[11:11] };
    end 
    if(N10387) begin
      { mem[4010:4010] } <= { data_i[10:10] };
    end 
    if(N10386) begin
      { mem[4009:4009] } <= { data_i[9:9] };
    end 
    if(N10385) begin
      { mem[4008:4008] } <= { data_i[8:8] };
    end 
    if(N10384) begin
      { mem[4007:4007] } <= { data_i[7:7] };
    end 
    if(N10383) begin
      { mem[4006:4006] } <= { data_i[6:6] };
    end 
    if(N10382) begin
      { mem[4005:4005] } <= { data_i[5:5] };
    end 
    if(N10381) begin
      { mem[4004:4004] } <= { data_i[4:4] };
    end 
    if(N10380) begin
      { mem[4003:4003] } <= { data_i[3:3] };
    end 
    if(N10379) begin
      { mem[4002:4002] } <= { data_i[2:2] };
    end 
    if(N10378) begin
      { mem[4001:4001] } <= { data_i[1:1] };
    end 
    if(N10377) begin
      { mem[4000:4000] } <= { data_i[0:0] };
    end 
    if(N10376) begin
      { mem[3999:3999] } <= { data_i[79:79] };
    end 
    if(N10375) begin
      { mem[3998:3998] } <= { data_i[78:78] };
    end 
    if(N10374) begin
      { mem[3997:3997] } <= { data_i[77:77] };
    end 
    if(N10373) begin
      { mem[3996:3996] } <= { data_i[76:76] };
    end 
    if(N10372) begin
      { mem[3995:3995] } <= { data_i[75:75] };
    end 
    if(N10371) begin
      { mem[3994:3994] } <= { data_i[74:74] };
    end 
    if(N10370) begin
      { mem[3993:3993] } <= { data_i[73:73] };
    end 
    if(N10369) begin
      { mem[3992:3992] } <= { data_i[72:72] };
    end 
    if(N10368) begin
      { mem[3991:3991] } <= { data_i[71:71] };
    end 
    if(N10367) begin
      { mem[3990:3990] } <= { data_i[70:70] };
    end 
    if(N10366) begin
      { mem[3989:3989] } <= { data_i[69:69] };
    end 
    if(N10365) begin
      { mem[3988:3988] } <= { data_i[68:68] };
    end 
    if(N10364) begin
      { mem[3987:3987] } <= { data_i[67:67] };
    end 
    if(N10363) begin
      { mem[3986:3986] } <= { data_i[66:66] };
    end 
    if(N10362) begin
      { mem[3985:3985] } <= { data_i[65:65] };
    end 
    if(N10361) begin
      { mem[3984:3984] } <= { data_i[64:64] };
    end 
    if(N10360) begin
      { mem[3983:3983] } <= { data_i[63:63] };
    end 
    if(N10359) begin
      { mem[3982:3982] } <= { data_i[62:62] };
    end 
    if(N10358) begin
      { mem[3981:3981] } <= { data_i[61:61] };
    end 
    if(N10357) begin
      { mem[3980:3980] } <= { data_i[60:60] };
    end 
    if(N10356) begin
      { mem[3979:3979] } <= { data_i[59:59] };
    end 
    if(N10355) begin
      { mem[3978:3978] } <= { data_i[58:58] };
    end 
    if(N10354) begin
      { mem[3977:3977] } <= { data_i[57:57] };
    end 
    if(N10353) begin
      { mem[3976:3976] } <= { data_i[56:56] };
    end 
    if(N10352) begin
      { mem[3975:3975] } <= { data_i[55:55] };
    end 
    if(N10351) begin
      { mem[3974:3974] } <= { data_i[54:54] };
    end 
    if(N10350) begin
      { mem[3973:3973] } <= { data_i[53:53] };
    end 
    if(N10349) begin
      { mem[3972:3972] } <= { data_i[52:52] };
    end 
    if(N10348) begin
      { mem[3971:3971] } <= { data_i[51:51] };
    end 
    if(N10347) begin
      { mem[3970:3970] } <= { data_i[50:50] };
    end 
    if(N10346) begin
      { mem[3969:3969] } <= { data_i[49:49] };
    end 
    if(N10345) begin
      { mem[3968:3968] } <= { data_i[48:48] };
    end 
    if(N10344) begin
      { mem[3967:3967] } <= { data_i[47:47] };
    end 
    if(N10343) begin
      { mem[3966:3966] } <= { data_i[46:46] };
    end 
    if(N10342) begin
      { mem[3965:3965] } <= { data_i[45:45] };
    end 
    if(N10341) begin
      { mem[3964:3964] } <= { data_i[44:44] };
    end 
    if(N10340) begin
      { mem[3963:3963] } <= { data_i[43:43] };
    end 
    if(N10339) begin
      { mem[3962:3962] } <= { data_i[42:42] };
    end 
    if(N10338) begin
      { mem[3961:3961] } <= { data_i[41:41] };
    end 
    if(N10337) begin
      { mem[3960:3960] } <= { data_i[40:40] };
    end 
    if(N10336) begin
      { mem[3959:3959] } <= { data_i[39:39] };
    end 
    if(N10335) begin
      { mem[3958:3958] } <= { data_i[38:38] };
    end 
    if(N10334) begin
      { mem[3957:3957] } <= { data_i[37:37] };
    end 
    if(N10333) begin
      { mem[3956:3956] } <= { data_i[36:36] };
    end 
    if(N10332) begin
      { mem[3955:3955] } <= { data_i[35:35] };
    end 
    if(N10331) begin
      { mem[3954:3954] } <= { data_i[34:34] };
    end 
    if(N10330) begin
      { mem[3953:3953] } <= { data_i[33:33] };
    end 
    if(N10329) begin
      { mem[3952:3952] } <= { data_i[32:32] };
    end 
    if(N10328) begin
      { mem[3951:3951] } <= { data_i[31:31] };
    end 
    if(N10327) begin
      { mem[3950:3950] } <= { data_i[30:30] };
    end 
    if(N10326) begin
      { mem[3949:3949] } <= { data_i[29:29] };
    end 
    if(N10325) begin
      { mem[3948:3948] } <= { data_i[28:28] };
    end 
    if(N10324) begin
      { mem[3947:3947] } <= { data_i[27:27] };
    end 
    if(N10323) begin
      { mem[3946:3946] } <= { data_i[26:26] };
    end 
    if(N10322) begin
      { mem[3945:3945] } <= { data_i[25:25] };
    end 
    if(N10321) begin
      { mem[3944:3944] } <= { data_i[24:24] };
    end 
    if(N10320) begin
      { mem[3943:3943] } <= { data_i[23:23] };
    end 
    if(N10319) begin
      { mem[3942:3942] } <= { data_i[22:22] };
    end 
    if(N10318) begin
      { mem[3941:3941] } <= { data_i[21:21] };
    end 
    if(N10317) begin
      { mem[3940:3940] } <= { data_i[20:20] };
    end 
    if(N10316) begin
      { mem[3939:3939] } <= { data_i[19:19] };
    end 
    if(N10315) begin
      { mem[3938:3938] } <= { data_i[18:18] };
    end 
    if(N10314) begin
      { mem[3937:3937] } <= { data_i[17:17] };
    end 
    if(N10313) begin
      { mem[3936:3936] } <= { data_i[16:16] };
    end 
    if(N10312) begin
      { mem[3935:3935] } <= { data_i[15:15] };
    end 
    if(N10311) begin
      { mem[3934:3934] } <= { data_i[14:14] };
    end 
    if(N10310) begin
      { mem[3933:3933] } <= { data_i[13:13] };
    end 
    if(N10309) begin
      { mem[3932:3932] } <= { data_i[12:12] };
    end 
    if(N10308) begin
      { mem[3931:3931] } <= { data_i[11:11] };
    end 
    if(N10307) begin
      { mem[3930:3930] } <= { data_i[10:10] };
    end 
    if(N10306) begin
      { mem[3929:3929] } <= { data_i[9:9] };
    end 
    if(N10305) begin
      { mem[3928:3928] } <= { data_i[8:8] };
    end 
    if(N10304) begin
      { mem[3927:3927] } <= { data_i[7:7] };
    end 
    if(N10303) begin
      { mem[3926:3926] } <= { data_i[6:6] };
    end 
    if(N10302) begin
      { mem[3925:3925] } <= { data_i[5:5] };
    end 
    if(N10301) begin
      { mem[3924:3924] } <= { data_i[4:4] };
    end 
    if(N10300) begin
      { mem[3923:3923] } <= { data_i[3:3] };
    end 
    if(N10299) begin
      { mem[3922:3922] } <= { data_i[2:2] };
    end 
    if(N10298) begin
      { mem[3921:3921] } <= { data_i[1:1] };
    end 
    if(N10297) begin
      { mem[3920:3920] } <= { data_i[0:0] };
    end 
    if(N10296) begin
      { mem[3919:3919] } <= { data_i[79:79] };
    end 
    if(N10295) begin
      { mem[3918:3918] } <= { data_i[78:78] };
    end 
    if(N10294) begin
      { mem[3917:3917] } <= { data_i[77:77] };
    end 
    if(N10293) begin
      { mem[3916:3916] } <= { data_i[76:76] };
    end 
    if(N10292) begin
      { mem[3915:3915] } <= { data_i[75:75] };
    end 
    if(N10291) begin
      { mem[3914:3914] } <= { data_i[74:74] };
    end 
    if(N10290) begin
      { mem[3913:3913] } <= { data_i[73:73] };
    end 
    if(N10289) begin
      { mem[3912:3912] } <= { data_i[72:72] };
    end 
    if(N10288) begin
      { mem[3911:3911] } <= { data_i[71:71] };
    end 
    if(N10287) begin
      { mem[3910:3910] } <= { data_i[70:70] };
    end 
    if(N10286) begin
      { mem[3909:3909] } <= { data_i[69:69] };
    end 
    if(N10285) begin
      { mem[3908:3908] } <= { data_i[68:68] };
    end 
    if(N10284) begin
      { mem[3907:3907] } <= { data_i[67:67] };
    end 
    if(N10283) begin
      { mem[3906:3906] } <= { data_i[66:66] };
    end 
    if(N10282) begin
      { mem[3905:3905] } <= { data_i[65:65] };
    end 
    if(N10281) begin
      { mem[3904:3904] } <= { data_i[64:64] };
    end 
    if(N10280) begin
      { mem[3903:3903] } <= { data_i[63:63] };
    end 
    if(N10279) begin
      { mem[3902:3902] } <= { data_i[62:62] };
    end 
    if(N10278) begin
      { mem[3901:3901] } <= { data_i[61:61] };
    end 
    if(N10277) begin
      { mem[3900:3900] } <= { data_i[60:60] };
    end 
    if(N10276) begin
      { mem[3899:3899] } <= { data_i[59:59] };
    end 
    if(N10275) begin
      { mem[3898:3898] } <= { data_i[58:58] };
    end 
    if(N10274) begin
      { mem[3897:3897] } <= { data_i[57:57] };
    end 
    if(N10273) begin
      { mem[3896:3896] } <= { data_i[56:56] };
    end 
    if(N10272) begin
      { mem[3895:3895] } <= { data_i[55:55] };
    end 
    if(N10271) begin
      { mem[3894:3894] } <= { data_i[54:54] };
    end 
    if(N10270) begin
      { mem[3893:3893] } <= { data_i[53:53] };
    end 
    if(N10269) begin
      { mem[3892:3892] } <= { data_i[52:52] };
    end 
    if(N10268) begin
      { mem[3891:3891] } <= { data_i[51:51] };
    end 
    if(N10267) begin
      { mem[3890:3890] } <= { data_i[50:50] };
    end 
    if(N10266) begin
      { mem[3889:3889] } <= { data_i[49:49] };
    end 
    if(N10265) begin
      { mem[3888:3888] } <= { data_i[48:48] };
    end 
    if(N10264) begin
      { mem[3887:3887] } <= { data_i[47:47] };
    end 
    if(N10263) begin
      { mem[3886:3886] } <= { data_i[46:46] };
    end 
    if(N10262) begin
      { mem[3885:3885] } <= { data_i[45:45] };
    end 
    if(N10261) begin
      { mem[3884:3884] } <= { data_i[44:44] };
    end 
    if(N10260) begin
      { mem[3883:3883] } <= { data_i[43:43] };
    end 
    if(N10259) begin
      { mem[3882:3882] } <= { data_i[42:42] };
    end 
    if(N10258) begin
      { mem[3881:3881] } <= { data_i[41:41] };
    end 
    if(N10257) begin
      { mem[3880:3880] } <= { data_i[40:40] };
    end 
    if(N10256) begin
      { mem[3879:3879] } <= { data_i[39:39] };
    end 
    if(N10255) begin
      { mem[3878:3878] } <= { data_i[38:38] };
    end 
    if(N10254) begin
      { mem[3877:3877] } <= { data_i[37:37] };
    end 
    if(N10253) begin
      { mem[3876:3876] } <= { data_i[36:36] };
    end 
    if(N10252) begin
      { mem[3875:3875] } <= { data_i[35:35] };
    end 
    if(N10251) begin
      { mem[3874:3874] } <= { data_i[34:34] };
    end 
    if(N10250) begin
      { mem[3873:3873] } <= { data_i[33:33] };
    end 
    if(N10249) begin
      { mem[3872:3872] } <= { data_i[32:32] };
    end 
    if(N10248) begin
      { mem[3871:3871] } <= { data_i[31:31] };
    end 
    if(N10247) begin
      { mem[3870:3870] } <= { data_i[30:30] };
    end 
    if(N10246) begin
      { mem[3869:3869] } <= { data_i[29:29] };
    end 
    if(N10245) begin
      { mem[3868:3868] } <= { data_i[28:28] };
    end 
    if(N10244) begin
      { mem[3867:3867] } <= { data_i[27:27] };
    end 
    if(N10243) begin
      { mem[3866:3866] } <= { data_i[26:26] };
    end 
    if(N10242) begin
      { mem[3865:3865] } <= { data_i[25:25] };
    end 
    if(N10241) begin
      { mem[3864:3864] } <= { data_i[24:24] };
    end 
    if(N10240) begin
      { mem[3863:3863] } <= { data_i[23:23] };
    end 
    if(N10239) begin
      { mem[3862:3862] } <= { data_i[22:22] };
    end 
    if(N10238) begin
      { mem[3861:3861] } <= { data_i[21:21] };
    end 
    if(N10237) begin
      { mem[3860:3860] } <= { data_i[20:20] };
    end 
    if(N10236) begin
      { mem[3859:3859] } <= { data_i[19:19] };
    end 
    if(N10235) begin
      { mem[3858:3858] } <= { data_i[18:18] };
    end 
    if(N10234) begin
      { mem[3857:3857] } <= { data_i[17:17] };
    end 
    if(N10233) begin
      { mem[3856:3856] } <= { data_i[16:16] };
    end 
    if(N10232) begin
      { mem[3855:3855] } <= { data_i[15:15] };
    end 
    if(N10231) begin
      { mem[3854:3854] } <= { data_i[14:14] };
    end 
    if(N10230) begin
      { mem[3853:3853] } <= { data_i[13:13] };
    end 
    if(N10229) begin
      { mem[3852:3852] } <= { data_i[12:12] };
    end 
    if(N10228) begin
      { mem[3851:3851] } <= { data_i[11:11] };
    end 
    if(N10227) begin
      { mem[3850:3850] } <= { data_i[10:10] };
    end 
    if(N10226) begin
      { mem[3849:3849] } <= { data_i[9:9] };
    end 
    if(N10225) begin
      { mem[3848:3848] } <= { data_i[8:8] };
    end 
    if(N10224) begin
      { mem[3847:3847] } <= { data_i[7:7] };
    end 
    if(N10223) begin
      { mem[3846:3846] } <= { data_i[6:6] };
    end 
    if(N10222) begin
      { mem[3845:3845] } <= { data_i[5:5] };
    end 
    if(N10221) begin
      { mem[3844:3844] } <= { data_i[4:4] };
    end 
    if(N10220) begin
      { mem[3843:3843] } <= { data_i[3:3] };
    end 
    if(N10219) begin
      { mem[3842:3842] } <= { data_i[2:2] };
    end 
    if(N10218) begin
      { mem[3841:3841] } <= { data_i[1:1] };
    end 
    if(N10217) begin
      { mem[3840:3840] } <= { data_i[0:0] };
    end 
    if(N10216) begin
      { mem[3839:3839] } <= { data_i[79:79] };
    end 
    if(N10215) begin
      { mem[3838:3838] } <= { data_i[78:78] };
    end 
    if(N10214) begin
      { mem[3837:3837] } <= { data_i[77:77] };
    end 
    if(N10213) begin
      { mem[3836:3836] } <= { data_i[76:76] };
    end 
    if(N10212) begin
      { mem[3835:3835] } <= { data_i[75:75] };
    end 
    if(N10211) begin
      { mem[3834:3834] } <= { data_i[74:74] };
    end 
    if(N10210) begin
      { mem[3833:3833] } <= { data_i[73:73] };
    end 
    if(N10209) begin
      { mem[3832:3832] } <= { data_i[72:72] };
    end 
    if(N10208) begin
      { mem[3831:3831] } <= { data_i[71:71] };
    end 
    if(N10207) begin
      { mem[3830:3830] } <= { data_i[70:70] };
    end 
    if(N10206) begin
      { mem[3829:3829] } <= { data_i[69:69] };
    end 
    if(N10205) begin
      { mem[3828:3828] } <= { data_i[68:68] };
    end 
    if(N10204) begin
      { mem[3827:3827] } <= { data_i[67:67] };
    end 
    if(N10203) begin
      { mem[3826:3826] } <= { data_i[66:66] };
    end 
    if(N10202) begin
      { mem[3825:3825] } <= { data_i[65:65] };
    end 
    if(N10201) begin
      { mem[3824:3824] } <= { data_i[64:64] };
    end 
    if(N10200) begin
      { mem[3823:3823] } <= { data_i[63:63] };
    end 
    if(N10199) begin
      { mem[3822:3822] } <= { data_i[62:62] };
    end 
    if(N10198) begin
      { mem[3821:3821] } <= { data_i[61:61] };
    end 
    if(N10197) begin
      { mem[3820:3820] } <= { data_i[60:60] };
    end 
    if(N10196) begin
      { mem[3819:3819] } <= { data_i[59:59] };
    end 
    if(N10195) begin
      { mem[3818:3818] } <= { data_i[58:58] };
    end 
    if(N10194) begin
      { mem[3817:3817] } <= { data_i[57:57] };
    end 
    if(N10193) begin
      { mem[3816:3816] } <= { data_i[56:56] };
    end 
    if(N10192) begin
      { mem[3815:3815] } <= { data_i[55:55] };
    end 
    if(N10191) begin
      { mem[3814:3814] } <= { data_i[54:54] };
    end 
    if(N10190) begin
      { mem[3813:3813] } <= { data_i[53:53] };
    end 
    if(N10189) begin
      { mem[3812:3812] } <= { data_i[52:52] };
    end 
    if(N10188) begin
      { mem[3811:3811] } <= { data_i[51:51] };
    end 
    if(N10187) begin
      { mem[3810:3810] } <= { data_i[50:50] };
    end 
    if(N10186) begin
      { mem[3809:3809] } <= { data_i[49:49] };
    end 
    if(N10185) begin
      { mem[3808:3808] } <= { data_i[48:48] };
    end 
    if(N10184) begin
      { mem[3807:3807] } <= { data_i[47:47] };
    end 
    if(N10183) begin
      { mem[3806:3806] } <= { data_i[46:46] };
    end 
    if(N10182) begin
      { mem[3805:3805] } <= { data_i[45:45] };
    end 
    if(N10181) begin
      { mem[3804:3804] } <= { data_i[44:44] };
    end 
    if(N10180) begin
      { mem[3803:3803] } <= { data_i[43:43] };
    end 
    if(N10179) begin
      { mem[3802:3802] } <= { data_i[42:42] };
    end 
    if(N10178) begin
      { mem[3801:3801] } <= { data_i[41:41] };
    end 
    if(N10177) begin
      { mem[3800:3800] } <= { data_i[40:40] };
    end 
    if(N10176) begin
      { mem[3799:3799] } <= { data_i[39:39] };
    end 
    if(N10175) begin
      { mem[3798:3798] } <= { data_i[38:38] };
    end 
    if(N10174) begin
      { mem[3797:3797] } <= { data_i[37:37] };
    end 
    if(N10173) begin
      { mem[3796:3796] } <= { data_i[36:36] };
    end 
    if(N10172) begin
      { mem[3795:3795] } <= { data_i[35:35] };
    end 
    if(N10171) begin
      { mem[3794:3794] } <= { data_i[34:34] };
    end 
    if(N10170) begin
      { mem[3793:3793] } <= { data_i[33:33] };
    end 
    if(N10169) begin
      { mem[3792:3792] } <= { data_i[32:32] };
    end 
    if(N10168) begin
      { mem[3791:3791] } <= { data_i[31:31] };
    end 
    if(N10167) begin
      { mem[3790:3790] } <= { data_i[30:30] };
    end 
    if(N10166) begin
      { mem[3789:3789] } <= { data_i[29:29] };
    end 
    if(N10165) begin
      { mem[3788:3788] } <= { data_i[28:28] };
    end 
    if(N10164) begin
      { mem[3787:3787] } <= { data_i[27:27] };
    end 
    if(N10163) begin
      { mem[3786:3786] } <= { data_i[26:26] };
    end 
    if(N10162) begin
      { mem[3785:3785] } <= { data_i[25:25] };
    end 
    if(N10161) begin
      { mem[3784:3784] } <= { data_i[24:24] };
    end 
    if(N10160) begin
      { mem[3783:3783] } <= { data_i[23:23] };
    end 
    if(N10159) begin
      { mem[3782:3782] } <= { data_i[22:22] };
    end 
    if(N10158) begin
      { mem[3781:3781] } <= { data_i[21:21] };
    end 
    if(N10157) begin
      { mem[3780:3780] } <= { data_i[20:20] };
    end 
    if(N10156) begin
      { mem[3779:3779] } <= { data_i[19:19] };
    end 
    if(N10155) begin
      { mem[3778:3778] } <= { data_i[18:18] };
    end 
    if(N10154) begin
      { mem[3777:3777] } <= { data_i[17:17] };
    end 
    if(N10153) begin
      { mem[3776:3776] } <= { data_i[16:16] };
    end 
    if(N10152) begin
      { mem[3775:3775] } <= { data_i[15:15] };
    end 
    if(N10151) begin
      { mem[3774:3774] } <= { data_i[14:14] };
    end 
    if(N10150) begin
      { mem[3773:3773] } <= { data_i[13:13] };
    end 
    if(N10149) begin
      { mem[3772:3772] } <= { data_i[12:12] };
    end 
    if(N10148) begin
      { mem[3771:3771] } <= { data_i[11:11] };
    end 
    if(N10147) begin
      { mem[3770:3770] } <= { data_i[10:10] };
    end 
    if(N10146) begin
      { mem[3769:3769] } <= { data_i[9:9] };
    end 
    if(N10145) begin
      { mem[3768:3768] } <= { data_i[8:8] };
    end 
    if(N10144) begin
      { mem[3767:3767] } <= { data_i[7:7] };
    end 
    if(N10143) begin
      { mem[3766:3766] } <= { data_i[6:6] };
    end 
    if(N10142) begin
      { mem[3765:3765] } <= { data_i[5:5] };
    end 
    if(N10141) begin
      { mem[3764:3764] } <= { data_i[4:4] };
    end 
    if(N10140) begin
      { mem[3763:3763] } <= { data_i[3:3] };
    end 
    if(N10139) begin
      { mem[3762:3762] } <= { data_i[2:2] };
    end 
    if(N10138) begin
      { mem[3761:3761] } <= { data_i[1:1] };
    end 
    if(N10137) begin
      { mem[3760:3760] } <= { data_i[0:0] };
    end 
    if(N10136) begin
      { mem[3759:3759] } <= { data_i[79:79] };
    end 
    if(N10135) begin
      { mem[3758:3758] } <= { data_i[78:78] };
    end 
    if(N10134) begin
      { mem[3757:3757] } <= { data_i[77:77] };
    end 
    if(N10133) begin
      { mem[3756:3756] } <= { data_i[76:76] };
    end 
    if(N10132) begin
      { mem[3755:3755] } <= { data_i[75:75] };
    end 
    if(N10131) begin
      { mem[3754:3754] } <= { data_i[74:74] };
    end 
    if(N10130) begin
      { mem[3753:3753] } <= { data_i[73:73] };
    end 
    if(N10129) begin
      { mem[3752:3752] } <= { data_i[72:72] };
    end 
    if(N10128) begin
      { mem[3751:3751] } <= { data_i[71:71] };
    end 
    if(N10127) begin
      { mem[3750:3750] } <= { data_i[70:70] };
    end 
    if(N10126) begin
      { mem[3749:3749] } <= { data_i[69:69] };
    end 
    if(N10125) begin
      { mem[3748:3748] } <= { data_i[68:68] };
    end 
    if(N10124) begin
      { mem[3747:3747] } <= { data_i[67:67] };
    end 
    if(N10123) begin
      { mem[3746:3746] } <= { data_i[66:66] };
    end 
    if(N10122) begin
      { mem[3745:3745] } <= { data_i[65:65] };
    end 
    if(N10121) begin
      { mem[3744:3744] } <= { data_i[64:64] };
    end 
    if(N10120) begin
      { mem[3743:3743] } <= { data_i[63:63] };
    end 
    if(N10119) begin
      { mem[3742:3742] } <= { data_i[62:62] };
    end 
    if(N10118) begin
      { mem[3741:3741] } <= { data_i[61:61] };
    end 
    if(N10117) begin
      { mem[3740:3740] } <= { data_i[60:60] };
    end 
    if(N10116) begin
      { mem[3739:3739] } <= { data_i[59:59] };
    end 
    if(N10115) begin
      { mem[3738:3738] } <= { data_i[58:58] };
    end 
    if(N10114) begin
      { mem[3737:3737] } <= { data_i[57:57] };
    end 
    if(N10113) begin
      { mem[3736:3736] } <= { data_i[56:56] };
    end 
    if(N10112) begin
      { mem[3735:3735] } <= { data_i[55:55] };
    end 
    if(N10111) begin
      { mem[3734:3734] } <= { data_i[54:54] };
    end 
    if(N10110) begin
      { mem[3733:3733] } <= { data_i[53:53] };
    end 
    if(N10109) begin
      { mem[3732:3732] } <= { data_i[52:52] };
    end 
    if(N10108) begin
      { mem[3731:3731] } <= { data_i[51:51] };
    end 
    if(N10107) begin
      { mem[3730:3730] } <= { data_i[50:50] };
    end 
    if(N10106) begin
      { mem[3729:3729] } <= { data_i[49:49] };
    end 
    if(N10105) begin
      { mem[3728:3728] } <= { data_i[48:48] };
    end 
    if(N10104) begin
      { mem[3727:3727] } <= { data_i[47:47] };
    end 
    if(N10103) begin
      { mem[3726:3726] } <= { data_i[46:46] };
    end 
    if(N10102) begin
      { mem[3725:3725] } <= { data_i[45:45] };
    end 
    if(N10101) begin
      { mem[3724:3724] } <= { data_i[44:44] };
    end 
    if(N10100) begin
      { mem[3723:3723] } <= { data_i[43:43] };
    end 
    if(N10099) begin
      { mem[3722:3722] } <= { data_i[42:42] };
    end 
    if(N10098) begin
      { mem[3721:3721] } <= { data_i[41:41] };
    end 
    if(N10097) begin
      { mem[3720:3720] } <= { data_i[40:40] };
    end 
    if(N10096) begin
      { mem[3719:3719] } <= { data_i[39:39] };
    end 
    if(N10095) begin
      { mem[3718:3718] } <= { data_i[38:38] };
    end 
    if(N10094) begin
      { mem[3717:3717] } <= { data_i[37:37] };
    end 
    if(N10093) begin
      { mem[3716:3716] } <= { data_i[36:36] };
    end 
    if(N10092) begin
      { mem[3715:3715] } <= { data_i[35:35] };
    end 
    if(N10091) begin
      { mem[3714:3714] } <= { data_i[34:34] };
    end 
    if(N10090) begin
      { mem[3713:3713] } <= { data_i[33:33] };
    end 
    if(N10089) begin
      { mem[3712:3712] } <= { data_i[32:32] };
    end 
    if(N10088) begin
      { mem[3711:3711] } <= { data_i[31:31] };
    end 
    if(N10087) begin
      { mem[3710:3710] } <= { data_i[30:30] };
    end 
    if(N10086) begin
      { mem[3709:3709] } <= { data_i[29:29] };
    end 
    if(N10085) begin
      { mem[3708:3708] } <= { data_i[28:28] };
    end 
    if(N10084) begin
      { mem[3707:3707] } <= { data_i[27:27] };
    end 
    if(N10083) begin
      { mem[3706:3706] } <= { data_i[26:26] };
    end 
    if(N10082) begin
      { mem[3705:3705] } <= { data_i[25:25] };
    end 
    if(N10081) begin
      { mem[3704:3704] } <= { data_i[24:24] };
    end 
    if(N10080) begin
      { mem[3703:3703] } <= { data_i[23:23] };
    end 
    if(N10079) begin
      { mem[3702:3702] } <= { data_i[22:22] };
    end 
    if(N10078) begin
      { mem[3701:3701] } <= { data_i[21:21] };
    end 
    if(N10077) begin
      { mem[3700:3700] } <= { data_i[20:20] };
    end 
    if(N10076) begin
      { mem[3699:3699] } <= { data_i[19:19] };
    end 
    if(N10075) begin
      { mem[3698:3698] } <= { data_i[18:18] };
    end 
    if(N10074) begin
      { mem[3697:3697] } <= { data_i[17:17] };
    end 
    if(N10073) begin
      { mem[3696:3696] } <= { data_i[16:16] };
    end 
    if(N10072) begin
      { mem[3695:3695] } <= { data_i[15:15] };
    end 
    if(N10071) begin
      { mem[3694:3694] } <= { data_i[14:14] };
    end 
    if(N10070) begin
      { mem[3693:3693] } <= { data_i[13:13] };
    end 
    if(N10069) begin
      { mem[3692:3692] } <= { data_i[12:12] };
    end 
    if(N10068) begin
      { mem[3691:3691] } <= { data_i[11:11] };
    end 
    if(N10067) begin
      { mem[3690:3690] } <= { data_i[10:10] };
    end 
    if(N10066) begin
      { mem[3689:3689] } <= { data_i[9:9] };
    end 
    if(N10065) begin
      { mem[3688:3688] } <= { data_i[8:8] };
    end 
    if(N10064) begin
      { mem[3687:3687] } <= { data_i[7:7] };
    end 
    if(N10063) begin
      { mem[3686:3686] } <= { data_i[6:6] };
    end 
    if(N10062) begin
      { mem[3685:3685] } <= { data_i[5:5] };
    end 
    if(N10061) begin
      { mem[3684:3684] } <= { data_i[4:4] };
    end 
    if(N10060) begin
      { mem[3683:3683] } <= { data_i[3:3] };
    end 
    if(N10059) begin
      { mem[3682:3682] } <= { data_i[2:2] };
    end 
    if(N10058) begin
      { mem[3681:3681] } <= { data_i[1:1] };
    end 
    if(N10057) begin
      { mem[3680:3680] } <= { data_i[0:0] };
    end 
    if(N10056) begin
      { mem[3679:3679] } <= { data_i[79:79] };
    end 
    if(N10055) begin
      { mem[3678:3678] } <= { data_i[78:78] };
    end 
    if(N10054) begin
      { mem[3677:3677] } <= { data_i[77:77] };
    end 
    if(N10053) begin
      { mem[3676:3676] } <= { data_i[76:76] };
    end 
    if(N10052) begin
      { mem[3675:3675] } <= { data_i[75:75] };
    end 
    if(N10051) begin
      { mem[3674:3674] } <= { data_i[74:74] };
    end 
    if(N10050) begin
      { mem[3673:3673] } <= { data_i[73:73] };
    end 
    if(N10049) begin
      { mem[3672:3672] } <= { data_i[72:72] };
    end 
    if(N10048) begin
      { mem[3671:3671] } <= { data_i[71:71] };
    end 
    if(N10047) begin
      { mem[3670:3670] } <= { data_i[70:70] };
    end 
    if(N10046) begin
      { mem[3669:3669] } <= { data_i[69:69] };
    end 
    if(N10045) begin
      { mem[3668:3668] } <= { data_i[68:68] };
    end 
    if(N10044) begin
      { mem[3667:3667] } <= { data_i[67:67] };
    end 
    if(N10043) begin
      { mem[3666:3666] } <= { data_i[66:66] };
    end 
    if(N10042) begin
      { mem[3665:3665] } <= { data_i[65:65] };
    end 
    if(N10041) begin
      { mem[3664:3664] } <= { data_i[64:64] };
    end 
    if(N10040) begin
      { mem[3663:3663] } <= { data_i[63:63] };
    end 
    if(N10039) begin
      { mem[3662:3662] } <= { data_i[62:62] };
    end 
    if(N10038) begin
      { mem[3661:3661] } <= { data_i[61:61] };
    end 
    if(N10037) begin
      { mem[3660:3660] } <= { data_i[60:60] };
    end 
    if(N10036) begin
      { mem[3659:3659] } <= { data_i[59:59] };
    end 
    if(N10035) begin
      { mem[3658:3658] } <= { data_i[58:58] };
    end 
    if(N10034) begin
      { mem[3657:3657] } <= { data_i[57:57] };
    end 
    if(N10033) begin
      { mem[3656:3656] } <= { data_i[56:56] };
    end 
    if(N10032) begin
      { mem[3655:3655] } <= { data_i[55:55] };
    end 
    if(N10031) begin
      { mem[3654:3654] } <= { data_i[54:54] };
    end 
    if(N10030) begin
      { mem[3653:3653] } <= { data_i[53:53] };
    end 
    if(N10029) begin
      { mem[3652:3652] } <= { data_i[52:52] };
    end 
    if(N10028) begin
      { mem[3651:3651] } <= { data_i[51:51] };
    end 
    if(N10027) begin
      { mem[3650:3650] } <= { data_i[50:50] };
    end 
    if(N10026) begin
      { mem[3649:3649] } <= { data_i[49:49] };
    end 
    if(N10025) begin
      { mem[3648:3648] } <= { data_i[48:48] };
    end 
    if(N10024) begin
      { mem[3647:3647] } <= { data_i[47:47] };
    end 
    if(N10023) begin
      { mem[3646:3646] } <= { data_i[46:46] };
    end 
    if(N10022) begin
      { mem[3645:3645] } <= { data_i[45:45] };
    end 
    if(N10021) begin
      { mem[3644:3644] } <= { data_i[44:44] };
    end 
    if(N10020) begin
      { mem[3643:3643] } <= { data_i[43:43] };
    end 
    if(N10019) begin
      { mem[3642:3642] } <= { data_i[42:42] };
    end 
    if(N10018) begin
      { mem[3641:3641] } <= { data_i[41:41] };
    end 
    if(N10017) begin
      { mem[3640:3640] } <= { data_i[40:40] };
    end 
    if(N10016) begin
      { mem[3639:3639] } <= { data_i[39:39] };
    end 
    if(N10015) begin
      { mem[3638:3638] } <= { data_i[38:38] };
    end 
    if(N10014) begin
      { mem[3637:3637] } <= { data_i[37:37] };
    end 
    if(N10013) begin
      { mem[3636:3636] } <= { data_i[36:36] };
    end 
    if(N10012) begin
      { mem[3635:3635] } <= { data_i[35:35] };
    end 
    if(N10011) begin
      { mem[3634:3634] } <= { data_i[34:34] };
    end 
    if(N10010) begin
      { mem[3633:3633] } <= { data_i[33:33] };
    end 
    if(N10009) begin
      { mem[3632:3632] } <= { data_i[32:32] };
    end 
    if(N10008) begin
      { mem[3631:3631] } <= { data_i[31:31] };
    end 
    if(N10007) begin
      { mem[3630:3630] } <= { data_i[30:30] };
    end 
    if(N10006) begin
      { mem[3629:3629] } <= { data_i[29:29] };
    end 
    if(N10005) begin
      { mem[3628:3628] } <= { data_i[28:28] };
    end 
    if(N10004) begin
      { mem[3627:3627] } <= { data_i[27:27] };
    end 
    if(N10003) begin
      { mem[3626:3626] } <= { data_i[26:26] };
    end 
    if(N10002) begin
      { mem[3625:3625] } <= { data_i[25:25] };
    end 
    if(N10001) begin
      { mem[3624:3624] } <= { data_i[24:24] };
    end 
    if(N10000) begin
      { mem[3623:3623] } <= { data_i[23:23] };
    end 
    if(N9999) begin
      { mem[3622:3622] } <= { data_i[22:22] };
    end 
    if(N9998) begin
      { mem[3621:3621] } <= { data_i[21:21] };
    end 
    if(N9997) begin
      { mem[3620:3620] } <= { data_i[20:20] };
    end 
    if(N9996) begin
      { mem[3619:3619] } <= { data_i[19:19] };
    end 
    if(N9995) begin
      { mem[3618:3618] } <= { data_i[18:18] };
    end 
    if(N9994) begin
      { mem[3617:3617] } <= { data_i[17:17] };
    end 
    if(N9993) begin
      { mem[3616:3616] } <= { data_i[16:16] };
    end 
    if(N9992) begin
      { mem[3615:3615] } <= { data_i[15:15] };
    end 
    if(N9991) begin
      { mem[3614:3614] } <= { data_i[14:14] };
    end 
    if(N9990) begin
      { mem[3613:3613] } <= { data_i[13:13] };
    end 
    if(N9989) begin
      { mem[3612:3612] } <= { data_i[12:12] };
    end 
    if(N9988) begin
      { mem[3611:3611] } <= { data_i[11:11] };
    end 
    if(N9987) begin
      { mem[3610:3610] } <= { data_i[10:10] };
    end 
    if(N9986) begin
      { mem[3609:3609] } <= { data_i[9:9] };
    end 
    if(N9985) begin
      { mem[3608:3608] } <= { data_i[8:8] };
    end 
    if(N9984) begin
      { mem[3607:3607] } <= { data_i[7:7] };
    end 
    if(N9983) begin
      { mem[3606:3606] } <= { data_i[6:6] };
    end 
    if(N9982) begin
      { mem[3605:3605] } <= { data_i[5:5] };
    end 
    if(N9981) begin
      { mem[3604:3604] } <= { data_i[4:4] };
    end 
    if(N9980) begin
      { mem[3603:3603] } <= { data_i[3:3] };
    end 
    if(N9979) begin
      { mem[3602:3602] } <= { data_i[2:2] };
    end 
    if(N9978) begin
      { mem[3601:3601] } <= { data_i[1:1] };
    end 
    if(N9977) begin
      { mem[3600:3600] } <= { data_i[0:0] };
    end 
    if(N9976) begin
      { mem[3599:3599] } <= { data_i[79:79] };
    end 
    if(N9975) begin
      { mem[3598:3598] } <= { data_i[78:78] };
    end 
    if(N9974) begin
      { mem[3597:3597] } <= { data_i[77:77] };
    end 
    if(N9973) begin
      { mem[3596:3596] } <= { data_i[76:76] };
    end 
    if(N9972) begin
      { mem[3595:3595] } <= { data_i[75:75] };
    end 
    if(N9971) begin
      { mem[3594:3594] } <= { data_i[74:74] };
    end 
    if(N9970) begin
      { mem[3593:3593] } <= { data_i[73:73] };
    end 
    if(N9969) begin
      { mem[3592:3592] } <= { data_i[72:72] };
    end 
    if(N9968) begin
      { mem[3591:3591] } <= { data_i[71:71] };
    end 
    if(N9967) begin
      { mem[3590:3590] } <= { data_i[70:70] };
    end 
    if(N9966) begin
      { mem[3589:3589] } <= { data_i[69:69] };
    end 
    if(N9965) begin
      { mem[3588:3588] } <= { data_i[68:68] };
    end 
    if(N9964) begin
      { mem[3587:3587] } <= { data_i[67:67] };
    end 
    if(N9963) begin
      { mem[3586:3586] } <= { data_i[66:66] };
    end 
    if(N9962) begin
      { mem[3585:3585] } <= { data_i[65:65] };
    end 
    if(N9961) begin
      { mem[3584:3584] } <= { data_i[64:64] };
    end 
    if(N9960) begin
      { mem[3583:3583] } <= { data_i[63:63] };
    end 
    if(N9959) begin
      { mem[3582:3582] } <= { data_i[62:62] };
    end 
    if(N9958) begin
      { mem[3581:3581] } <= { data_i[61:61] };
    end 
    if(N9957) begin
      { mem[3580:3580] } <= { data_i[60:60] };
    end 
    if(N9956) begin
      { mem[3579:3579] } <= { data_i[59:59] };
    end 
    if(N9955) begin
      { mem[3578:3578] } <= { data_i[58:58] };
    end 
    if(N9954) begin
      { mem[3577:3577] } <= { data_i[57:57] };
    end 
    if(N9953) begin
      { mem[3576:3576] } <= { data_i[56:56] };
    end 
    if(N9952) begin
      { mem[3575:3575] } <= { data_i[55:55] };
    end 
    if(N9951) begin
      { mem[3574:3574] } <= { data_i[54:54] };
    end 
    if(N9950) begin
      { mem[3573:3573] } <= { data_i[53:53] };
    end 
    if(N9949) begin
      { mem[3572:3572] } <= { data_i[52:52] };
    end 
    if(N9948) begin
      { mem[3571:3571] } <= { data_i[51:51] };
    end 
    if(N9947) begin
      { mem[3570:3570] } <= { data_i[50:50] };
    end 
    if(N9946) begin
      { mem[3569:3569] } <= { data_i[49:49] };
    end 
    if(N9945) begin
      { mem[3568:3568] } <= { data_i[48:48] };
    end 
    if(N9944) begin
      { mem[3567:3567] } <= { data_i[47:47] };
    end 
    if(N9943) begin
      { mem[3566:3566] } <= { data_i[46:46] };
    end 
    if(N9942) begin
      { mem[3565:3565] } <= { data_i[45:45] };
    end 
    if(N9941) begin
      { mem[3564:3564] } <= { data_i[44:44] };
    end 
    if(N9940) begin
      { mem[3563:3563] } <= { data_i[43:43] };
    end 
    if(N9939) begin
      { mem[3562:3562] } <= { data_i[42:42] };
    end 
    if(N9938) begin
      { mem[3561:3561] } <= { data_i[41:41] };
    end 
    if(N9937) begin
      { mem[3560:3560] } <= { data_i[40:40] };
    end 
    if(N9936) begin
      { mem[3559:3559] } <= { data_i[39:39] };
    end 
    if(N9935) begin
      { mem[3558:3558] } <= { data_i[38:38] };
    end 
    if(N9934) begin
      { mem[3557:3557] } <= { data_i[37:37] };
    end 
    if(N9933) begin
      { mem[3556:3556] } <= { data_i[36:36] };
    end 
    if(N9932) begin
      { mem[3555:3555] } <= { data_i[35:35] };
    end 
    if(N9931) begin
      { mem[3554:3554] } <= { data_i[34:34] };
    end 
    if(N9930) begin
      { mem[3553:3553] } <= { data_i[33:33] };
    end 
    if(N9929) begin
      { mem[3552:3552] } <= { data_i[32:32] };
    end 
    if(N9928) begin
      { mem[3551:3551] } <= { data_i[31:31] };
    end 
    if(N9927) begin
      { mem[3550:3550] } <= { data_i[30:30] };
    end 
    if(N9926) begin
      { mem[3549:3549] } <= { data_i[29:29] };
    end 
    if(N9925) begin
      { mem[3548:3548] } <= { data_i[28:28] };
    end 
    if(N9924) begin
      { mem[3547:3547] } <= { data_i[27:27] };
    end 
    if(N9923) begin
      { mem[3546:3546] } <= { data_i[26:26] };
    end 
    if(N9922) begin
      { mem[3545:3545] } <= { data_i[25:25] };
    end 
    if(N9921) begin
      { mem[3544:3544] } <= { data_i[24:24] };
    end 
    if(N9920) begin
      { mem[3543:3543] } <= { data_i[23:23] };
    end 
    if(N9919) begin
      { mem[3542:3542] } <= { data_i[22:22] };
    end 
    if(N9918) begin
      { mem[3541:3541] } <= { data_i[21:21] };
    end 
    if(N9917) begin
      { mem[3540:3540] } <= { data_i[20:20] };
    end 
    if(N9916) begin
      { mem[3539:3539] } <= { data_i[19:19] };
    end 
    if(N9915) begin
      { mem[3538:3538] } <= { data_i[18:18] };
    end 
    if(N9914) begin
      { mem[3537:3537] } <= { data_i[17:17] };
    end 
    if(N9913) begin
      { mem[3536:3536] } <= { data_i[16:16] };
    end 
    if(N9912) begin
      { mem[3535:3535] } <= { data_i[15:15] };
    end 
    if(N9911) begin
      { mem[3534:3534] } <= { data_i[14:14] };
    end 
    if(N9910) begin
      { mem[3533:3533] } <= { data_i[13:13] };
    end 
    if(N9909) begin
      { mem[3532:3532] } <= { data_i[12:12] };
    end 
    if(N9908) begin
      { mem[3531:3531] } <= { data_i[11:11] };
    end 
    if(N9907) begin
      { mem[3530:3530] } <= { data_i[10:10] };
    end 
    if(N9906) begin
      { mem[3529:3529] } <= { data_i[9:9] };
    end 
    if(N9905) begin
      { mem[3528:3528] } <= { data_i[8:8] };
    end 
    if(N9904) begin
      { mem[3527:3527] } <= { data_i[7:7] };
    end 
    if(N9903) begin
      { mem[3526:3526] } <= { data_i[6:6] };
    end 
    if(N9902) begin
      { mem[3525:3525] } <= { data_i[5:5] };
    end 
    if(N9901) begin
      { mem[3524:3524] } <= { data_i[4:4] };
    end 
    if(N9900) begin
      { mem[3523:3523] } <= { data_i[3:3] };
    end 
    if(N9899) begin
      { mem[3522:3522] } <= { data_i[2:2] };
    end 
    if(N9898) begin
      { mem[3521:3521] } <= { data_i[1:1] };
    end 
    if(N9897) begin
      { mem[3520:3520] } <= { data_i[0:0] };
    end 
    if(N9896) begin
      { mem[3519:3519] } <= { data_i[79:79] };
    end 
    if(N9895) begin
      { mem[3518:3518] } <= { data_i[78:78] };
    end 
    if(N9894) begin
      { mem[3517:3517] } <= { data_i[77:77] };
    end 
    if(N9893) begin
      { mem[3516:3516] } <= { data_i[76:76] };
    end 
    if(N9892) begin
      { mem[3515:3515] } <= { data_i[75:75] };
    end 
    if(N9891) begin
      { mem[3514:3514] } <= { data_i[74:74] };
    end 
    if(N9890) begin
      { mem[3513:3513] } <= { data_i[73:73] };
    end 
    if(N9889) begin
      { mem[3512:3512] } <= { data_i[72:72] };
    end 
    if(N9888) begin
      { mem[3511:3511] } <= { data_i[71:71] };
    end 
    if(N9887) begin
      { mem[3510:3510] } <= { data_i[70:70] };
    end 
    if(N9886) begin
      { mem[3509:3509] } <= { data_i[69:69] };
    end 
    if(N9885) begin
      { mem[3508:3508] } <= { data_i[68:68] };
    end 
    if(N9884) begin
      { mem[3507:3507] } <= { data_i[67:67] };
    end 
    if(N9883) begin
      { mem[3506:3506] } <= { data_i[66:66] };
    end 
    if(N9882) begin
      { mem[3505:3505] } <= { data_i[65:65] };
    end 
    if(N9881) begin
      { mem[3504:3504] } <= { data_i[64:64] };
    end 
    if(N9880) begin
      { mem[3503:3503] } <= { data_i[63:63] };
    end 
    if(N9879) begin
      { mem[3502:3502] } <= { data_i[62:62] };
    end 
    if(N9878) begin
      { mem[3501:3501] } <= { data_i[61:61] };
    end 
    if(N9877) begin
      { mem[3500:3500] } <= { data_i[60:60] };
    end 
    if(N9876) begin
      { mem[3499:3499] } <= { data_i[59:59] };
    end 
    if(N9875) begin
      { mem[3498:3498] } <= { data_i[58:58] };
    end 
    if(N9874) begin
      { mem[3497:3497] } <= { data_i[57:57] };
    end 
    if(N9873) begin
      { mem[3496:3496] } <= { data_i[56:56] };
    end 
    if(N9872) begin
      { mem[3495:3495] } <= { data_i[55:55] };
    end 
    if(N9871) begin
      { mem[3494:3494] } <= { data_i[54:54] };
    end 
    if(N9870) begin
      { mem[3493:3493] } <= { data_i[53:53] };
    end 
    if(N9869) begin
      { mem[3492:3492] } <= { data_i[52:52] };
    end 
    if(N9868) begin
      { mem[3491:3491] } <= { data_i[51:51] };
    end 
    if(N9867) begin
      { mem[3490:3490] } <= { data_i[50:50] };
    end 
    if(N9866) begin
      { mem[3489:3489] } <= { data_i[49:49] };
    end 
    if(N9865) begin
      { mem[3488:3488] } <= { data_i[48:48] };
    end 
    if(N9864) begin
      { mem[3487:3487] } <= { data_i[47:47] };
    end 
    if(N9863) begin
      { mem[3486:3486] } <= { data_i[46:46] };
    end 
    if(N9862) begin
      { mem[3485:3485] } <= { data_i[45:45] };
    end 
    if(N9861) begin
      { mem[3484:3484] } <= { data_i[44:44] };
    end 
    if(N9860) begin
      { mem[3483:3483] } <= { data_i[43:43] };
    end 
    if(N9859) begin
      { mem[3482:3482] } <= { data_i[42:42] };
    end 
    if(N9858) begin
      { mem[3481:3481] } <= { data_i[41:41] };
    end 
    if(N9857) begin
      { mem[3480:3480] } <= { data_i[40:40] };
    end 
    if(N9856) begin
      { mem[3479:3479] } <= { data_i[39:39] };
    end 
    if(N9855) begin
      { mem[3478:3478] } <= { data_i[38:38] };
    end 
    if(N9854) begin
      { mem[3477:3477] } <= { data_i[37:37] };
    end 
    if(N9853) begin
      { mem[3476:3476] } <= { data_i[36:36] };
    end 
    if(N9852) begin
      { mem[3475:3475] } <= { data_i[35:35] };
    end 
    if(N9851) begin
      { mem[3474:3474] } <= { data_i[34:34] };
    end 
    if(N9850) begin
      { mem[3473:3473] } <= { data_i[33:33] };
    end 
    if(N9849) begin
      { mem[3472:3472] } <= { data_i[32:32] };
    end 
    if(N9848) begin
      { mem[3471:3471] } <= { data_i[31:31] };
    end 
    if(N9847) begin
      { mem[3470:3470] } <= { data_i[30:30] };
    end 
    if(N9846) begin
      { mem[3469:3469] } <= { data_i[29:29] };
    end 
    if(N9845) begin
      { mem[3468:3468] } <= { data_i[28:28] };
    end 
    if(N9844) begin
      { mem[3467:3467] } <= { data_i[27:27] };
    end 
    if(N9843) begin
      { mem[3466:3466] } <= { data_i[26:26] };
    end 
    if(N9842) begin
      { mem[3465:3465] } <= { data_i[25:25] };
    end 
    if(N9841) begin
      { mem[3464:3464] } <= { data_i[24:24] };
    end 
    if(N9840) begin
      { mem[3463:3463] } <= { data_i[23:23] };
    end 
    if(N9839) begin
      { mem[3462:3462] } <= { data_i[22:22] };
    end 
    if(N9838) begin
      { mem[3461:3461] } <= { data_i[21:21] };
    end 
    if(N9837) begin
      { mem[3460:3460] } <= { data_i[20:20] };
    end 
    if(N9836) begin
      { mem[3459:3459] } <= { data_i[19:19] };
    end 
    if(N9835) begin
      { mem[3458:3458] } <= { data_i[18:18] };
    end 
    if(N9834) begin
      { mem[3457:3457] } <= { data_i[17:17] };
    end 
    if(N9833) begin
      { mem[3456:3456] } <= { data_i[16:16] };
    end 
    if(N9832) begin
      { mem[3455:3455] } <= { data_i[15:15] };
    end 
    if(N9831) begin
      { mem[3454:3454] } <= { data_i[14:14] };
    end 
    if(N9830) begin
      { mem[3453:3453] } <= { data_i[13:13] };
    end 
    if(N9829) begin
      { mem[3452:3452] } <= { data_i[12:12] };
    end 
    if(N9828) begin
      { mem[3451:3451] } <= { data_i[11:11] };
    end 
    if(N9827) begin
      { mem[3450:3450] } <= { data_i[10:10] };
    end 
    if(N9826) begin
      { mem[3449:3449] } <= { data_i[9:9] };
    end 
    if(N9825) begin
      { mem[3448:3448] } <= { data_i[8:8] };
    end 
    if(N9824) begin
      { mem[3447:3447] } <= { data_i[7:7] };
    end 
    if(N9823) begin
      { mem[3446:3446] } <= { data_i[6:6] };
    end 
    if(N9822) begin
      { mem[3445:3445] } <= { data_i[5:5] };
    end 
    if(N9821) begin
      { mem[3444:3444] } <= { data_i[4:4] };
    end 
    if(N9820) begin
      { mem[3443:3443] } <= { data_i[3:3] };
    end 
    if(N9819) begin
      { mem[3442:3442] } <= { data_i[2:2] };
    end 
    if(N9818) begin
      { mem[3441:3441] } <= { data_i[1:1] };
    end 
    if(N9817) begin
      { mem[3440:3440] } <= { data_i[0:0] };
    end 
    if(N9816) begin
      { mem[3439:3439] } <= { data_i[79:79] };
    end 
    if(N9815) begin
      { mem[3438:3438] } <= { data_i[78:78] };
    end 
    if(N9814) begin
      { mem[3437:3437] } <= { data_i[77:77] };
    end 
    if(N9813) begin
      { mem[3436:3436] } <= { data_i[76:76] };
    end 
    if(N9812) begin
      { mem[3435:3435] } <= { data_i[75:75] };
    end 
    if(N9811) begin
      { mem[3434:3434] } <= { data_i[74:74] };
    end 
    if(N9810) begin
      { mem[3433:3433] } <= { data_i[73:73] };
    end 
    if(N9809) begin
      { mem[3432:3432] } <= { data_i[72:72] };
    end 
    if(N9808) begin
      { mem[3431:3431] } <= { data_i[71:71] };
    end 
    if(N9807) begin
      { mem[3430:3430] } <= { data_i[70:70] };
    end 
    if(N9806) begin
      { mem[3429:3429] } <= { data_i[69:69] };
    end 
    if(N9805) begin
      { mem[3428:3428] } <= { data_i[68:68] };
    end 
    if(N9804) begin
      { mem[3427:3427] } <= { data_i[67:67] };
    end 
    if(N9803) begin
      { mem[3426:3426] } <= { data_i[66:66] };
    end 
    if(N9802) begin
      { mem[3425:3425] } <= { data_i[65:65] };
    end 
    if(N9801) begin
      { mem[3424:3424] } <= { data_i[64:64] };
    end 
    if(N9800) begin
      { mem[3423:3423] } <= { data_i[63:63] };
    end 
    if(N9799) begin
      { mem[3422:3422] } <= { data_i[62:62] };
    end 
    if(N9798) begin
      { mem[3421:3421] } <= { data_i[61:61] };
    end 
    if(N9797) begin
      { mem[3420:3420] } <= { data_i[60:60] };
    end 
    if(N9796) begin
      { mem[3419:3419] } <= { data_i[59:59] };
    end 
    if(N9795) begin
      { mem[3418:3418] } <= { data_i[58:58] };
    end 
    if(N9794) begin
      { mem[3417:3417] } <= { data_i[57:57] };
    end 
    if(N9793) begin
      { mem[3416:3416] } <= { data_i[56:56] };
    end 
    if(N9792) begin
      { mem[3415:3415] } <= { data_i[55:55] };
    end 
    if(N9791) begin
      { mem[3414:3414] } <= { data_i[54:54] };
    end 
    if(N9790) begin
      { mem[3413:3413] } <= { data_i[53:53] };
    end 
    if(N9789) begin
      { mem[3412:3412] } <= { data_i[52:52] };
    end 
    if(N9788) begin
      { mem[3411:3411] } <= { data_i[51:51] };
    end 
    if(N9787) begin
      { mem[3410:3410] } <= { data_i[50:50] };
    end 
    if(N9786) begin
      { mem[3409:3409] } <= { data_i[49:49] };
    end 
    if(N9785) begin
      { mem[3408:3408] } <= { data_i[48:48] };
    end 
    if(N9784) begin
      { mem[3407:3407] } <= { data_i[47:47] };
    end 
    if(N9783) begin
      { mem[3406:3406] } <= { data_i[46:46] };
    end 
    if(N9782) begin
      { mem[3405:3405] } <= { data_i[45:45] };
    end 
    if(N9781) begin
      { mem[3404:3404] } <= { data_i[44:44] };
    end 
    if(N9780) begin
      { mem[3403:3403] } <= { data_i[43:43] };
    end 
    if(N9779) begin
      { mem[3402:3402] } <= { data_i[42:42] };
    end 
    if(N9778) begin
      { mem[3401:3401] } <= { data_i[41:41] };
    end 
    if(N9777) begin
      { mem[3400:3400] } <= { data_i[40:40] };
    end 
    if(N9776) begin
      { mem[3399:3399] } <= { data_i[39:39] };
    end 
    if(N9775) begin
      { mem[3398:3398] } <= { data_i[38:38] };
    end 
    if(N9774) begin
      { mem[3397:3397] } <= { data_i[37:37] };
    end 
    if(N9773) begin
      { mem[3396:3396] } <= { data_i[36:36] };
    end 
    if(N9772) begin
      { mem[3395:3395] } <= { data_i[35:35] };
    end 
    if(N9771) begin
      { mem[3394:3394] } <= { data_i[34:34] };
    end 
    if(N9770) begin
      { mem[3393:3393] } <= { data_i[33:33] };
    end 
    if(N9769) begin
      { mem[3392:3392] } <= { data_i[32:32] };
    end 
    if(N9768) begin
      { mem[3391:3391] } <= { data_i[31:31] };
    end 
    if(N9767) begin
      { mem[3390:3390] } <= { data_i[30:30] };
    end 
    if(N9766) begin
      { mem[3389:3389] } <= { data_i[29:29] };
    end 
    if(N9765) begin
      { mem[3388:3388] } <= { data_i[28:28] };
    end 
    if(N9764) begin
      { mem[3387:3387] } <= { data_i[27:27] };
    end 
    if(N9763) begin
      { mem[3386:3386] } <= { data_i[26:26] };
    end 
    if(N9762) begin
      { mem[3385:3385] } <= { data_i[25:25] };
    end 
    if(N9761) begin
      { mem[3384:3384] } <= { data_i[24:24] };
    end 
    if(N9760) begin
      { mem[3383:3383] } <= { data_i[23:23] };
    end 
    if(N9759) begin
      { mem[3382:3382] } <= { data_i[22:22] };
    end 
    if(N9758) begin
      { mem[3381:3381] } <= { data_i[21:21] };
    end 
    if(N9757) begin
      { mem[3380:3380] } <= { data_i[20:20] };
    end 
    if(N9756) begin
      { mem[3379:3379] } <= { data_i[19:19] };
    end 
    if(N9755) begin
      { mem[3378:3378] } <= { data_i[18:18] };
    end 
    if(N9754) begin
      { mem[3377:3377] } <= { data_i[17:17] };
    end 
    if(N9753) begin
      { mem[3376:3376] } <= { data_i[16:16] };
    end 
    if(N9752) begin
      { mem[3375:3375] } <= { data_i[15:15] };
    end 
    if(N9751) begin
      { mem[3374:3374] } <= { data_i[14:14] };
    end 
    if(N9750) begin
      { mem[3373:3373] } <= { data_i[13:13] };
    end 
    if(N9749) begin
      { mem[3372:3372] } <= { data_i[12:12] };
    end 
    if(N9748) begin
      { mem[3371:3371] } <= { data_i[11:11] };
    end 
    if(N9747) begin
      { mem[3370:3370] } <= { data_i[10:10] };
    end 
    if(N9746) begin
      { mem[3369:3369] } <= { data_i[9:9] };
    end 
    if(N9745) begin
      { mem[3368:3368] } <= { data_i[8:8] };
    end 
    if(N9744) begin
      { mem[3367:3367] } <= { data_i[7:7] };
    end 
    if(N9743) begin
      { mem[3366:3366] } <= { data_i[6:6] };
    end 
    if(N9742) begin
      { mem[3365:3365] } <= { data_i[5:5] };
    end 
    if(N9741) begin
      { mem[3364:3364] } <= { data_i[4:4] };
    end 
    if(N9740) begin
      { mem[3363:3363] } <= { data_i[3:3] };
    end 
    if(N9739) begin
      { mem[3362:3362] } <= { data_i[2:2] };
    end 
    if(N9738) begin
      { mem[3361:3361] } <= { data_i[1:1] };
    end 
    if(N9737) begin
      { mem[3360:3360] } <= { data_i[0:0] };
    end 
    if(N9736) begin
      { mem[3359:3359] } <= { data_i[79:79] };
    end 
    if(N9735) begin
      { mem[3358:3358] } <= { data_i[78:78] };
    end 
    if(N9734) begin
      { mem[3357:3357] } <= { data_i[77:77] };
    end 
    if(N9733) begin
      { mem[3356:3356] } <= { data_i[76:76] };
    end 
    if(N9732) begin
      { mem[3355:3355] } <= { data_i[75:75] };
    end 
    if(N9731) begin
      { mem[3354:3354] } <= { data_i[74:74] };
    end 
    if(N9730) begin
      { mem[3353:3353] } <= { data_i[73:73] };
    end 
    if(N9729) begin
      { mem[3352:3352] } <= { data_i[72:72] };
    end 
    if(N9728) begin
      { mem[3351:3351] } <= { data_i[71:71] };
    end 
    if(N9727) begin
      { mem[3350:3350] } <= { data_i[70:70] };
    end 
    if(N9726) begin
      { mem[3349:3349] } <= { data_i[69:69] };
    end 
    if(N9725) begin
      { mem[3348:3348] } <= { data_i[68:68] };
    end 
    if(N9724) begin
      { mem[3347:3347] } <= { data_i[67:67] };
    end 
    if(N9723) begin
      { mem[3346:3346] } <= { data_i[66:66] };
    end 
    if(N9722) begin
      { mem[3345:3345] } <= { data_i[65:65] };
    end 
    if(N9721) begin
      { mem[3344:3344] } <= { data_i[64:64] };
    end 
    if(N9720) begin
      { mem[3343:3343] } <= { data_i[63:63] };
    end 
    if(N9719) begin
      { mem[3342:3342] } <= { data_i[62:62] };
    end 
    if(N9718) begin
      { mem[3341:3341] } <= { data_i[61:61] };
    end 
    if(N9717) begin
      { mem[3340:3340] } <= { data_i[60:60] };
    end 
    if(N9716) begin
      { mem[3339:3339] } <= { data_i[59:59] };
    end 
    if(N9715) begin
      { mem[3338:3338] } <= { data_i[58:58] };
    end 
    if(N9714) begin
      { mem[3337:3337] } <= { data_i[57:57] };
    end 
    if(N9713) begin
      { mem[3336:3336] } <= { data_i[56:56] };
    end 
    if(N9712) begin
      { mem[3335:3335] } <= { data_i[55:55] };
    end 
    if(N9711) begin
      { mem[3334:3334] } <= { data_i[54:54] };
    end 
    if(N9710) begin
      { mem[3333:3333] } <= { data_i[53:53] };
    end 
    if(N9709) begin
      { mem[3332:3332] } <= { data_i[52:52] };
    end 
    if(N9708) begin
      { mem[3331:3331] } <= { data_i[51:51] };
    end 
    if(N9707) begin
      { mem[3330:3330] } <= { data_i[50:50] };
    end 
    if(N9706) begin
      { mem[3329:3329] } <= { data_i[49:49] };
    end 
    if(N9705) begin
      { mem[3328:3328] } <= { data_i[48:48] };
    end 
    if(N9704) begin
      { mem[3327:3327] } <= { data_i[47:47] };
    end 
    if(N9703) begin
      { mem[3326:3326] } <= { data_i[46:46] };
    end 
    if(N9702) begin
      { mem[3325:3325] } <= { data_i[45:45] };
    end 
    if(N9701) begin
      { mem[3324:3324] } <= { data_i[44:44] };
    end 
    if(N9700) begin
      { mem[3323:3323] } <= { data_i[43:43] };
    end 
    if(N9699) begin
      { mem[3322:3322] } <= { data_i[42:42] };
    end 
    if(N9698) begin
      { mem[3321:3321] } <= { data_i[41:41] };
    end 
    if(N9697) begin
      { mem[3320:3320] } <= { data_i[40:40] };
    end 
    if(N9696) begin
      { mem[3319:3319] } <= { data_i[39:39] };
    end 
    if(N9695) begin
      { mem[3318:3318] } <= { data_i[38:38] };
    end 
    if(N9694) begin
      { mem[3317:3317] } <= { data_i[37:37] };
    end 
    if(N9693) begin
      { mem[3316:3316] } <= { data_i[36:36] };
    end 
    if(N9692) begin
      { mem[3315:3315] } <= { data_i[35:35] };
    end 
    if(N9691) begin
      { mem[3314:3314] } <= { data_i[34:34] };
    end 
    if(N9690) begin
      { mem[3313:3313] } <= { data_i[33:33] };
    end 
    if(N9689) begin
      { mem[3312:3312] } <= { data_i[32:32] };
    end 
    if(N9688) begin
      { mem[3311:3311] } <= { data_i[31:31] };
    end 
    if(N9687) begin
      { mem[3310:3310] } <= { data_i[30:30] };
    end 
    if(N9686) begin
      { mem[3309:3309] } <= { data_i[29:29] };
    end 
    if(N9685) begin
      { mem[3308:3308] } <= { data_i[28:28] };
    end 
    if(N9684) begin
      { mem[3307:3307] } <= { data_i[27:27] };
    end 
    if(N9683) begin
      { mem[3306:3306] } <= { data_i[26:26] };
    end 
    if(N9682) begin
      { mem[3305:3305] } <= { data_i[25:25] };
    end 
    if(N9681) begin
      { mem[3304:3304] } <= { data_i[24:24] };
    end 
    if(N9680) begin
      { mem[3303:3303] } <= { data_i[23:23] };
    end 
    if(N9679) begin
      { mem[3302:3302] } <= { data_i[22:22] };
    end 
    if(N9678) begin
      { mem[3301:3301] } <= { data_i[21:21] };
    end 
    if(N9677) begin
      { mem[3300:3300] } <= { data_i[20:20] };
    end 
    if(N9676) begin
      { mem[3299:3299] } <= { data_i[19:19] };
    end 
    if(N9675) begin
      { mem[3298:3298] } <= { data_i[18:18] };
    end 
    if(N9674) begin
      { mem[3297:3297] } <= { data_i[17:17] };
    end 
    if(N9673) begin
      { mem[3296:3296] } <= { data_i[16:16] };
    end 
    if(N9672) begin
      { mem[3295:3295] } <= { data_i[15:15] };
    end 
    if(N9671) begin
      { mem[3294:3294] } <= { data_i[14:14] };
    end 
    if(N9670) begin
      { mem[3293:3293] } <= { data_i[13:13] };
    end 
    if(N9669) begin
      { mem[3292:3292] } <= { data_i[12:12] };
    end 
    if(N9668) begin
      { mem[3291:3291] } <= { data_i[11:11] };
    end 
    if(N9667) begin
      { mem[3290:3290] } <= { data_i[10:10] };
    end 
    if(N9666) begin
      { mem[3289:3289] } <= { data_i[9:9] };
    end 
    if(N9665) begin
      { mem[3288:3288] } <= { data_i[8:8] };
    end 
    if(N9664) begin
      { mem[3287:3287] } <= { data_i[7:7] };
    end 
    if(N9663) begin
      { mem[3286:3286] } <= { data_i[6:6] };
    end 
    if(N9662) begin
      { mem[3285:3285] } <= { data_i[5:5] };
    end 
    if(N9661) begin
      { mem[3284:3284] } <= { data_i[4:4] };
    end 
    if(N9660) begin
      { mem[3283:3283] } <= { data_i[3:3] };
    end 
    if(N9659) begin
      { mem[3282:3282] } <= { data_i[2:2] };
    end 
    if(N9658) begin
      { mem[3281:3281] } <= { data_i[1:1] };
    end 
    if(N9657) begin
      { mem[3280:3280] } <= { data_i[0:0] };
    end 
    if(N9656) begin
      { mem[3279:3279] } <= { data_i[79:79] };
    end 
    if(N9655) begin
      { mem[3278:3278] } <= { data_i[78:78] };
    end 
    if(N9654) begin
      { mem[3277:3277] } <= { data_i[77:77] };
    end 
    if(N9653) begin
      { mem[3276:3276] } <= { data_i[76:76] };
    end 
    if(N9652) begin
      { mem[3275:3275] } <= { data_i[75:75] };
    end 
    if(N9651) begin
      { mem[3274:3274] } <= { data_i[74:74] };
    end 
    if(N9650) begin
      { mem[3273:3273] } <= { data_i[73:73] };
    end 
    if(N9649) begin
      { mem[3272:3272] } <= { data_i[72:72] };
    end 
    if(N9648) begin
      { mem[3271:3271] } <= { data_i[71:71] };
    end 
    if(N9647) begin
      { mem[3270:3270] } <= { data_i[70:70] };
    end 
    if(N9646) begin
      { mem[3269:3269] } <= { data_i[69:69] };
    end 
    if(N9645) begin
      { mem[3268:3268] } <= { data_i[68:68] };
    end 
    if(N9644) begin
      { mem[3267:3267] } <= { data_i[67:67] };
    end 
    if(N9643) begin
      { mem[3266:3266] } <= { data_i[66:66] };
    end 
    if(N9642) begin
      { mem[3265:3265] } <= { data_i[65:65] };
    end 
    if(N9641) begin
      { mem[3264:3264] } <= { data_i[64:64] };
    end 
    if(N9640) begin
      { mem[3263:3263] } <= { data_i[63:63] };
    end 
    if(N9639) begin
      { mem[3262:3262] } <= { data_i[62:62] };
    end 
    if(N9638) begin
      { mem[3261:3261] } <= { data_i[61:61] };
    end 
    if(N9637) begin
      { mem[3260:3260] } <= { data_i[60:60] };
    end 
    if(N9636) begin
      { mem[3259:3259] } <= { data_i[59:59] };
    end 
    if(N9635) begin
      { mem[3258:3258] } <= { data_i[58:58] };
    end 
    if(N9634) begin
      { mem[3257:3257] } <= { data_i[57:57] };
    end 
    if(N9633) begin
      { mem[3256:3256] } <= { data_i[56:56] };
    end 
    if(N9632) begin
      { mem[3255:3255] } <= { data_i[55:55] };
    end 
    if(N9631) begin
      { mem[3254:3254] } <= { data_i[54:54] };
    end 
    if(N9630) begin
      { mem[3253:3253] } <= { data_i[53:53] };
    end 
    if(N9629) begin
      { mem[3252:3252] } <= { data_i[52:52] };
    end 
    if(N9628) begin
      { mem[3251:3251] } <= { data_i[51:51] };
    end 
    if(N9627) begin
      { mem[3250:3250] } <= { data_i[50:50] };
    end 
    if(N9626) begin
      { mem[3249:3249] } <= { data_i[49:49] };
    end 
    if(N9625) begin
      { mem[3248:3248] } <= { data_i[48:48] };
    end 
    if(N9624) begin
      { mem[3247:3247] } <= { data_i[47:47] };
    end 
    if(N9623) begin
      { mem[3246:3246] } <= { data_i[46:46] };
    end 
    if(N9622) begin
      { mem[3245:3245] } <= { data_i[45:45] };
    end 
    if(N9621) begin
      { mem[3244:3244] } <= { data_i[44:44] };
    end 
    if(N9620) begin
      { mem[3243:3243] } <= { data_i[43:43] };
    end 
    if(N9619) begin
      { mem[3242:3242] } <= { data_i[42:42] };
    end 
    if(N9618) begin
      { mem[3241:3241] } <= { data_i[41:41] };
    end 
    if(N9617) begin
      { mem[3240:3240] } <= { data_i[40:40] };
    end 
    if(N9616) begin
      { mem[3239:3239] } <= { data_i[39:39] };
    end 
    if(N9615) begin
      { mem[3238:3238] } <= { data_i[38:38] };
    end 
    if(N9614) begin
      { mem[3237:3237] } <= { data_i[37:37] };
    end 
    if(N9613) begin
      { mem[3236:3236] } <= { data_i[36:36] };
    end 
    if(N9612) begin
      { mem[3235:3235] } <= { data_i[35:35] };
    end 
    if(N9611) begin
      { mem[3234:3234] } <= { data_i[34:34] };
    end 
    if(N9610) begin
      { mem[3233:3233] } <= { data_i[33:33] };
    end 
    if(N9609) begin
      { mem[3232:3232] } <= { data_i[32:32] };
    end 
    if(N9608) begin
      { mem[3231:3231] } <= { data_i[31:31] };
    end 
    if(N9607) begin
      { mem[3230:3230] } <= { data_i[30:30] };
    end 
    if(N9606) begin
      { mem[3229:3229] } <= { data_i[29:29] };
    end 
    if(N9605) begin
      { mem[3228:3228] } <= { data_i[28:28] };
    end 
    if(N9604) begin
      { mem[3227:3227] } <= { data_i[27:27] };
    end 
    if(N9603) begin
      { mem[3226:3226] } <= { data_i[26:26] };
    end 
    if(N9602) begin
      { mem[3225:3225] } <= { data_i[25:25] };
    end 
    if(N9601) begin
      { mem[3224:3224] } <= { data_i[24:24] };
    end 
    if(N9600) begin
      { mem[3223:3223] } <= { data_i[23:23] };
    end 
    if(N9599) begin
      { mem[3222:3222] } <= { data_i[22:22] };
    end 
    if(N9598) begin
      { mem[3221:3221] } <= { data_i[21:21] };
    end 
    if(N9597) begin
      { mem[3220:3220] } <= { data_i[20:20] };
    end 
    if(N9596) begin
      { mem[3219:3219] } <= { data_i[19:19] };
    end 
    if(N9595) begin
      { mem[3218:3218] } <= { data_i[18:18] };
    end 
    if(N9594) begin
      { mem[3217:3217] } <= { data_i[17:17] };
    end 
    if(N9593) begin
      { mem[3216:3216] } <= { data_i[16:16] };
    end 
    if(N9592) begin
      { mem[3215:3215] } <= { data_i[15:15] };
    end 
    if(N9591) begin
      { mem[3214:3214] } <= { data_i[14:14] };
    end 
    if(N9590) begin
      { mem[3213:3213] } <= { data_i[13:13] };
    end 
    if(N9589) begin
      { mem[3212:3212] } <= { data_i[12:12] };
    end 
    if(N9588) begin
      { mem[3211:3211] } <= { data_i[11:11] };
    end 
    if(N9587) begin
      { mem[3210:3210] } <= { data_i[10:10] };
    end 
    if(N9586) begin
      { mem[3209:3209] } <= { data_i[9:9] };
    end 
    if(N9585) begin
      { mem[3208:3208] } <= { data_i[8:8] };
    end 
    if(N9584) begin
      { mem[3207:3207] } <= { data_i[7:7] };
    end 
    if(N9583) begin
      { mem[3206:3206] } <= { data_i[6:6] };
    end 
    if(N9582) begin
      { mem[3205:3205] } <= { data_i[5:5] };
    end 
    if(N9581) begin
      { mem[3204:3204] } <= { data_i[4:4] };
    end 
    if(N9580) begin
      { mem[3203:3203] } <= { data_i[3:3] };
    end 
    if(N9579) begin
      { mem[3202:3202] } <= { data_i[2:2] };
    end 
    if(N9578) begin
      { mem[3201:3201] } <= { data_i[1:1] };
    end 
    if(N9577) begin
      { mem[3200:3200] } <= { data_i[0:0] };
    end 
    if(N9576) begin
      { mem[3199:3199] } <= { data_i[79:79] };
    end 
    if(N9575) begin
      { mem[3198:3198] } <= { data_i[78:78] };
    end 
    if(N9574) begin
      { mem[3197:3197] } <= { data_i[77:77] };
    end 
    if(N9573) begin
      { mem[3196:3196] } <= { data_i[76:76] };
    end 
    if(N9572) begin
      { mem[3195:3195] } <= { data_i[75:75] };
    end 
    if(N9571) begin
      { mem[3194:3194] } <= { data_i[74:74] };
    end 
    if(N9570) begin
      { mem[3193:3193] } <= { data_i[73:73] };
    end 
    if(N9569) begin
      { mem[3192:3192] } <= { data_i[72:72] };
    end 
    if(N9568) begin
      { mem[3191:3191] } <= { data_i[71:71] };
    end 
    if(N9567) begin
      { mem[3190:3190] } <= { data_i[70:70] };
    end 
    if(N9566) begin
      { mem[3189:3189] } <= { data_i[69:69] };
    end 
    if(N9565) begin
      { mem[3188:3188] } <= { data_i[68:68] };
    end 
    if(N9564) begin
      { mem[3187:3187] } <= { data_i[67:67] };
    end 
    if(N9563) begin
      { mem[3186:3186] } <= { data_i[66:66] };
    end 
    if(N9562) begin
      { mem[3185:3185] } <= { data_i[65:65] };
    end 
    if(N9561) begin
      { mem[3184:3184] } <= { data_i[64:64] };
    end 
    if(N9560) begin
      { mem[3183:3183] } <= { data_i[63:63] };
    end 
    if(N9559) begin
      { mem[3182:3182] } <= { data_i[62:62] };
    end 
    if(N9558) begin
      { mem[3181:3181] } <= { data_i[61:61] };
    end 
    if(N9557) begin
      { mem[3180:3180] } <= { data_i[60:60] };
    end 
    if(N9556) begin
      { mem[3179:3179] } <= { data_i[59:59] };
    end 
    if(N9555) begin
      { mem[3178:3178] } <= { data_i[58:58] };
    end 
    if(N9554) begin
      { mem[3177:3177] } <= { data_i[57:57] };
    end 
    if(N9553) begin
      { mem[3176:3176] } <= { data_i[56:56] };
    end 
    if(N9552) begin
      { mem[3175:3175] } <= { data_i[55:55] };
    end 
    if(N9551) begin
      { mem[3174:3174] } <= { data_i[54:54] };
    end 
    if(N9550) begin
      { mem[3173:3173] } <= { data_i[53:53] };
    end 
    if(N9549) begin
      { mem[3172:3172] } <= { data_i[52:52] };
    end 
    if(N9548) begin
      { mem[3171:3171] } <= { data_i[51:51] };
    end 
    if(N9547) begin
      { mem[3170:3170] } <= { data_i[50:50] };
    end 
    if(N9546) begin
      { mem[3169:3169] } <= { data_i[49:49] };
    end 
    if(N9545) begin
      { mem[3168:3168] } <= { data_i[48:48] };
    end 
    if(N9544) begin
      { mem[3167:3167] } <= { data_i[47:47] };
    end 
    if(N9543) begin
      { mem[3166:3166] } <= { data_i[46:46] };
    end 
    if(N9542) begin
      { mem[3165:3165] } <= { data_i[45:45] };
    end 
    if(N9541) begin
      { mem[3164:3164] } <= { data_i[44:44] };
    end 
    if(N9540) begin
      { mem[3163:3163] } <= { data_i[43:43] };
    end 
    if(N9539) begin
      { mem[3162:3162] } <= { data_i[42:42] };
    end 
    if(N9538) begin
      { mem[3161:3161] } <= { data_i[41:41] };
    end 
    if(N9537) begin
      { mem[3160:3160] } <= { data_i[40:40] };
    end 
    if(N9536) begin
      { mem[3159:3159] } <= { data_i[39:39] };
    end 
    if(N9535) begin
      { mem[3158:3158] } <= { data_i[38:38] };
    end 
    if(N9534) begin
      { mem[3157:3157] } <= { data_i[37:37] };
    end 
    if(N9533) begin
      { mem[3156:3156] } <= { data_i[36:36] };
    end 
    if(N9532) begin
      { mem[3155:3155] } <= { data_i[35:35] };
    end 
    if(N9531) begin
      { mem[3154:3154] } <= { data_i[34:34] };
    end 
    if(N9530) begin
      { mem[3153:3153] } <= { data_i[33:33] };
    end 
    if(N9529) begin
      { mem[3152:3152] } <= { data_i[32:32] };
    end 
    if(N9528) begin
      { mem[3151:3151] } <= { data_i[31:31] };
    end 
    if(N9527) begin
      { mem[3150:3150] } <= { data_i[30:30] };
    end 
    if(N9526) begin
      { mem[3149:3149] } <= { data_i[29:29] };
    end 
    if(N9525) begin
      { mem[3148:3148] } <= { data_i[28:28] };
    end 
    if(N9524) begin
      { mem[3147:3147] } <= { data_i[27:27] };
    end 
    if(N9523) begin
      { mem[3146:3146] } <= { data_i[26:26] };
    end 
    if(N9522) begin
      { mem[3145:3145] } <= { data_i[25:25] };
    end 
    if(N9521) begin
      { mem[3144:3144] } <= { data_i[24:24] };
    end 
    if(N9520) begin
      { mem[3143:3143] } <= { data_i[23:23] };
    end 
    if(N9519) begin
      { mem[3142:3142] } <= { data_i[22:22] };
    end 
    if(N9518) begin
      { mem[3141:3141] } <= { data_i[21:21] };
    end 
    if(N9517) begin
      { mem[3140:3140] } <= { data_i[20:20] };
    end 
    if(N9516) begin
      { mem[3139:3139] } <= { data_i[19:19] };
    end 
    if(N9515) begin
      { mem[3138:3138] } <= { data_i[18:18] };
    end 
    if(N9514) begin
      { mem[3137:3137] } <= { data_i[17:17] };
    end 
    if(N9513) begin
      { mem[3136:3136] } <= { data_i[16:16] };
    end 
    if(N9512) begin
      { mem[3135:3135] } <= { data_i[15:15] };
    end 
    if(N9511) begin
      { mem[3134:3134] } <= { data_i[14:14] };
    end 
    if(N9510) begin
      { mem[3133:3133] } <= { data_i[13:13] };
    end 
    if(N9509) begin
      { mem[3132:3132] } <= { data_i[12:12] };
    end 
    if(N9508) begin
      { mem[3131:3131] } <= { data_i[11:11] };
    end 
    if(N9507) begin
      { mem[3130:3130] } <= { data_i[10:10] };
    end 
    if(N9506) begin
      { mem[3129:3129] } <= { data_i[9:9] };
    end 
    if(N9505) begin
      { mem[3128:3128] } <= { data_i[8:8] };
    end 
    if(N9504) begin
      { mem[3127:3127] } <= { data_i[7:7] };
    end 
    if(N9503) begin
      { mem[3126:3126] } <= { data_i[6:6] };
    end 
    if(N9502) begin
      { mem[3125:3125] } <= { data_i[5:5] };
    end 
    if(N9501) begin
      { mem[3124:3124] } <= { data_i[4:4] };
    end 
    if(N9500) begin
      { mem[3123:3123] } <= { data_i[3:3] };
    end 
    if(N9499) begin
      { mem[3122:3122] } <= { data_i[2:2] };
    end 
    if(N9498) begin
      { mem[3121:3121] } <= { data_i[1:1] };
    end 
    if(N9497) begin
      { mem[3120:3120] } <= { data_i[0:0] };
    end 
    if(N9496) begin
      { mem[3119:3119] } <= { data_i[79:79] };
    end 
    if(N9495) begin
      { mem[3118:3118] } <= { data_i[78:78] };
    end 
    if(N9494) begin
      { mem[3117:3117] } <= { data_i[77:77] };
    end 
    if(N9493) begin
      { mem[3116:3116] } <= { data_i[76:76] };
    end 
    if(N9492) begin
      { mem[3115:3115] } <= { data_i[75:75] };
    end 
    if(N9491) begin
      { mem[3114:3114] } <= { data_i[74:74] };
    end 
    if(N9490) begin
      { mem[3113:3113] } <= { data_i[73:73] };
    end 
    if(N9489) begin
      { mem[3112:3112] } <= { data_i[72:72] };
    end 
    if(N9488) begin
      { mem[3111:3111] } <= { data_i[71:71] };
    end 
    if(N9487) begin
      { mem[3110:3110] } <= { data_i[70:70] };
    end 
    if(N9486) begin
      { mem[3109:3109] } <= { data_i[69:69] };
    end 
    if(N9485) begin
      { mem[3108:3108] } <= { data_i[68:68] };
    end 
    if(N9484) begin
      { mem[3107:3107] } <= { data_i[67:67] };
    end 
    if(N9483) begin
      { mem[3106:3106] } <= { data_i[66:66] };
    end 
    if(N9482) begin
      { mem[3105:3105] } <= { data_i[65:65] };
    end 
    if(N9481) begin
      { mem[3104:3104] } <= { data_i[64:64] };
    end 
    if(N9480) begin
      { mem[3103:3103] } <= { data_i[63:63] };
    end 
    if(N9479) begin
      { mem[3102:3102] } <= { data_i[62:62] };
    end 
    if(N9478) begin
      { mem[3101:3101] } <= { data_i[61:61] };
    end 
    if(N9477) begin
      { mem[3100:3100] } <= { data_i[60:60] };
    end 
    if(N9476) begin
      { mem[3099:3099] } <= { data_i[59:59] };
    end 
    if(N9475) begin
      { mem[3098:3098] } <= { data_i[58:58] };
    end 
    if(N9474) begin
      { mem[3097:3097] } <= { data_i[57:57] };
    end 
    if(N9473) begin
      { mem[3096:3096] } <= { data_i[56:56] };
    end 
    if(N9472) begin
      { mem[3095:3095] } <= { data_i[55:55] };
    end 
    if(N9471) begin
      { mem[3094:3094] } <= { data_i[54:54] };
    end 
    if(N9470) begin
      { mem[3093:3093] } <= { data_i[53:53] };
    end 
    if(N9469) begin
      { mem[3092:3092] } <= { data_i[52:52] };
    end 
    if(N9468) begin
      { mem[3091:3091] } <= { data_i[51:51] };
    end 
    if(N9467) begin
      { mem[3090:3090] } <= { data_i[50:50] };
    end 
    if(N9466) begin
      { mem[3089:3089] } <= { data_i[49:49] };
    end 
    if(N9465) begin
      { mem[3088:3088] } <= { data_i[48:48] };
    end 
    if(N9464) begin
      { mem[3087:3087] } <= { data_i[47:47] };
    end 
    if(N9463) begin
      { mem[3086:3086] } <= { data_i[46:46] };
    end 
    if(N9462) begin
      { mem[3085:3085] } <= { data_i[45:45] };
    end 
    if(N9461) begin
      { mem[3084:3084] } <= { data_i[44:44] };
    end 
    if(N9460) begin
      { mem[3083:3083] } <= { data_i[43:43] };
    end 
    if(N9459) begin
      { mem[3082:3082] } <= { data_i[42:42] };
    end 
    if(N9458) begin
      { mem[3081:3081] } <= { data_i[41:41] };
    end 
    if(N9457) begin
      { mem[3080:3080] } <= { data_i[40:40] };
    end 
    if(N9456) begin
      { mem[3079:3079] } <= { data_i[39:39] };
    end 
    if(N9455) begin
      { mem[3078:3078] } <= { data_i[38:38] };
    end 
    if(N9454) begin
      { mem[3077:3077] } <= { data_i[37:37] };
    end 
    if(N9453) begin
      { mem[3076:3076] } <= { data_i[36:36] };
    end 
    if(N9452) begin
      { mem[3075:3075] } <= { data_i[35:35] };
    end 
    if(N9451) begin
      { mem[3074:3074] } <= { data_i[34:34] };
    end 
    if(N9450) begin
      { mem[3073:3073] } <= { data_i[33:33] };
    end 
    if(N9449) begin
      { mem[3072:3072] } <= { data_i[32:32] };
    end 
    if(N9448) begin
      { mem[3071:3071] } <= { data_i[31:31] };
    end 
    if(N9447) begin
      { mem[3070:3070] } <= { data_i[30:30] };
    end 
    if(N9446) begin
      { mem[3069:3069] } <= { data_i[29:29] };
    end 
    if(N9445) begin
      { mem[3068:3068] } <= { data_i[28:28] };
    end 
    if(N9444) begin
      { mem[3067:3067] } <= { data_i[27:27] };
    end 
    if(N9443) begin
      { mem[3066:3066] } <= { data_i[26:26] };
    end 
    if(N9442) begin
      { mem[3065:3065] } <= { data_i[25:25] };
    end 
    if(N9441) begin
      { mem[3064:3064] } <= { data_i[24:24] };
    end 
    if(N9440) begin
      { mem[3063:3063] } <= { data_i[23:23] };
    end 
    if(N9439) begin
      { mem[3062:3062] } <= { data_i[22:22] };
    end 
    if(N9438) begin
      { mem[3061:3061] } <= { data_i[21:21] };
    end 
    if(N9437) begin
      { mem[3060:3060] } <= { data_i[20:20] };
    end 
    if(N9436) begin
      { mem[3059:3059] } <= { data_i[19:19] };
    end 
    if(N9435) begin
      { mem[3058:3058] } <= { data_i[18:18] };
    end 
    if(N9434) begin
      { mem[3057:3057] } <= { data_i[17:17] };
    end 
    if(N9433) begin
      { mem[3056:3056] } <= { data_i[16:16] };
    end 
    if(N9432) begin
      { mem[3055:3055] } <= { data_i[15:15] };
    end 
    if(N9431) begin
      { mem[3054:3054] } <= { data_i[14:14] };
    end 
    if(N9430) begin
      { mem[3053:3053] } <= { data_i[13:13] };
    end 
    if(N9429) begin
      { mem[3052:3052] } <= { data_i[12:12] };
    end 
    if(N9428) begin
      { mem[3051:3051] } <= { data_i[11:11] };
    end 
    if(N9427) begin
      { mem[3050:3050] } <= { data_i[10:10] };
    end 
    if(N9426) begin
      { mem[3049:3049] } <= { data_i[9:9] };
    end 
    if(N9425) begin
      { mem[3048:3048] } <= { data_i[8:8] };
    end 
    if(N9424) begin
      { mem[3047:3047] } <= { data_i[7:7] };
    end 
    if(N9423) begin
      { mem[3046:3046] } <= { data_i[6:6] };
    end 
    if(N9422) begin
      { mem[3045:3045] } <= { data_i[5:5] };
    end 
    if(N9421) begin
      { mem[3044:3044] } <= { data_i[4:4] };
    end 
    if(N9420) begin
      { mem[3043:3043] } <= { data_i[3:3] };
    end 
    if(N9419) begin
      { mem[3042:3042] } <= { data_i[2:2] };
    end 
    if(N9418) begin
      { mem[3041:3041] } <= { data_i[1:1] };
    end 
    if(N9417) begin
      { mem[3040:3040] } <= { data_i[0:0] };
    end 
    if(N9416) begin
      { mem[3039:3039] } <= { data_i[79:79] };
    end 
    if(N9415) begin
      { mem[3038:3038] } <= { data_i[78:78] };
    end 
    if(N9414) begin
      { mem[3037:3037] } <= { data_i[77:77] };
    end 
    if(N9413) begin
      { mem[3036:3036] } <= { data_i[76:76] };
    end 
    if(N9412) begin
      { mem[3035:3035] } <= { data_i[75:75] };
    end 
    if(N9411) begin
      { mem[3034:3034] } <= { data_i[74:74] };
    end 
    if(N9410) begin
      { mem[3033:3033] } <= { data_i[73:73] };
    end 
    if(N9409) begin
      { mem[3032:3032] } <= { data_i[72:72] };
    end 
    if(N9408) begin
      { mem[3031:3031] } <= { data_i[71:71] };
    end 
    if(N9407) begin
      { mem[3030:3030] } <= { data_i[70:70] };
    end 
    if(N9406) begin
      { mem[3029:3029] } <= { data_i[69:69] };
    end 
    if(N9405) begin
      { mem[3028:3028] } <= { data_i[68:68] };
    end 
    if(N9404) begin
      { mem[3027:3027] } <= { data_i[67:67] };
    end 
    if(N9403) begin
      { mem[3026:3026] } <= { data_i[66:66] };
    end 
    if(N9402) begin
      { mem[3025:3025] } <= { data_i[65:65] };
    end 
    if(N9401) begin
      { mem[3024:3024] } <= { data_i[64:64] };
    end 
    if(N9400) begin
      { mem[3023:3023] } <= { data_i[63:63] };
    end 
    if(N9399) begin
      { mem[3022:3022] } <= { data_i[62:62] };
    end 
    if(N9398) begin
      { mem[3021:3021] } <= { data_i[61:61] };
    end 
    if(N9397) begin
      { mem[3020:3020] } <= { data_i[60:60] };
    end 
    if(N9396) begin
      { mem[3019:3019] } <= { data_i[59:59] };
    end 
    if(N9395) begin
      { mem[3018:3018] } <= { data_i[58:58] };
    end 
    if(N9394) begin
      { mem[3017:3017] } <= { data_i[57:57] };
    end 
    if(N9393) begin
      { mem[3016:3016] } <= { data_i[56:56] };
    end 
    if(N9392) begin
      { mem[3015:3015] } <= { data_i[55:55] };
    end 
    if(N9391) begin
      { mem[3014:3014] } <= { data_i[54:54] };
    end 
    if(N9390) begin
      { mem[3013:3013] } <= { data_i[53:53] };
    end 
    if(N9389) begin
      { mem[3012:3012] } <= { data_i[52:52] };
    end 
    if(N9388) begin
      { mem[3011:3011] } <= { data_i[51:51] };
    end 
    if(N9387) begin
      { mem[3010:3010] } <= { data_i[50:50] };
    end 
    if(N9386) begin
      { mem[3009:3009] } <= { data_i[49:49] };
    end 
    if(N9385) begin
      { mem[3008:3008] } <= { data_i[48:48] };
    end 
    if(N9384) begin
      { mem[3007:3007] } <= { data_i[47:47] };
    end 
    if(N9383) begin
      { mem[3006:3006] } <= { data_i[46:46] };
    end 
    if(N9382) begin
      { mem[3005:3005] } <= { data_i[45:45] };
    end 
    if(N9381) begin
      { mem[3004:3004] } <= { data_i[44:44] };
    end 
    if(N9380) begin
      { mem[3003:3003] } <= { data_i[43:43] };
    end 
    if(N9379) begin
      { mem[3002:3002] } <= { data_i[42:42] };
    end 
    if(N9378) begin
      { mem[3001:3001] } <= { data_i[41:41] };
    end 
    if(N9377) begin
      { mem[3000:3000] } <= { data_i[40:40] };
    end 
    if(N9376) begin
      { mem[2999:2999] } <= { data_i[39:39] };
    end 
    if(N9375) begin
      { mem[2998:2998] } <= { data_i[38:38] };
    end 
    if(N9374) begin
      { mem[2997:2997] } <= { data_i[37:37] };
    end 
    if(N9373) begin
      { mem[2996:2996] } <= { data_i[36:36] };
    end 
    if(N9372) begin
      { mem[2995:2995] } <= { data_i[35:35] };
    end 
    if(N9371) begin
      { mem[2994:2994] } <= { data_i[34:34] };
    end 
    if(N9370) begin
      { mem[2993:2993] } <= { data_i[33:33] };
    end 
    if(N9369) begin
      { mem[2992:2992] } <= { data_i[32:32] };
    end 
    if(N9368) begin
      { mem[2991:2991] } <= { data_i[31:31] };
    end 
    if(N9367) begin
      { mem[2990:2990] } <= { data_i[30:30] };
    end 
    if(N9366) begin
      { mem[2989:2989] } <= { data_i[29:29] };
    end 
    if(N9365) begin
      { mem[2988:2988] } <= { data_i[28:28] };
    end 
    if(N9364) begin
      { mem[2987:2987] } <= { data_i[27:27] };
    end 
    if(N9363) begin
      { mem[2986:2986] } <= { data_i[26:26] };
    end 
    if(N9362) begin
      { mem[2985:2985] } <= { data_i[25:25] };
    end 
    if(N9361) begin
      { mem[2984:2984] } <= { data_i[24:24] };
    end 
    if(N9360) begin
      { mem[2983:2983] } <= { data_i[23:23] };
    end 
    if(N9359) begin
      { mem[2982:2982] } <= { data_i[22:22] };
    end 
    if(N9358) begin
      { mem[2981:2981] } <= { data_i[21:21] };
    end 
    if(N9357) begin
      { mem[2980:2980] } <= { data_i[20:20] };
    end 
    if(N9356) begin
      { mem[2979:2979] } <= { data_i[19:19] };
    end 
    if(N9355) begin
      { mem[2978:2978] } <= { data_i[18:18] };
    end 
    if(N9354) begin
      { mem[2977:2977] } <= { data_i[17:17] };
    end 
    if(N9353) begin
      { mem[2976:2976] } <= { data_i[16:16] };
    end 
    if(N9352) begin
      { mem[2975:2975] } <= { data_i[15:15] };
    end 
    if(N9351) begin
      { mem[2974:2974] } <= { data_i[14:14] };
    end 
    if(N9350) begin
      { mem[2973:2973] } <= { data_i[13:13] };
    end 
    if(N9349) begin
      { mem[2972:2972] } <= { data_i[12:12] };
    end 
    if(N9348) begin
      { mem[2971:2971] } <= { data_i[11:11] };
    end 
    if(N9347) begin
      { mem[2970:2970] } <= { data_i[10:10] };
    end 
    if(N9346) begin
      { mem[2969:2969] } <= { data_i[9:9] };
    end 
    if(N9345) begin
      { mem[2968:2968] } <= { data_i[8:8] };
    end 
    if(N9344) begin
      { mem[2967:2967] } <= { data_i[7:7] };
    end 
    if(N9343) begin
      { mem[2966:2966] } <= { data_i[6:6] };
    end 
    if(N9342) begin
      { mem[2965:2965] } <= { data_i[5:5] };
    end 
    if(N9341) begin
      { mem[2964:2964] } <= { data_i[4:4] };
    end 
    if(N9340) begin
      { mem[2963:2963] } <= { data_i[3:3] };
    end 
    if(N9339) begin
      { mem[2962:2962] } <= { data_i[2:2] };
    end 
    if(N9338) begin
      { mem[2961:2961] } <= { data_i[1:1] };
    end 
    if(N9337) begin
      { mem[2960:2960] } <= { data_i[0:0] };
    end 
    if(N9336) begin
      { mem[2959:2959] } <= { data_i[79:79] };
    end 
    if(N9335) begin
      { mem[2958:2958] } <= { data_i[78:78] };
    end 
    if(N9334) begin
      { mem[2957:2957] } <= { data_i[77:77] };
    end 
    if(N9333) begin
      { mem[2956:2956] } <= { data_i[76:76] };
    end 
    if(N9332) begin
      { mem[2955:2955] } <= { data_i[75:75] };
    end 
    if(N9331) begin
      { mem[2954:2954] } <= { data_i[74:74] };
    end 
    if(N9330) begin
      { mem[2953:2953] } <= { data_i[73:73] };
    end 
    if(N9329) begin
      { mem[2952:2952] } <= { data_i[72:72] };
    end 
    if(N9328) begin
      { mem[2951:2951] } <= { data_i[71:71] };
    end 
    if(N9327) begin
      { mem[2950:2950] } <= { data_i[70:70] };
    end 
    if(N9326) begin
      { mem[2949:2949] } <= { data_i[69:69] };
    end 
    if(N9325) begin
      { mem[2948:2948] } <= { data_i[68:68] };
    end 
    if(N9324) begin
      { mem[2947:2947] } <= { data_i[67:67] };
    end 
    if(N9323) begin
      { mem[2946:2946] } <= { data_i[66:66] };
    end 
    if(N9322) begin
      { mem[2945:2945] } <= { data_i[65:65] };
    end 
    if(N9321) begin
      { mem[2944:2944] } <= { data_i[64:64] };
    end 
    if(N9320) begin
      { mem[2943:2943] } <= { data_i[63:63] };
    end 
    if(N9319) begin
      { mem[2942:2942] } <= { data_i[62:62] };
    end 
    if(N9318) begin
      { mem[2941:2941] } <= { data_i[61:61] };
    end 
    if(N9317) begin
      { mem[2940:2940] } <= { data_i[60:60] };
    end 
    if(N9316) begin
      { mem[2939:2939] } <= { data_i[59:59] };
    end 
    if(N9315) begin
      { mem[2938:2938] } <= { data_i[58:58] };
    end 
    if(N9314) begin
      { mem[2937:2937] } <= { data_i[57:57] };
    end 
    if(N9313) begin
      { mem[2936:2936] } <= { data_i[56:56] };
    end 
    if(N9312) begin
      { mem[2935:2935] } <= { data_i[55:55] };
    end 
    if(N9311) begin
      { mem[2934:2934] } <= { data_i[54:54] };
    end 
    if(N9310) begin
      { mem[2933:2933] } <= { data_i[53:53] };
    end 
    if(N9309) begin
      { mem[2932:2932] } <= { data_i[52:52] };
    end 
    if(N9308) begin
      { mem[2931:2931] } <= { data_i[51:51] };
    end 
    if(N9307) begin
      { mem[2930:2930] } <= { data_i[50:50] };
    end 
    if(N9306) begin
      { mem[2929:2929] } <= { data_i[49:49] };
    end 
    if(N9305) begin
      { mem[2928:2928] } <= { data_i[48:48] };
    end 
    if(N9304) begin
      { mem[2927:2927] } <= { data_i[47:47] };
    end 
    if(N9303) begin
      { mem[2926:2926] } <= { data_i[46:46] };
    end 
    if(N9302) begin
      { mem[2925:2925] } <= { data_i[45:45] };
    end 
    if(N9301) begin
      { mem[2924:2924] } <= { data_i[44:44] };
    end 
    if(N9300) begin
      { mem[2923:2923] } <= { data_i[43:43] };
    end 
    if(N9299) begin
      { mem[2922:2922] } <= { data_i[42:42] };
    end 
    if(N9298) begin
      { mem[2921:2921] } <= { data_i[41:41] };
    end 
    if(N9297) begin
      { mem[2920:2920] } <= { data_i[40:40] };
    end 
    if(N9296) begin
      { mem[2919:2919] } <= { data_i[39:39] };
    end 
    if(N9295) begin
      { mem[2918:2918] } <= { data_i[38:38] };
    end 
    if(N9294) begin
      { mem[2917:2917] } <= { data_i[37:37] };
    end 
    if(N9293) begin
      { mem[2916:2916] } <= { data_i[36:36] };
    end 
    if(N9292) begin
      { mem[2915:2915] } <= { data_i[35:35] };
    end 
    if(N9291) begin
      { mem[2914:2914] } <= { data_i[34:34] };
    end 
    if(N9290) begin
      { mem[2913:2913] } <= { data_i[33:33] };
    end 
    if(N9289) begin
      { mem[2912:2912] } <= { data_i[32:32] };
    end 
    if(N9288) begin
      { mem[2911:2911] } <= { data_i[31:31] };
    end 
    if(N9287) begin
      { mem[2910:2910] } <= { data_i[30:30] };
    end 
    if(N9286) begin
      { mem[2909:2909] } <= { data_i[29:29] };
    end 
    if(N9285) begin
      { mem[2908:2908] } <= { data_i[28:28] };
    end 
    if(N9284) begin
      { mem[2907:2907] } <= { data_i[27:27] };
    end 
    if(N9283) begin
      { mem[2906:2906] } <= { data_i[26:26] };
    end 
    if(N9282) begin
      { mem[2905:2905] } <= { data_i[25:25] };
    end 
    if(N9281) begin
      { mem[2904:2904] } <= { data_i[24:24] };
    end 
    if(N9280) begin
      { mem[2903:2903] } <= { data_i[23:23] };
    end 
    if(N9279) begin
      { mem[2902:2902] } <= { data_i[22:22] };
    end 
    if(N9278) begin
      { mem[2901:2901] } <= { data_i[21:21] };
    end 
    if(N9277) begin
      { mem[2900:2900] } <= { data_i[20:20] };
    end 
    if(N9276) begin
      { mem[2899:2899] } <= { data_i[19:19] };
    end 
    if(N9275) begin
      { mem[2898:2898] } <= { data_i[18:18] };
    end 
    if(N9274) begin
      { mem[2897:2897] } <= { data_i[17:17] };
    end 
    if(N9273) begin
      { mem[2896:2896] } <= { data_i[16:16] };
    end 
    if(N9272) begin
      { mem[2895:2895] } <= { data_i[15:15] };
    end 
    if(N9271) begin
      { mem[2894:2894] } <= { data_i[14:14] };
    end 
    if(N9270) begin
      { mem[2893:2893] } <= { data_i[13:13] };
    end 
    if(N9269) begin
      { mem[2892:2892] } <= { data_i[12:12] };
    end 
    if(N9268) begin
      { mem[2891:2891] } <= { data_i[11:11] };
    end 
    if(N9267) begin
      { mem[2890:2890] } <= { data_i[10:10] };
    end 
    if(N9266) begin
      { mem[2889:2889] } <= { data_i[9:9] };
    end 
    if(N9265) begin
      { mem[2888:2888] } <= { data_i[8:8] };
    end 
    if(N9264) begin
      { mem[2887:2887] } <= { data_i[7:7] };
    end 
    if(N9263) begin
      { mem[2886:2886] } <= { data_i[6:6] };
    end 
    if(N9262) begin
      { mem[2885:2885] } <= { data_i[5:5] };
    end 
    if(N9261) begin
      { mem[2884:2884] } <= { data_i[4:4] };
    end 
    if(N9260) begin
      { mem[2883:2883] } <= { data_i[3:3] };
    end 
    if(N9259) begin
      { mem[2882:2882] } <= { data_i[2:2] };
    end 
    if(N9258) begin
      { mem[2881:2881] } <= { data_i[1:1] };
    end 
    if(N9257) begin
      { mem[2880:2880] } <= { data_i[0:0] };
    end 
    if(N9256) begin
      { mem[2879:2879] } <= { data_i[79:79] };
    end 
    if(N9255) begin
      { mem[2878:2878] } <= { data_i[78:78] };
    end 
    if(N9254) begin
      { mem[2877:2877] } <= { data_i[77:77] };
    end 
    if(N9253) begin
      { mem[2876:2876] } <= { data_i[76:76] };
    end 
    if(N9252) begin
      { mem[2875:2875] } <= { data_i[75:75] };
    end 
    if(N9251) begin
      { mem[2874:2874] } <= { data_i[74:74] };
    end 
    if(N9250) begin
      { mem[2873:2873] } <= { data_i[73:73] };
    end 
    if(N9249) begin
      { mem[2872:2872] } <= { data_i[72:72] };
    end 
    if(N9248) begin
      { mem[2871:2871] } <= { data_i[71:71] };
    end 
    if(N9247) begin
      { mem[2870:2870] } <= { data_i[70:70] };
    end 
    if(N9246) begin
      { mem[2869:2869] } <= { data_i[69:69] };
    end 
    if(N9245) begin
      { mem[2868:2868] } <= { data_i[68:68] };
    end 
    if(N9244) begin
      { mem[2867:2867] } <= { data_i[67:67] };
    end 
    if(N9243) begin
      { mem[2866:2866] } <= { data_i[66:66] };
    end 
    if(N9242) begin
      { mem[2865:2865] } <= { data_i[65:65] };
    end 
    if(N9241) begin
      { mem[2864:2864] } <= { data_i[64:64] };
    end 
    if(N9240) begin
      { mem[2863:2863] } <= { data_i[63:63] };
    end 
    if(N9239) begin
      { mem[2862:2862] } <= { data_i[62:62] };
    end 
    if(N9238) begin
      { mem[2861:2861] } <= { data_i[61:61] };
    end 
    if(N9237) begin
      { mem[2860:2860] } <= { data_i[60:60] };
    end 
    if(N9236) begin
      { mem[2859:2859] } <= { data_i[59:59] };
    end 
    if(N9235) begin
      { mem[2858:2858] } <= { data_i[58:58] };
    end 
    if(N9234) begin
      { mem[2857:2857] } <= { data_i[57:57] };
    end 
    if(N9233) begin
      { mem[2856:2856] } <= { data_i[56:56] };
    end 
    if(N9232) begin
      { mem[2855:2855] } <= { data_i[55:55] };
    end 
    if(N9231) begin
      { mem[2854:2854] } <= { data_i[54:54] };
    end 
    if(N9230) begin
      { mem[2853:2853] } <= { data_i[53:53] };
    end 
    if(N9229) begin
      { mem[2852:2852] } <= { data_i[52:52] };
    end 
    if(N9228) begin
      { mem[2851:2851] } <= { data_i[51:51] };
    end 
    if(N9227) begin
      { mem[2850:2850] } <= { data_i[50:50] };
    end 
    if(N9226) begin
      { mem[2849:2849] } <= { data_i[49:49] };
    end 
    if(N9225) begin
      { mem[2848:2848] } <= { data_i[48:48] };
    end 
    if(N9224) begin
      { mem[2847:2847] } <= { data_i[47:47] };
    end 
    if(N9223) begin
      { mem[2846:2846] } <= { data_i[46:46] };
    end 
    if(N9222) begin
      { mem[2845:2845] } <= { data_i[45:45] };
    end 
    if(N9221) begin
      { mem[2844:2844] } <= { data_i[44:44] };
    end 
    if(N9220) begin
      { mem[2843:2843] } <= { data_i[43:43] };
    end 
    if(N9219) begin
      { mem[2842:2842] } <= { data_i[42:42] };
    end 
    if(N9218) begin
      { mem[2841:2841] } <= { data_i[41:41] };
    end 
    if(N9217) begin
      { mem[2840:2840] } <= { data_i[40:40] };
    end 
    if(N9216) begin
      { mem[2839:2839] } <= { data_i[39:39] };
    end 
    if(N9215) begin
      { mem[2838:2838] } <= { data_i[38:38] };
    end 
    if(N9214) begin
      { mem[2837:2837] } <= { data_i[37:37] };
    end 
    if(N9213) begin
      { mem[2836:2836] } <= { data_i[36:36] };
    end 
    if(N9212) begin
      { mem[2835:2835] } <= { data_i[35:35] };
    end 
    if(N9211) begin
      { mem[2834:2834] } <= { data_i[34:34] };
    end 
    if(N9210) begin
      { mem[2833:2833] } <= { data_i[33:33] };
    end 
    if(N9209) begin
      { mem[2832:2832] } <= { data_i[32:32] };
    end 
    if(N9208) begin
      { mem[2831:2831] } <= { data_i[31:31] };
    end 
    if(N9207) begin
      { mem[2830:2830] } <= { data_i[30:30] };
    end 
    if(N9206) begin
      { mem[2829:2829] } <= { data_i[29:29] };
    end 
    if(N9205) begin
      { mem[2828:2828] } <= { data_i[28:28] };
    end 
    if(N9204) begin
      { mem[2827:2827] } <= { data_i[27:27] };
    end 
    if(N9203) begin
      { mem[2826:2826] } <= { data_i[26:26] };
    end 
    if(N9202) begin
      { mem[2825:2825] } <= { data_i[25:25] };
    end 
    if(N9201) begin
      { mem[2824:2824] } <= { data_i[24:24] };
    end 
    if(N9200) begin
      { mem[2823:2823] } <= { data_i[23:23] };
    end 
    if(N9199) begin
      { mem[2822:2822] } <= { data_i[22:22] };
    end 
    if(N9198) begin
      { mem[2821:2821] } <= { data_i[21:21] };
    end 
    if(N9197) begin
      { mem[2820:2820] } <= { data_i[20:20] };
    end 
    if(N9196) begin
      { mem[2819:2819] } <= { data_i[19:19] };
    end 
    if(N9195) begin
      { mem[2818:2818] } <= { data_i[18:18] };
    end 
    if(N9194) begin
      { mem[2817:2817] } <= { data_i[17:17] };
    end 
    if(N9193) begin
      { mem[2816:2816] } <= { data_i[16:16] };
    end 
    if(N9192) begin
      { mem[2815:2815] } <= { data_i[15:15] };
    end 
    if(N9191) begin
      { mem[2814:2814] } <= { data_i[14:14] };
    end 
    if(N9190) begin
      { mem[2813:2813] } <= { data_i[13:13] };
    end 
    if(N9189) begin
      { mem[2812:2812] } <= { data_i[12:12] };
    end 
    if(N9188) begin
      { mem[2811:2811] } <= { data_i[11:11] };
    end 
    if(N9187) begin
      { mem[2810:2810] } <= { data_i[10:10] };
    end 
    if(N9186) begin
      { mem[2809:2809] } <= { data_i[9:9] };
    end 
    if(N9185) begin
      { mem[2808:2808] } <= { data_i[8:8] };
    end 
    if(N9184) begin
      { mem[2807:2807] } <= { data_i[7:7] };
    end 
    if(N9183) begin
      { mem[2806:2806] } <= { data_i[6:6] };
    end 
    if(N9182) begin
      { mem[2805:2805] } <= { data_i[5:5] };
    end 
    if(N9181) begin
      { mem[2804:2804] } <= { data_i[4:4] };
    end 
    if(N9180) begin
      { mem[2803:2803] } <= { data_i[3:3] };
    end 
    if(N9179) begin
      { mem[2802:2802] } <= { data_i[2:2] };
    end 
    if(N9178) begin
      { mem[2801:2801] } <= { data_i[1:1] };
    end 
    if(N9177) begin
      { mem[2800:2800] } <= { data_i[0:0] };
    end 
    if(N9176) begin
      { mem[2799:2799] } <= { data_i[79:79] };
    end 
    if(N9175) begin
      { mem[2798:2798] } <= { data_i[78:78] };
    end 
    if(N9174) begin
      { mem[2797:2797] } <= { data_i[77:77] };
    end 
    if(N9173) begin
      { mem[2796:2796] } <= { data_i[76:76] };
    end 
    if(N9172) begin
      { mem[2795:2795] } <= { data_i[75:75] };
    end 
    if(N9171) begin
      { mem[2794:2794] } <= { data_i[74:74] };
    end 
    if(N9170) begin
      { mem[2793:2793] } <= { data_i[73:73] };
    end 
    if(N9169) begin
      { mem[2792:2792] } <= { data_i[72:72] };
    end 
    if(N9168) begin
      { mem[2791:2791] } <= { data_i[71:71] };
    end 
    if(N9167) begin
      { mem[2790:2790] } <= { data_i[70:70] };
    end 
    if(N9166) begin
      { mem[2789:2789] } <= { data_i[69:69] };
    end 
    if(N9165) begin
      { mem[2788:2788] } <= { data_i[68:68] };
    end 
    if(N9164) begin
      { mem[2787:2787] } <= { data_i[67:67] };
    end 
    if(N9163) begin
      { mem[2786:2786] } <= { data_i[66:66] };
    end 
    if(N9162) begin
      { mem[2785:2785] } <= { data_i[65:65] };
    end 
    if(N9161) begin
      { mem[2784:2784] } <= { data_i[64:64] };
    end 
    if(N9160) begin
      { mem[2783:2783] } <= { data_i[63:63] };
    end 
    if(N9159) begin
      { mem[2782:2782] } <= { data_i[62:62] };
    end 
    if(N9158) begin
      { mem[2781:2781] } <= { data_i[61:61] };
    end 
    if(N9157) begin
      { mem[2780:2780] } <= { data_i[60:60] };
    end 
    if(N9156) begin
      { mem[2779:2779] } <= { data_i[59:59] };
    end 
    if(N9155) begin
      { mem[2778:2778] } <= { data_i[58:58] };
    end 
    if(N9154) begin
      { mem[2777:2777] } <= { data_i[57:57] };
    end 
    if(N9153) begin
      { mem[2776:2776] } <= { data_i[56:56] };
    end 
    if(N9152) begin
      { mem[2775:2775] } <= { data_i[55:55] };
    end 
    if(N9151) begin
      { mem[2774:2774] } <= { data_i[54:54] };
    end 
    if(N9150) begin
      { mem[2773:2773] } <= { data_i[53:53] };
    end 
    if(N9149) begin
      { mem[2772:2772] } <= { data_i[52:52] };
    end 
    if(N9148) begin
      { mem[2771:2771] } <= { data_i[51:51] };
    end 
    if(N9147) begin
      { mem[2770:2770] } <= { data_i[50:50] };
    end 
    if(N9146) begin
      { mem[2769:2769] } <= { data_i[49:49] };
    end 
    if(N9145) begin
      { mem[2768:2768] } <= { data_i[48:48] };
    end 
    if(N9144) begin
      { mem[2767:2767] } <= { data_i[47:47] };
    end 
    if(N9143) begin
      { mem[2766:2766] } <= { data_i[46:46] };
    end 
    if(N9142) begin
      { mem[2765:2765] } <= { data_i[45:45] };
    end 
    if(N9141) begin
      { mem[2764:2764] } <= { data_i[44:44] };
    end 
    if(N9140) begin
      { mem[2763:2763] } <= { data_i[43:43] };
    end 
    if(N9139) begin
      { mem[2762:2762] } <= { data_i[42:42] };
    end 
    if(N9138) begin
      { mem[2761:2761] } <= { data_i[41:41] };
    end 
    if(N9137) begin
      { mem[2760:2760] } <= { data_i[40:40] };
    end 
    if(N9136) begin
      { mem[2759:2759] } <= { data_i[39:39] };
    end 
    if(N9135) begin
      { mem[2758:2758] } <= { data_i[38:38] };
    end 
    if(N9134) begin
      { mem[2757:2757] } <= { data_i[37:37] };
    end 
    if(N9133) begin
      { mem[2756:2756] } <= { data_i[36:36] };
    end 
    if(N9132) begin
      { mem[2755:2755] } <= { data_i[35:35] };
    end 
    if(N9131) begin
      { mem[2754:2754] } <= { data_i[34:34] };
    end 
    if(N9130) begin
      { mem[2753:2753] } <= { data_i[33:33] };
    end 
    if(N9129) begin
      { mem[2752:2752] } <= { data_i[32:32] };
    end 
    if(N9128) begin
      { mem[2751:2751] } <= { data_i[31:31] };
    end 
    if(N9127) begin
      { mem[2750:2750] } <= { data_i[30:30] };
    end 
    if(N9126) begin
      { mem[2749:2749] } <= { data_i[29:29] };
    end 
    if(N9125) begin
      { mem[2748:2748] } <= { data_i[28:28] };
    end 
    if(N9124) begin
      { mem[2747:2747] } <= { data_i[27:27] };
    end 
    if(N9123) begin
      { mem[2746:2746] } <= { data_i[26:26] };
    end 
    if(N9122) begin
      { mem[2745:2745] } <= { data_i[25:25] };
    end 
    if(N9121) begin
      { mem[2744:2744] } <= { data_i[24:24] };
    end 
    if(N9120) begin
      { mem[2743:2743] } <= { data_i[23:23] };
    end 
    if(N9119) begin
      { mem[2742:2742] } <= { data_i[22:22] };
    end 
    if(N9118) begin
      { mem[2741:2741] } <= { data_i[21:21] };
    end 
    if(N9117) begin
      { mem[2740:2740] } <= { data_i[20:20] };
    end 
    if(N9116) begin
      { mem[2739:2739] } <= { data_i[19:19] };
    end 
    if(N9115) begin
      { mem[2738:2738] } <= { data_i[18:18] };
    end 
    if(N9114) begin
      { mem[2737:2737] } <= { data_i[17:17] };
    end 
    if(N9113) begin
      { mem[2736:2736] } <= { data_i[16:16] };
    end 
    if(N9112) begin
      { mem[2735:2735] } <= { data_i[15:15] };
    end 
    if(N9111) begin
      { mem[2734:2734] } <= { data_i[14:14] };
    end 
    if(N9110) begin
      { mem[2733:2733] } <= { data_i[13:13] };
    end 
    if(N9109) begin
      { mem[2732:2732] } <= { data_i[12:12] };
    end 
    if(N9108) begin
      { mem[2731:2731] } <= { data_i[11:11] };
    end 
    if(N9107) begin
      { mem[2730:2730] } <= { data_i[10:10] };
    end 
    if(N9106) begin
      { mem[2729:2729] } <= { data_i[9:9] };
    end 
    if(N9105) begin
      { mem[2728:2728] } <= { data_i[8:8] };
    end 
    if(N9104) begin
      { mem[2727:2727] } <= { data_i[7:7] };
    end 
    if(N9103) begin
      { mem[2726:2726] } <= { data_i[6:6] };
    end 
    if(N9102) begin
      { mem[2725:2725] } <= { data_i[5:5] };
    end 
    if(N9101) begin
      { mem[2724:2724] } <= { data_i[4:4] };
    end 
    if(N9100) begin
      { mem[2723:2723] } <= { data_i[3:3] };
    end 
    if(N9099) begin
      { mem[2722:2722] } <= { data_i[2:2] };
    end 
    if(N9098) begin
      { mem[2721:2721] } <= { data_i[1:1] };
    end 
    if(N9097) begin
      { mem[2720:2720] } <= { data_i[0:0] };
    end 
    if(N9096) begin
      { mem[2719:2719] } <= { data_i[79:79] };
    end 
    if(N9095) begin
      { mem[2718:2718] } <= { data_i[78:78] };
    end 
    if(N9094) begin
      { mem[2717:2717] } <= { data_i[77:77] };
    end 
    if(N9093) begin
      { mem[2716:2716] } <= { data_i[76:76] };
    end 
    if(N9092) begin
      { mem[2715:2715] } <= { data_i[75:75] };
    end 
    if(N9091) begin
      { mem[2714:2714] } <= { data_i[74:74] };
    end 
    if(N9090) begin
      { mem[2713:2713] } <= { data_i[73:73] };
    end 
    if(N9089) begin
      { mem[2712:2712] } <= { data_i[72:72] };
    end 
    if(N9088) begin
      { mem[2711:2711] } <= { data_i[71:71] };
    end 
    if(N9087) begin
      { mem[2710:2710] } <= { data_i[70:70] };
    end 
    if(N9086) begin
      { mem[2709:2709] } <= { data_i[69:69] };
    end 
    if(N9085) begin
      { mem[2708:2708] } <= { data_i[68:68] };
    end 
    if(N9084) begin
      { mem[2707:2707] } <= { data_i[67:67] };
    end 
    if(N9083) begin
      { mem[2706:2706] } <= { data_i[66:66] };
    end 
    if(N9082) begin
      { mem[2705:2705] } <= { data_i[65:65] };
    end 
    if(N9081) begin
      { mem[2704:2704] } <= { data_i[64:64] };
    end 
    if(N9080) begin
      { mem[2703:2703] } <= { data_i[63:63] };
    end 
    if(N9079) begin
      { mem[2702:2702] } <= { data_i[62:62] };
    end 
    if(N9078) begin
      { mem[2701:2701] } <= { data_i[61:61] };
    end 
    if(N9077) begin
      { mem[2700:2700] } <= { data_i[60:60] };
    end 
    if(N9076) begin
      { mem[2699:2699] } <= { data_i[59:59] };
    end 
    if(N9075) begin
      { mem[2698:2698] } <= { data_i[58:58] };
    end 
    if(N9074) begin
      { mem[2697:2697] } <= { data_i[57:57] };
    end 
    if(N9073) begin
      { mem[2696:2696] } <= { data_i[56:56] };
    end 
    if(N9072) begin
      { mem[2695:2695] } <= { data_i[55:55] };
    end 
    if(N9071) begin
      { mem[2694:2694] } <= { data_i[54:54] };
    end 
    if(N9070) begin
      { mem[2693:2693] } <= { data_i[53:53] };
    end 
    if(N9069) begin
      { mem[2692:2692] } <= { data_i[52:52] };
    end 
    if(N9068) begin
      { mem[2691:2691] } <= { data_i[51:51] };
    end 
    if(N9067) begin
      { mem[2690:2690] } <= { data_i[50:50] };
    end 
    if(N9066) begin
      { mem[2689:2689] } <= { data_i[49:49] };
    end 
    if(N9065) begin
      { mem[2688:2688] } <= { data_i[48:48] };
    end 
    if(N9064) begin
      { mem[2687:2687] } <= { data_i[47:47] };
    end 
    if(N9063) begin
      { mem[2686:2686] } <= { data_i[46:46] };
    end 
    if(N9062) begin
      { mem[2685:2685] } <= { data_i[45:45] };
    end 
    if(N9061) begin
      { mem[2684:2684] } <= { data_i[44:44] };
    end 
    if(N9060) begin
      { mem[2683:2683] } <= { data_i[43:43] };
    end 
    if(N9059) begin
      { mem[2682:2682] } <= { data_i[42:42] };
    end 
    if(N9058) begin
      { mem[2681:2681] } <= { data_i[41:41] };
    end 
    if(N9057) begin
      { mem[2680:2680] } <= { data_i[40:40] };
    end 
    if(N9056) begin
      { mem[2679:2679] } <= { data_i[39:39] };
    end 
    if(N9055) begin
      { mem[2678:2678] } <= { data_i[38:38] };
    end 
    if(N9054) begin
      { mem[2677:2677] } <= { data_i[37:37] };
    end 
    if(N9053) begin
      { mem[2676:2676] } <= { data_i[36:36] };
    end 
    if(N9052) begin
      { mem[2675:2675] } <= { data_i[35:35] };
    end 
    if(N9051) begin
      { mem[2674:2674] } <= { data_i[34:34] };
    end 
    if(N9050) begin
      { mem[2673:2673] } <= { data_i[33:33] };
    end 
    if(N9049) begin
      { mem[2672:2672] } <= { data_i[32:32] };
    end 
    if(N9048) begin
      { mem[2671:2671] } <= { data_i[31:31] };
    end 
    if(N9047) begin
      { mem[2670:2670] } <= { data_i[30:30] };
    end 
    if(N9046) begin
      { mem[2669:2669] } <= { data_i[29:29] };
    end 
    if(N9045) begin
      { mem[2668:2668] } <= { data_i[28:28] };
    end 
    if(N9044) begin
      { mem[2667:2667] } <= { data_i[27:27] };
    end 
    if(N9043) begin
      { mem[2666:2666] } <= { data_i[26:26] };
    end 
    if(N9042) begin
      { mem[2665:2665] } <= { data_i[25:25] };
    end 
    if(N9041) begin
      { mem[2664:2664] } <= { data_i[24:24] };
    end 
    if(N9040) begin
      { mem[2663:2663] } <= { data_i[23:23] };
    end 
    if(N9039) begin
      { mem[2662:2662] } <= { data_i[22:22] };
    end 
    if(N9038) begin
      { mem[2661:2661] } <= { data_i[21:21] };
    end 
    if(N9037) begin
      { mem[2660:2660] } <= { data_i[20:20] };
    end 
    if(N9036) begin
      { mem[2659:2659] } <= { data_i[19:19] };
    end 
    if(N9035) begin
      { mem[2658:2658] } <= { data_i[18:18] };
    end 
    if(N9034) begin
      { mem[2657:2657] } <= { data_i[17:17] };
    end 
    if(N9033) begin
      { mem[2656:2656] } <= { data_i[16:16] };
    end 
    if(N9032) begin
      { mem[2655:2655] } <= { data_i[15:15] };
    end 
    if(N9031) begin
      { mem[2654:2654] } <= { data_i[14:14] };
    end 
    if(N9030) begin
      { mem[2653:2653] } <= { data_i[13:13] };
    end 
    if(N9029) begin
      { mem[2652:2652] } <= { data_i[12:12] };
    end 
    if(N9028) begin
      { mem[2651:2651] } <= { data_i[11:11] };
    end 
    if(N9027) begin
      { mem[2650:2650] } <= { data_i[10:10] };
    end 
    if(N9026) begin
      { mem[2649:2649] } <= { data_i[9:9] };
    end 
    if(N9025) begin
      { mem[2648:2648] } <= { data_i[8:8] };
    end 
    if(N9024) begin
      { mem[2647:2647] } <= { data_i[7:7] };
    end 
    if(N9023) begin
      { mem[2646:2646] } <= { data_i[6:6] };
    end 
    if(N9022) begin
      { mem[2645:2645] } <= { data_i[5:5] };
    end 
    if(N9021) begin
      { mem[2644:2644] } <= { data_i[4:4] };
    end 
    if(N9020) begin
      { mem[2643:2643] } <= { data_i[3:3] };
    end 
    if(N9019) begin
      { mem[2642:2642] } <= { data_i[2:2] };
    end 
    if(N9018) begin
      { mem[2641:2641] } <= { data_i[1:1] };
    end 
    if(N9017) begin
      { mem[2640:2640] } <= { data_i[0:0] };
    end 
    if(N9016) begin
      { mem[2639:2639] } <= { data_i[79:79] };
    end 
    if(N9015) begin
      { mem[2638:2638] } <= { data_i[78:78] };
    end 
    if(N9014) begin
      { mem[2637:2637] } <= { data_i[77:77] };
    end 
    if(N9013) begin
      { mem[2636:2636] } <= { data_i[76:76] };
    end 
    if(N9012) begin
      { mem[2635:2635] } <= { data_i[75:75] };
    end 
    if(N9011) begin
      { mem[2634:2634] } <= { data_i[74:74] };
    end 
    if(N9010) begin
      { mem[2633:2633] } <= { data_i[73:73] };
    end 
    if(N9009) begin
      { mem[2632:2632] } <= { data_i[72:72] };
    end 
    if(N9008) begin
      { mem[2631:2631] } <= { data_i[71:71] };
    end 
    if(N9007) begin
      { mem[2630:2630] } <= { data_i[70:70] };
    end 
    if(N9006) begin
      { mem[2629:2629] } <= { data_i[69:69] };
    end 
    if(N9005) begin
      { mem[2628:2628] } <= { data_i[68:68] };
    end 
    if(N9004) begin
      { mem[2627:2627] } <= { data_i[67:67] };
    end 
    if(N9003) begin
      { mem[2626:2626] } <= { data_i[66:66] };
    end 
    if(N9002) begin
      { mem[2625:2625] } <= { data_i[65:65] };
    end 
    if(N9001) begin
      { mem[2624:2624] } <= { data_i[64:64] };
    end 
    if(N9000) begin
      { mem[2623:2623] } <= { data_i[63:63] };
    end 
    if(N8999) begin
      { mem[2622:2622] } <= { data_i[62:62] };
    end 
    if(N8998) begin
      { mem[2621:2621] } <= { data_i[61:61] };
    end 
    if(N8997) begin
      { mem[2620:2620] } <= { data_i[60:60] };
    end 
    if(N8996) begin
      { mem[2619:2619] } <= { data_i[59:59] };
    end 
    if(N8995) begin
      { mem[2618:2618] } <= { data_i[58:58] };
    end 
    if(N8994) begin
      { mem[2617:2617] } <= { data_i[57:57] };
    end 
    if(N8993) begin
      { mem[2616:2616] } <= { data_i[56:56] };
    end 
    if(N8992) begin
      { mem[2615:2615] } <= { data_i[55:55] };
    end 
    if(N8991) begin
      { mem[2614:2614] } <= { data_i[54:54] };
    end 
    if(N8990) begin
      { mem[2613:2613] } <= { data_i[53:53] };
    end 
    if(N8989) begin
      { mem[2612:2612] } <= { data_i[52:52] };
    end 
    if(N8988) begin
      { mem[2611:2611] } <= { data_i[51:51] };
    end 
    if(N8987) begin
      { mem[2610:2610] } <= { data_i[50:50] };
    end 
    if(N8986) begin
      { mem[2609:2609] } <= { data_i[49:49] };
    end 
    if(N8985) begin
      { mem[2608:2608] } <= { data_i[48:48] };
    end 
    if(N8984) begin
      { mem[2607:2607] } <= { data_i[47:47] };
    end 
    if(N8983) begin
      { mem[2606:2606] } <= { data_i[46:46] };
    end 
    if(N8982) begin
      { mem[2605:2605] } <= { data_i[45:45] };
    end 
    if(N8981) begin
      { mem[2604:2604] } <= { data_i[44:44] };
    end 
    if(N8980) begin
      { mem[2603:2603] } <= { data_i[43:43] };
    end 
    if(N8979) begin
      { mem[2602:2602] } <= { data_i[42:42] };
    end 
    if(N8978) begin
      { mem[2601:2601] } <= { data_i[41:41] };
    end 
    if(N8977) begin
      { mem[2600:2600] } <= { data_i[40:40] };
    end 
    if(N8976) begin
      { mem[2599:2599] } <= { data_i[39:39] };
    end 
    if(N8975) begin
      { mem[2598:2598] } <= { data_i[38:38] };
    end 
    if(N8974) begin
      { mem[2597:2597] } <= { data_i[37:37] };
    end 
    if(N8973) begin
      { mem[2596:2596] } <= { data_i[36:36] };
    end 
    if(N8972) begin
      { mem[2595:2595] } <= { data_i[35:35] };
    end 
    if(N8971) begin
      { mem[2594:2594] } <= { data_i[34:34] };
    end 
    if(N8970) begin
      { mem[2593:2593] } <= { data_i[33:33] };
    end 
    if(N8969) begin
      { mem[2592:2592] } <= { data_i[32:32] };
    end 
    if(N8968) begin
      { mem[2591:2591] } <= { data_i[31:31] };
    end 
    if(N8967) begin
      { mem[2590:2590] } <= { data_i[30:30] };
    end 
    if(N8966) begin
      { mem[2589:2589] } <= { data_i[29:29] };
    end 
    if(N8965) begin
      { mem[2588:2588] } <= { data_i[28:28] };
    end 
    if(N8964) begin
      { mem[2587:2587] } <= { data_i[27:27] };
    end 
    if(N8963) begin
      { mem[2586:2586] } <= { data_i[26:26] };
    end 
    if(N8962) begin
      { mem[2585:2585] } <= { data_i[25:25] };
    end 
    if(N8961) begin
      { mem[2584:2584] } <= { data_i[24:24] };
    end 
    if(N8960) begin
      { mem[2583:2583] } <= { data_i[23:23] };
    end 
    if(N8959) begin
      { mem[2582:2582] } <= { data_i[22:22] };
    end 
    if(N8958) begin
      { mem[2581:2581] } <= { data_i[21:21] };
    end 
    if(N8957) begin
      { mem[2580:2580] } <= { data_i[20:20] };
    end 
    if(N8956) begin
      { mem[2579:2579] } <= { data_i[19:19] };
    end 
    if(N8955) begin
      { mem[2578:2578] } <= { data_i[18:18] };
    end 
    if(N8954) begin
      { mem[2577:2577] } <= { data_i[17:17] };
    end 
    if(N8953) begin
      { mem[2576:2576] } <= { data_i[16:16] };
    end 
    if(N8952) begin
      { mem[2575:2575] } <= { data_i[15:15] };
    end 
    if(N8951) begin
      { mem[2574:2574] } <= { data_i[14:14] };
    end 
    if(N8950) begin
      { mem[2573:2573] } <= { data_i[13:13] };
    end 
    if(N8949) begin
      { mem[2572:2572] } <= { data_i[12:12] };
    end 
    if(N8948) begin
      { mem[2571:2571] } <= { data_i[11:11] };
    end 
    if(N8947) begin
      { mem[2570:2570] } <= { data_i[10:10] };
    end 
    if(N8946) begin
      { mem[2569:2569] } <= { data_i[9:9] };
    end 
    if(N8945) begin
      { mem[2568:2568] } <= { data_i[8:8] };
    end 
    if(N8944) begin
      { mem[2567:2567] } <= { data_i[7:7] };
    end 
    if(N8943) begin
      { mem[2566:2566] } <= { data_i[6:6] };
    end 
    if(N8942) begin
      { mem[2565:2565] } <= { data_i[5:5] };
    end 
    if(N8941) begin
      { mem[2564:2564] } <= { data_i[4:4] };
    end 
    if(N8940) begin
      { mem[2563:2563] } <= { data_i[3:3] };
    end 
    if(N8939) begin
      { mem[2562:2562] } <= { data_i[2:2] };
    end 
    if(N8938) begin
      { mem[2561:2561] } <= { data_i[1:1] };
    end 
    if(N8937) begin
      { mem[2560:2560] } <= { data_i[0:0] };
    end 
    if(N8936) begin
      { mem[2559:2559] } <= { data_i[79:79] };
    end 
    if(N8935) begin
      { mem[2558:2558] } <= { data_i[78:78] };
    end 
    if(N8934) begin
      { mem[2557:2557] } <= { data_i[77:77] };
    end 
    if(N8933) begin
      { mem[2556:2556] } <= { data_i[76:76] };
    end 
    if(N8932) begin
      { mem[2555:2555] } <= { data_i[75:75] };
    end 
    if(N8931) begin
      { mem[2554:2554] } <= { data_i[74:74] };
    end 
    if(N8930) begin
      { mem[2553:2553] } <= { data_i[73:73] };
    end 
    if(N8929) begin
      { mem[2552:2552] } <= { data_i[72:72] };
    end 
    if(N8928) begin
      { mem[2551:2551] } <= { data_i[71:71] };
    end 
    if(N8927) begin
      { mem[2550:2550] } <= { data_i[70:70] };
    end 
    if(N8926) begin
      { mem[2549:2549] } <= { data_i[69:69] };
    end 
    if(N8925) begin
      { mem[2548:2548] } <= { data_i[68:68] };
    end 
    if(N8924) begin
      { mem[2547:2547] } <= { data_i[67:67] };
    end 
    if(N8923) begin
      { mem[2546:2546] } <= { data_i[66:66] };
    end 
    if(N8922) begin
      { mem[2545:2545] } <= { data_i[65:65] };
    end 
    if(N8921) begin
      { mem[2544:2544] } <= { data_i[64:64] };
    end 
    if(N8920) begin
      { mem[2543:2543] } <= { data_i[63:63] };
    end 
    if(N8919) begin
      { mem[2542:2542] } <= { data_i[62:62] };
    end 
    if(N8918) begin
      { mem[2541:2541] } <= { data_i[61:61] };
    end 
    if(N8917) begin
      { mem[2540:2540] } <= { data_i[60:60] };
    end 
    if(N8916) begin
      { mem[2539:2539] } <= { data_i[59:59] };
    end 
    if(N8915) begin
      { mem[2538:2538] } <= { data_i[58:58] };
    end 
    if(N8914) begin
      { mem[2537:2537] } <= { data_i[57:57] };
    end 
    if(N8913) begin
      { mem[2536:2536] } <= { data_i[56:56] };
    end 
    if(N8912) begin
      { mem[2535:2535] } <= { data_i[55:55] };
    end 
    if(N8911) begin
      { mem[2534:2534] } <= { data_i[54:54] };
    end 
    if(N8910) begin
      { mem[2533:2533] } <= { data_i[53:53] };
    end 
    if(N8909) begin
      { mem[2532:2532] } <= { data_i[52:52] };
    end 
    if(N8908) begin
      { mem[2531:2531] } <= { data_i[51:51] };
    end 
    if(N8907) begin
      { mem[2530:2530] } <= { data_i[50:50] };
    end 
    if(N8906) begin
      { mem[2529:2529] } <= { data_i[49:49] };
    end 
    if(N8905) begin
      { mem[2528:2528] } <= { data_i[48:48] };
    end 
    if(N8904) begin
      { mem[2527:2527] } <= { data_i[47:47] };
    end 
    if(N8903) begin
      { mem[2526:2526] } <= { data_i[46:46] };
    end 
    if(N8902) begin
      { mem[2525:2525] } <= { data_i[45:45] };
    end 
    if(N8901) begin
      { mem[2524:2524] } <= { data_i[44:44] };
    end 
    if(N8900) begin
      { mem[2523:2523] } <= { data_i[43:43] };
    end 
    if(N8899) begin
      { mem[2522:2522] } <= { data_i[42:42] };
    end 
    if(N8898) begin
      { mem[2521:2521] } <= { data_i[41:41] };
    end 
    if(N8897) begin
      { mem[2520:2520] } <= { data_i[40:40] };
    end 
    if(N8896) begin
      { mem[2519:2519] } <= { data_i[39:39] };
    end 
    if(N8895) begin
      { mem[2518:2518] } <= { data_i[38:38] };
    end 
    if(N8894) begin
      { mem[2517:2517] } <= { data_i[37:37] };
    end 
    if(N8893) begin
      { mem[2516:2516] } <= { data_i[36:36] };
    end 
    if(N8892) begin
      { mem[2515:2515] } <= { data_i[35:35] };
    end 
    if(N8891) begin
      { mem[2514:2514] } <= { data_i[34:34] };
    end 
    if(N8890) begin
      { mem[2513:2513] } <= { data_i[33:33] };
    end 
    if(N8889) begin
      { mem[2512:2512] } <= { data_i[32:32] };
    end 
    if(N8888) begin
      { mem[2511:2511] } <= { data_i[31:31] };
    end 
    if(N8887) begin
      { mem[2510:2510] } <= { data_i[30:30] };
    end 
    if(N8886) begin
      { mem[2509:2509] } <= { data_i[29:29] };
    end 
    if(N8885) begin
      { mem[2508:2508] } <= { data_i[28:28] };
    end 
    if(N8884) begin
      { mem[2507:2507] } <= { data_i[27:27] };
    end 
    if(N8883) begin
      { mem[2506:2506] } <= { data_i[26:26] };
    end 
    if(N8882) begin
      { mem[2505:2505] } <= { data_i[25:25] };
    end 
    if(N8881) begin
      { mem[2504:2504] } <= { data_i[24:24] };
    end 
    if(N8880) begin
      { mem[2503:2503] } <= { data_i[23:23] };
    end 
    if(N8879) begin
      { mem[2502:2502] } <= { data_i[22:22] };
    end 
    if(N8878) begin
      { mem[2501:2501] } <= { data_i[21:21] };
    end 
    if(N8877) begin
      { mem[2500:2500] } <= { data_i[20:20] };
    end 
    if(N8876) begin
      { mem[2499:2499] } <= { data_i[19:19] };
    end 
    if(N8875) begin
      { mem[2498:2498] } <= { data_i[18:18] };
    end 
    if(N8874) begin
      { mem[2497:2497] } <= { data_i[17:17] };
    end 
    if(N8873) begin
      { mem[2496:2496] } <= { data_i[16:16] };
    end 
    if(N8872) begin
      { mem[2495:2495] } <= { data_i[15:15] };
    end 
    if(N8871) begin
      { mem[2494:2494] } <= { data_i[14:14] };
    end 
    if(N8870) begin
      { mem[2493:2493] } <= { data_i[13:13] };
    end 
    if(N8869) begin
      { mem[2492:2492] } <= { data_i[12:12] };
    end 
    if(N8868) begin
      { mem[2491:2491] } <= { data_i[11:11] };
    end 
    if(N8867) begin
      { mem[2490:2490] } <= { data_i[10:10] };
    end 
    if(N8866) begin
      { mem[2489:2489] } <= { data_i[9:9] };
    end 
    if(N8865) begin
      { mem[2488:2488] } <= { data_i[8:8] };
    end 
    if(N8864) begin
      { mem[2487:2487] } <= { data_i[7:7] };
    end 
    if(N8863) begin
      { mem[2486:2486] } <= { data_i[6:6] };
    end 
    if(N8862) begin
      { mem[2485:2485] } <= { data_i[5:5] };
    end 
    if(N8861) begin
      { mem[2484:2484] } <= { data_i[4:4] };
    end 
    if(N8860) begin
      { mem[2483:2483] } <= { data_i[3:3] };
    end 
    if(N8859) begin
      { mem[2482:2482] } <= { data_i[2:2] };
    end 
    if(N8858) begin
      { mem[2481:2481] } <= { data_i[1:1] };
    end 
    if(N8857) begin
      { mem[2480:2480] } <= { data_i[0:0] };
    end 
    if(N8856) begin
      { mem[2479:2479] } <= { data_i[79:79] };
    end 
    if(N8855) begin
      { mem[2478:2478] } <= { data_i[78:78] };
    end 
    if(N8854) begin
      { mem[2477:2477] } <= { data_i[77:77] };
    end 
    if(N8853) begin
      { mem[2476:2476] } <= { data_i[76:76] };
    end 
    if(N8852) begin
      { mem[2475:2475] } <= { data_i[75:75] };
    end 
    if(N8851) begin
      { mem[2474:2474] } <= { data_i[74:74] };
    end 
    if(N8850) begin
      { mem[2473:2473] } <= { data_i[73:73] };
    end 
    if(N8849) begin
      { mem[2472:2472] } <= { data_i[72:72] };
    end 
    if(N8848) begin
      { mem[2471:2471] } <= { data_i[71:71] };
    end 
    if(N8847) begin
      { mem[2470:2470] } <= { data_i[70:70] };
    end 
    if(N8846) begin
      { mem[2469:2469] } <= { data_i[69:69] };
    end 
    if(N8845) begin
      { mem[2468:2468] } <= { data_i[68:68] };
    end 
    if(N8844) begin
      { mem[2467:2467] } <= { data_i[67:67] };
    end 
    if(N8843) begin
      { mem[2466:2466] } <= { data_i[66:66] };
    end 
    if(N8842) begin
      { mem[2465:2465] } <= { data_i[65:65] };
    end 
    if(N8841) begin
      { mem[2464:2464] } <= { data_i[64:64] };
    end 
    if(N8840) begin
      { mem[2463:2463] } <= { data_i[63:63] };
    end 
    if(N8839) begin
      { mem[2462:2462] } <= { data_i[62:62] };
    end 
    if(N8838) begin
      { mem[2461:2461] } <= { data_i[61:61] };
    end 
    if(N8837) begin
      { mem[2460:2460] } <= { data_i[60:60] };
    end 
    if(N8836) begin
      { mem[2459:2459] } <= { data_i[59:59] };
    end 
    if(N8835) begin
      { mem[2458:2458] } <= { data_i[58:58] };
    end 
    if(N8834) begin
      { mem[2457:2457] } <= { data_i[57:57] };
    end 
    if(N8833) begin
      { mem[2456:2456] } <= { data_i[56:56] };
    end 
    if(N8832) begin
      { mem[2455:2455] } <= { data_i[55:55] };
    end 
    if(N8831) begin
      { mem[2454:2454] } <= { data_i[54:54] };
    end 
    if(N8830) begin
      { mem[2453:2453] } <= { data_i[53:53] };
    end 
    if(N8829) begin
      { mem[2452:2452] } <= { data_i[52:52] };
    end 
    if(N8828) begin
      { mem[2451:2451] } <= { data_i[51:51] };
    end 
    if(N8827) begin
      { mem[2450:2450] } <= { data_i[50:50] };
    end 
    if(N8826) begin
      { mem[2449:2449] } <= { data_i[49:49] };
    end 
    if(N8825) begin
      { mem[2448:2448] } <= { data_i[48:48] };
    end 
    if(N8824) begin
      { mem[2447:2447] } <= { data_i[47:47] };
    end 
    if(N8823) begin
      { mem[2446:2446] } <= { data_i[46:46] };
    end 
    if(N8822) begin
      { mem[2445:2445] } <= { data_i[45:45] };
    end 
    if(N8821) begin
      { mem[2444:2444] } <= { data_i[44:44] };
    end 
    if(N8820) begin
      { mem[2443:2443] } <= { data_i[43:43] };
    end 
    if(N8819) begin
      { mem[2442:2442] } <= { data_i[42:42] };
    end 
    if(N8818) begin
      { mem[2441:2441] } <= { data_i[41:41] };
    end 
    if(N8817) begin
      { mem[2440:2440] } <= { data_i[40:40] };
    end 
    if(N8816) begin
      { mem[2439:2439] } <= { data_i[39:39] };
    end 
    if(N8815) begin
      { mem[2438:2438] } <= { data_i[38:38] };
    end 
    if(N8814) begin
      { mem[2437:2437] } <= { data_i[37:37] };
    end 
    if(N8813) begin
      { mem[2436:2436] } <= { data_i[36:36] };
    end 
    if(N8812) begin
      { mem[2435:2435] } <= { data_i[35:35] };
    end 
    if(N8811) begin
      { mem[2434:2434] } <= { data_i[34:34] };
    end 
    if(N8810) begin
      { mem[2433:2433] } <= { data_i[33:33] };
    end 
    if(N8809) begin
      { mem[2432:2432] } <= { data_i[32:32] };
    end 
    if(N8808) begin
      { mem[2431:2431] } <= { data_i[31:31] };
    end 
    if(N8807) begin
      { mem[2430:2430] } <= { data_i[30:30] };
    end 
    if(N8806) begin
      { mem[2429:2429] } <= { data_i[29:29] };
    end 
    if(N8805) begin
      { mem[2428:2428] } <= { data_i[28:28] };
    end 
    if(N8804) begin
      { mem[2427:2427] } <= { data_i[27:27] };
    end 
    if(N8803) begin
      { mem[2426:2426] } <= { data_i[26:26] };
    end 
    if(N8802) begin
      { mem[2425:2425] } <= { data_i[25:25] };
    end 
    if(N8801) begin
      { mem[2424:2424] } <= { data_i[24:24] };
    end 
    if(N8800) begin
      { mem[2423:2423] } <= { data_i[23:23] };
    end 
    if(N8799) begin
      { mem[2422:2422] } <= { data_i[22:22] };
    end 
    if(N8798) begin
      { mem[2421:2421] } <= { data_i[21:21] };
    end 
    if(N8797) begin
      { mem[2420:2420] } <= { data_i[20:20] };
    end 
    if(N8796) begin
      { mem[2419:2419] } <= { data_i[19:19] };
    end 
    if(N8795) begin
      { mem[2418:2418] } <= { data_i[18:18] };
    end 
    if(N8794) begin
      { mem[2417:2417] } <= { data_i[17:17] };
    end 
    if(N8793) begin
      { mem[2416:2416] } <= { data_i[16:16] };
    end 
    if(N8792) begin
      { mem[2415:2415] } <= { data_i[15:15] };
    end 
    if(N8791) begin
      { mem[2414:2414] } <= { data_i[14:14] };
    end 
    if(N8790) begin
      { mem[2413:2413] } <= { data_i[13:13] };
    end 
    if(N8789) begin
      { mem[2412:2412] } <= { data_i[12:12] };
    end 
    if(N8788) begin
      { mem[2411:2411] } <= { data_i[11:11] };
    end 
    if(N8787) begin
      { mem[2410:2410] } <= { data_i[10:10] };
    end 
    if(N8786) begin
      { mem[2409:2409] } <= { data_i[9:9] };
    end 
    if(N8785) begin
      { mem[2408:2408] } <= { data_i[8:8] };
    end 
    if(N8784) begin
      { mem[2407:2407] } <= { data_i[7:7] };
    end 
    if(N8783) begin
      { mem[2406:2406] } <= { data_i[6:6] };
    end 
    if(N8782) begin
      { mem[2405:2405] } <= { data_i[5:5] };
    end 
    if(N8781) begin
      { mem[2404:2404] } <= { data_i[4:4] };
    end 
    if(N8780) begin
      { mem[2403:2403] } <= { data_i[3:3] };
    end 
    if(N8779) begin
      { mem[2402:2402] } <= { data_i[2:2] };
    end 
    if(N8778) begin
      { mem[2401:2401] } <= { data_i[1:1] };
    end 
    if(N8777) begin
      { mem[2400:2400] } <= { data_i[0:0] };
    end 
    if(N8776) begin
      { mem[2399:2399] } <= { data_i[79:79] };
    end 
    if(N8775) begin
      { mem[2398:2398] } <= { data_i[78:78] };
    end 
    if(N8774) begin
      { mem[2397:2397] } <= { data_i[77:77] };
    end 
    if(N8773) begin
      { mem[2396:2396] } <= { data_i[76:76] };
    end 
    if(N8772) begin
      { mem[2395:2395] } <= { data_i[75:75] };
    end 
    if(N8771) begin
      { mem[2394:2394] } <= { data_i[74:74] };
    end 
    if(N8770) begin
      { mem[2393:2393] } <= { data_i[73:73] };
    end 
    if(N8769) begin
      { mem[2392:2392] } <= { data_i[72:72] };
    end 
    if(N8768) begin
      { mem[2391:2391] } <= { data_i[71:71] };
    end 
    if(N8767) begin
      { mem[2390:2390] } <= { data_i[70:70] };
    end 
    if(N8766) begin
      { mem[2389:2389] } <= { data_i[69:69] };
    end 
    if(N8765) begin
      { mem[2388:2388] } <= { data_i[68:68] };
    end 
    if(N8764) begin
      { mem[2387:2387] } <= { data_i[67:67] };
    end 
    if(N8763) begin
      { mem[2386:2386] } <= { data_i[66:66] };
    end 
    if(N8762) begin
      { mem[2385:2385] } <= { data_i[65:65] };
    end 
    if(N8761) begin
      { mem[2384:2384] } <= { data_i[64:64] };
    end 
    if(N8760) begin
      { mem[2383:2383] } <= { data_i[63:63] };
    end 
    if(N8759) begin
      { mem[2382:2382] } <= { data_i[62:62] };
    end 
    if(N8758) begin
      { mem[2381:2381] } <= { data_i[61:61] };
    end 
    if(N8757) begin
      { mem[2380:2380] } <= { data_i[60:60] };
    end 
    if(N8756) begin
      { mem[2379:2379] } <= { data_i[59:59] };
    end 
    if(N8755) begin
      { mem[2378:2378] } <= { data_i[58:58] };
    end 
    if(N8754) begin
      { mem[2377:2377] } <= { data_i[57:57] };
    end 
    if(N8753) begin
      { mem[2376:2376] } <= { data_i[56:56] };
    end 
    if(N8752) begin
      { mem[2375:2375] } <= { data_i[55:55] };
    end 
    if(N8751) begin
      { mem[2374:2374] } <= { data_i[54:54] };
    end 
    if(N8750) begin
      { mem[2373:2373] } <= { data_i[53:53] };
    end 
    if(N8749) begin
      { mem[2372:2372] } <= { data_i[52:52] };
    end 
    if(N8748) begin
      { mem[2371:2371] } <= { data_i[51:51] };
    end 
    if(N8747) begin
      { mem[2370:2370] } <= { data_i[50:50] };
    end 
    if(N8746) begin
      { mem[2369:2369] } <= { data_i[49:49] };
    end 
    if(N8745) begin
      { mem[2368:2368] } <= { data_i[48:48] };
    end 
    if(N8744) begin
      { mem[2367:2367] } <= { data_i[47:47] };
    end 
    if(N8743) begin
      { mem[2366:2366] } <= { data_i[46:46] };
    end 
    if(N8742) begin
      { mem[2365:2365] } <= { data_i[45:45] };
    end 
    if(N8741) begin
      { mem[2364:2364] } <= { data_i[44:44] };
    end 
    if(N8740) begin
      { mem[2363:2363] } <= { data_i[43:43] };
    end 
    if(N8739) begin
      { mem[2362:2362] } <= { data_i[42:42] };
    end 
    if(N8738) begin
      { mem[2361:2361] } <= { data_i[41:41] };
    end 
    if(N8737) begin
      { mem[2360:2360] } <= { data_i[40:40] };
    end 
    if(N8736) begin
      { mem[2359:2359] } <= { data_i[39:39] };
    end 
    if(N8735) begin
      { mem[2358:2358] } <= { data_i[38:38] };
    end 
    if(N8734) begin
      { mem[2357:2357] } <= { data_i[37:37] };
    end 
    if(N8733) begin
      { mem[2356:2356] } <= { data_i[36:36] };
    end 
    if(N8732) begin
      { mem[2355:2355] } <= { data_i[35:35] };
    end 
    if(N8731) begin
      { mem[2354:2354] } <= { data_i[34:34] };
    end 
    if(N8730) begin
      { mem[2353:2353] } <= { data_i[33:33] };
    end 
    if(N8729) begin
      { mem[2352:2352] } <= { data_i[32:32] };
    end 
    if(N8728) begin
      { mem[2351:2351] } <= { data_i[31:31] };
    end 
    if(N8727) begin
      { mem[2350:2350] } <= { data_i[30:30] };
    end 
    if(N8726) begin
      { mem[2349:2349] } <= { data_i[29:29] };
    end 
    if(N8725) begin
      { mem[2348:2348] } <= { data_i[28:28] };
    end 
    if(N8724) begin
      { mem[2347:2347] } <= { data_i[27:27] };
    end 
    if(N8723) begin
      { mem[2346:2346] } <= { data_i[26:26] };
    end 
    if(N8722) begin
      { mem[2345:2345] } <= { data_i[25:25] };
    end 
    if(N8721) begin
      { mem[2344:2344] } <= { data_i[24:24] };
    end 
    if(N8720) begin
      { mem[2343:2343] } <= { data_i[23:23] };
    end 
    if(N8719) begin
      { mem[2342:2342] } <= { data_i[22:22] };
    end 
    if(N8718) begin
      { mem[2341:2341] } <= { data_i[21:21] };
    end 
    if(N8717) begin
      { mem[2340:2340] } <= { data_i[20:20] };
    end 
    if(N8716) begin
      { mem[2339:2339] } <= { data_i[19:19] };
    end 
    if(N8715) begin
      { mem[2338:2338] } <= { data_i[18:18] };
    end 
    if(N8714) begin
      { mem[2337:2337] } <= { data_i[17:17] };
    end 
    if(N8713) begin
      { mem[2336:2336] } <= { data_i[16:16] };
    end 
    if(N8712) begin
      { mem[2335:2335] } <= { data_i[15:15] };
    end 
    if(N8711) begin
      { mem[2334:2334] } <= { data_i[14:14] };
    end 
    if(N8710) begin
      { mem[2333:2333] } <= { data_i[13:13] };
    end 
    if(N8709) begin
      { mem[2332:2332] } <= { data_i[12:12] };
    end 
    if(N8708) begin
      { mem[2331:2331] } <= { data_i[11:11] };
    end 
    if(N8707) begin
      { mem[2330:2330] } <= { data_i[10:10] };
    end 
    if(N8706) begin
      { mem[2329:2329] } <= { data_i[9:9] };
    end 
    if(N8705) begin
      { mem[2328:2328] } <= { data_i[8:8] };
    end 
    if(N8704) begin
      { mem[2327:2327] } <= { data_i[7:7] };
    end 
    if(N8703) begin
      { mem[2326:2326] } <= { data_i[6:6] };
    end 
    if(N8702) begin
      { mem[2325:2325] } <= { data_i[5:5] };
    end 
    if(N8701) begin
      { mem[2324:2324] } <= { data_i[4:4] };
    end 
    if(N8700) begin
      { mem[2323:2323] } <= { data_i[3:3] };
    end 
    if(N8699) begin
      { mem[2322:2322] } <= { data_i[2:2] };
    end 
    if(N8698) begin
      { mem[2321:2321] } <= { data_i[1:1] };
    end 
    if(N8697) begin
      { mem[2320:2320] } <= { data_i[0:0] };
    end 
    if(N8696) begin
      { mem[2319:2319] } <= { data_i[79:79] };
    end 
    if(N8695) begin
      { mem[2318:2318] } <= { data_i[78:78] };
    end 
    if(N8694) begin
      { mem[2317:2317] } <= { data_i[77:77] };
    end 
    if(N8693) begin
      { mem[2316:2316] } <= { data_i[76:76] };
    end 
    if(N8692) begin
      { mem[2315:2315] } <= { data_i[75:75] };
    end 
    if(N8691) begin
      { mem[2314:2314] } <= { data_i[74:74] };
    end 
    if(N8690) begin
      { mem[2313:2313] } <= { data_i[73:73] };
    end 
    if(N8689) begin
      { mem[2312:2312] } <= { data_i[72:72] };
    end 
    if(N8688) begin
      { mem[2311:2311] } <= { data_i[71:71] };
    end 
    if(N8687) begin
      { mem[2310:2310] } <= { data_i[70:70] };
    end 
    if(N8686) begin
      { mem[2309:2309] } <= { data_i[69:69] };
    end 
    if(N8685) begin
      { mem[2308:2308] } <= { data_i[68:68] };
    end 
    if(N8684) begin
      { mem[2307:2307] } <= { data_i[67:67] };
    end 
    if(N8683) begin
      { mem[2306:2306] } <= { data_i[66:66] };
    end 
    if(N8682) begin
      { mem[2305:2305] } <= { data_i[65:65] };
    end 
    if(N8681) begin
      { mem[2304:2304] } <= { data_i[64:64] };
    end 
    if(N8680) begin
      { mem[2303:2303] } <= { data_i[63:63] };
    end 
    if(N8679) begin
      { mem[2302:2302] } <= { data_i[62:62] };
    end 
    if(N8678) begin
      { mem[2301:2301] } <= { data_i[61:61] };
    end 
    if(N8677) begin
      { mem[2300:2300] } <= { data_i[60:60] };
    end 
    if(N8676) begin
      { mem[2299:2299] } <= { data_i[59:59] };
    end 
    if(N8675) begin
      { mem[2298:2298] } <= { data_i[58:58] };
    end 
    if(N8674) begin
      { mem[2297:2297] } <= { data_i[57:57] };
    end 
    if(N8673) begin
      { mem[2296:2296] } <= { data_i[56:56] };
    end 
    if(N8672) begin
      { mem[2295:2295] } <= { data_i[55:55] };
    end 
    if(N8671) begin
      { mem[2294:2294] } <= { data_i[54:54] };
    end 
    if(N8670) begin
      { mem[2293:2293] } <= { data_i[53:53] };
    end 
    if(N8669) begin
      { mem[2292:2292] } <= { data_i[52:52] };
    end 
    if(N8668) begin
      { mem[2291:2291] } <= { data_i[51:51] };
    end 
    if(N8667) begin
      { mem[2290:2290] } <= { data_i[50:50] };
    end 
    if(N8666) begin
      { mem[2289:2289] } <= { data_i[49:49] };
    end 
    if(N8665) begin
      { mem[2288:2288] } <= { data_i[48:48] };
    end 
    if(N8664) begin
      { mem[2287:2287] } <= { data_i[47:47] };
    end 
    if(N8663) begin
      { mem[2286:2286] } <= { data_i[46:46] };
    end 
    if(N8662) begin
      { mem[2285:2285] } <= { data_i[45:45] };
    end 
    if(N8661) begin
      { mem[2284:2284] } <= { data_i[44:44] };
    end 
    if(N8660) begin
      { mem[2283:2283] } <= { data_i[43:43] };
    end 
    if(N8659) begin
      { mem[2282:2282] } <= { data_i[42:42] };
    end 
    if(N8658) begin
      { mem[2281:2281] } <= { data_i[41:41] };
    end 
    if(N8657) begin
      { mem[2280:2280] } <= { data_i[40:40] };
    end 
    if(N8656) begin
      { mem[2279:2279] } <= { data_i[39:39] };
    end 
    if(N8655) begin
      { mem[2278:2278] } <= { data_i[38:38] };
    end 
    if(N8654) begin
      { mem[2277:2277] } <= { data_i[37:37] };
    end 
    if(N8653) begin
      { mem[2276:2276] } <= { data_i[36:36] };
    end 
    if(N8652) begin
      { mem[2275:2275] } <= { data_i[35:35] };
    end 
    if(N8651) begin
      { mem[2274:2274] } <= { data_i[34:34] };
    end 
    if(N8650) begin
      { mem[2273:2273] } <= { data_i[33:33] };
    end 
    if(N8649) begin
      { mem[2272:2272] } <= { data_i[32:32] };
    end 
    if(N8648) begin
      { mem[2271:2271] } <= { data_i[31:31] };
    end 
    if(N8647) begin
      { mem[2270:2270] } <= { data_i[30:30] };
    end 
    if(N8646) begin
      { mem[2269:2269] } <= { data_i[29:29] };
    end 
    if(N8645) begin
      { mem[2268:2268] } <= { data_i[28:28] };
    end 
    if(N8644) begin
      { mem[2267:2267] } <= { data_i[27:27] };
    end 
    if(N8643) begin
      { mem[2266:2266] } <= { data_i[26:26] };
    end 
    if(N8642) begin
      { mem[2265:2265] } <= { data_i[25:25] };
    end 
    if(N8641) begin
      { mem[2264:2264] } <= { data_i[24:24] };
    end 
    if(N8640) begin
      { mem[2263:2263] } <= { data_i[23:23] };
    end 
    if(N8639) begin
      { mem[2262:2262] } <= { data_i[22:22] };
    end 
    if(N8638) begin
      { mem[2261:2261] } <= { data_i[21:21] };
    end 
    if(N8637) begin
      { mem[2260:2260] } <= { data_i[20:20] };
    end 
    if(N8636) begin
      { mem[2259:2259] } <= { data_i[19:19] };
    end 
    if(N8635) begin
      { mem[2258:2258] } <= { data_i[18:18] };
    end 
    if(N8634) begin
      { mem[2257:2257] } <= { data_i[17:17] };
    end 
    if(N8633) begin
      { mem[2256:2256] } <= { data_i[16:16] };
    end 
    if(N8632) begin
      { mem[2255:2255] } <= { data_i[15:15] };
    end 
    if(N8631) begin
      { mem[2254:2254] } <= { data_i[14:14] };
    end 
    if(N8630) begin
      { mem[2253:2253] } <= { data_i[13:13] };
    end 
    if(N8629) begin
      { mem[2252:2252] } <= { data_i[12:12] };
    end 
    if(N8628) begin
      { mem[2251:2251] } <= { data_i[11:11] };
    end 
    if(N8627) begin
      { mem[2250:2250] } <= { data_i[10:10] };
    end 
    if(N8626) begin
      { mem[2249:2249] } <= { data_i[9:9] };
    end 
    if(N8625) begin
      { mem[2248:2248] } <= { data_i[8:8] };
    end 
    if(N8624) begin
      { mem[2247:2247] } <= { data_i[7:7] };
    end 
    if(N8623) begin
      { mem[2246:2246] } <= { data_i[6:6] };
    end 
    if(N8622) begin
      { mem[2245:2245] } <= { data_i[5:5] };
    end 
    if(N8621) begin
      { mem[2244:2244] } <= { data_i[4:4] };
    end 
    if(N8620) begin
      { mem[2243:2243] } <= { data_i[3:3] };
    end 
    if(N8619) begin
      { mem[2242:2242] } <= { data_i[2:2] };
    end 
    if(N8618) begin
      { mem[2241:2241] } <= { data_i[1:1] };
    end 
    if(N8617) begin
      { mem[2240:2240] } <= { data_i[0:0] };
    end 
    if(N8616) begin
      { mem[2239:2239] } <= { data_i[79:79] };
    end 
    if(N8615) begin
      { mem[2238:2238] } <= { data_i[78:78] };
    end 
    if(N8614) begin
      { mem[2237:2237] } <= { data_i[77:77] };
    end 
    if(N8613) begin
      { mem[2236:2236] } <= { data_i[76:76] };
    end 
    if(N8612) begin
      { mem[2235:2235] } <= { data_i[75:75] };
    end 
    if(N8611) begin
      { mem[2234:2234] } <= { data_i[74:74] };
    end 
    if(N8610) begin
      { mem[2233:2233] } <= { data_i[73:73] };
    end 
    if(N8609) begin
      { mem[2232:2232] } <= { data_i[72:72] };
    end 
    if(N8608) begin
      { mem[2231:2231] } <= { data_i[71:71] };
    end 
    if(N8607) begin
      { mem[2230:2230] } <= { data_i[70:70] };
    end 
    if(N8606) begin
      { mem[2229:2229] } <= { data_i[69:69] };
    end 
    if(N8605) begin
      { mem[2228:2228] } <= { data_i[68:68] };
    end 
    if(N8604) begin
      { mem[2227:2227] } <= { data_i[67:67] };
    end 
    if(N8603) begin
      { mem[2226:2226] } <= { data_i[66:66] };
    end 
    if(N8602) begin
      { mem[2225:2225] } <= { data_i[65:65] };
    end 
    if(N8601) begin
      { mem[2224:2224] } <= { data_i[64:64] };
    end 
    if(N8600) begin
      { mem[2223:2223] } <= { data_i[63:63] };
    end 
    if(N8599) begin
      { mem[2222:2222] } <= { data_i[62:62] };
    end 
    if(N8598) begin
      { mem[2221:2221] } <= { data_i[61:61] };
    end 
    if(N8597) begin
      { mem[2220:2220] } <= { data_i[60:60] };
    end 
    if(N8596) begin
      { mem[2219:2219] } <= { data_i[59:59] };
    end 
    if(N8595) begin
      { mem[2218:2218] } <= { data_i[58:58] };
    end 
    if(N8594) begin
      { mem[2217:2217] } <= { data_i[57:57] };
    end 
    if(N8593) begin
      { mem[2216:2216] } <= { data_i[56:56] };
    end 
    if(N8592) begin
      { mem[2215:2215] } <= { data_i[55:55] };
    end 
    if(N8591) begin
      { mem[2214:2214] } <= { data_i[54:54] };
    end 
    if(N8590) begin
      { mem[2213:2213] } <= { data_i[53:53] };
    end 
    if(N8589) begin
      { mem[2212:2212] } <= { data_i[52:52] };
    end 
    if(N8588) begin
      { mem[2211:2211] } <= { data_i[51:51] };
    end 
    if(N8587) begin
      { mem[2210:2210] } <= { data_i[50:50] };
    end 
    if(N8586) begin
      { mem[2209:2209] } <= { data_i[49:49] };
    end 
    if(N8585) begin
      { mem[2208:2208] } <= { data_i[48:48] };
    end 
    if(N8584) begin
      { mem[2207:2207] } <= { data_i[47:47] };
    end 
    if(N8583) begin
      { mem[2206:2206] } <= { data_i[46:46] };
    end 
    if(N8582) begin
      { mem[2205:2205] } <= { data_i[45:45] };
    end 
    if(N8581) begin
      { mem[2204:2204] } <= { data_i[44:44] };
    end 
    if(N8580) begin
      { mem[2203:2203] } <= { data_i[43:43] };
    end 
    if(N8579) begin
      { mem[2202:2202] } <= { data_i[42:42] };
    end 
    if(N8578) begin
      { mem[2201:2201] } <= { data_i[41:41] };
    end 
    if(N8577) begin
      { mem[2200:2200] } <= { data_i[40:40] };
    end 
    if(N8576) begin
      { mem[2199:2199] } <= { data_i[39:39] };
    end 
    if(N8575) begin
      { mem[2198:2198] } <= { data_i[38:38] };
    end 
    if(N8574) begin
      { mem[2197:2197] } <= { data_i[37:37] };
    end 
    if(N8573) begin
      { mem[2196:2196] } <= { data_i[36:36] };
    end 
    if(N8572) begin
      { mem[2195:2195] } <= { data_i[35:35] };
    end 
    if(N8571) begin
      { mem[2194:2194] } <= { data_i[34:34] };
    end 
    if(N8570) begin
      { mem[2193:2193] } <= { data_i[33:33] };
    end 
    if(N8569) begin
      { mem[2192:2192] } <= { data_i[32:32] };
    end 
    if(N8568) begin
      { mem[2191:2191] } <= { data_i[31:31] };
    end 
    if(N8567) begin
      { mem[2190:2190] } <= { data_i[30:30] };
    end 
    if(N8566) begin
      { mem[2189:2189] } <= { data_i[29:29] };
    end 
    if(N8565) begin
      { mem[2188:2188] } <= { data_i[28:28] };
    end 
    if(N8564) begin
      { mem[2187:2187] } <= { data_i[27:27] };
    end 
    if(N8563) begin
      { mem[2186:2186] } <= { data_i[26:26] };
    end 
    if(N8562) begin
      { mem[2185:2185] } <= { data_i[25:25] };
    end 
    if(N8561) begin
      { mem[2184:2184] } <= { data_i[24:24] };
    end 
    if(N8560) begin
      { mem[2183:2183] } <= { data_i[23:23] };
    end 
    if(N8559) begin
      { mem[2182:2182] } <= { data_i[22:22] };
    end 
    if(N8558) begin
      { mem[2181:2181] } <= { data_i[21:21] };
    end 
    if(N8557) begin
      { mem[2180:2180] } <= { data_i[20:20] };
    end 
    if(N8556) begin
      { mem[2179:2179] } <= { data_i[19:19] };
    end 
    if(N8555) begin
      { mem[2178:2178] } <= { data_i[18:18] };
    end 
    if(N8554) begin
      { mem[2177:2177] } <= { data_i[17:17] };
    end 
    if(N8553) begin
      { mem[2176:2176] } <= { data_i[16:16] };
    end 
    if(N8552) begin
      { mem[2175:2175] } <= { data_i[15:15] };
    end 
    if(N8551) begin
      { mem[2174:2174] } <= { data_i[14:14] };
    end 
    if(N8550) begin
      { mem[2173:2173] } <= { data_i[13:13] };
    end 
    if(N8549) begin
      { mem[2172:2172] } <= { data_i[12:12] };
    end 
    if(N8548) begin
      { mem[2171:2171] } <= { data_i[11:11] };
    end 
    if(N8547) begin
      { mem[2170:2170] } <= { data_i[10:10] };
    end 
    if(N8546) begin
      { mem[2169:2169] } <= { data_i[9:9] };
    end 
    if(N8545) begin
      { mem[2168:2168] } <= { data_i[8:8] };
    end 
    if(N8544) begin
      { mem[2167:2167] } <= { data_i[7:7] };
    end 
    if(N8543) begin
      { mem[2166:2166] } <= { data_i[6:6] };
    end 
    if(N8542) begin
      { mem[2165:2165] } <= { data_i[5:5] };
    end 
    if(N8541) begin
      { mem[2164:2164] } <= { data_i[4:4] };
    end 
    if(N8540) begin
      { mem[2163:2163] } <= { data_i[3:3] };
    end 
    if(N8539) begin
      { mem[2162:2162] } <= { data_i[2:2] };
    end 
    if(N8538) begin
      { mem[2161:2161] } <= { data_i[1:1] };
    end 
    if(N8537) begin
      { mem[2160:2160] } <= { data_i[0:0] };
    end 
    if(N8536) begin
      { mem[2159:2159] } <= { data_i[79:79] };
    end 
    if(N8535) begin
      { mem[2158:2158] } <= { data_i[78:78] };
    end 
    if(N8534) begin
      { mem[2157:2157] } <= { data_i[77:77] };
    end 
    if(N8533) begin
      { mem[2156:2156] } <= { data_i[76:76] };
    end 
    if(N8532) begin
      { mem[2155:2155] } <= { data_i[75:75] };
    end 
    if(N8531) begin
      { mem[2154:2154] } <= { data_i[74:74] };
    end 
    if(N8530) begin
      { mem[2153:2153] } <= { data_i[73:73] };
    end 
    if(N8529) begin
      { mem[2152:2152] } <= { data_i[72:72] };
    end 
    if(N8528) begin
      { mem[2151:2151] } <= { data_i[71:71] };
    end 
    if(N8527) begin
      { mem[2150:2150] } <= { data_i[70:70] };
    end 
    if(N8526) begin
      { mem[2149:2149] } <= { data_i[69:69] };
    end 
    if(N8525) begin
      { mem[2148:2148] } <= { data_i[68:68] };
    end 
    if(N8524) begin
      { mem[2147:2147] } <= { data_i[67:67] };
    end 
    if(N8523) begin
      { mem[2146:2146] } <= { data_i[66:66] };
    end 
    if(N8522) begin
      { mem[2145:2145] } <= { data_i[65:65] };
    end 
    if(N8521) begin
      { mem[2144:2144] } <= { data_i[64:64] };
    end 
    if(N8520) begin
      { mem[2143:2143] } <= { data_i[63:63] };
    end 
    if(N8519) begin
      { mem[2142:2142] } <= { data_i[62:62] };
    end 
    if(N8518) begin
      { mem[2141:2141] } <= { data_i[61:61] };
    end 
    if(N8517) begin
      { mem[2140:2140] } <= { data_i[60:60] };
    end 
    if(N8516) begin
      { mem[2139:2139] } <= { data_i[59:59] };
    end 
    if(N8515) begin
      { mem[2138:2138] } <= { data_i[58:58] };
    end 
    if(N8514) begin
      { mem[2137:2137] } <= { data_i[57:57] };
    end 
    if(N8513) begin
      { mem[2136:2136] } <= { data_i[56:56] };
    end 
    if(N8512) begin
      { mem[2135:2135] } <= { data_i[55:55] };
    end 
    if(N8511) begin
      { mem[2134:2134] } <= { data_i[54:54] };
    end 
    if(N8510) begin
      { mem[2133:2133] } <= { data_i[53:53] };
    end 
    if(N8509) begin
      { mem[2132:2132] } <= { data_i[52:52] };
    end 
    if(N8508) begin
      { mem[2131:2131] } <= { data_i[51:51] };
    end 
    if(N8507) begin
      { mem[2130:2130] } <= { data_i[50:50] };
    end 
    if(N8506) begin
      { mem[2129:2129] } <= { data_i[49:49] };
    end 
    if(N8505) begin
      { mem[2128:2128] } <= { data_i[48:48] };
    end 
    if(N8504) begin
      { mem[2127:2127] } <= { data_i[47:47] };
    end 
    if(N8503) begin
      { mem[2126:2126] } <= { data_i[46:46] };
    end 
    if(N8502) begin
      { mem[2125:2125] } <= { data_i[45:45] };
    end 
    if(N8501) begin
      { mem[2124:2124] } <= { data_i[44:44] };
    end 
    if(N8500) begin
      { mem[2123:2123] } <= { data_i[43:43] };
    end 
    if(N8499) begin
      { mem[2122:2122] } <= { data_i[42:42] };
    end 
    if(N8498) begin
      { mem[2121:2121] } <= { data_i[41:41] };
    end 
    if(N8497) begin
      { mem[2120:2120] } <= { data_i[40:40] };
    end 
    if(N8496) begin
      { mem[2119:2119] } <= { data_i[39:39] };
    end 
    if(N8495) begin
      { mem[2118:2118] } <= { data_i[38:38] };
    end 
    if(N8494) begin
      { mem[2117:2117] } <= { data_i[37:37] };
    end 
    if(N8493) begin
      { mem[2116:2116] } <= { data_i[36:36] };
    end 
    if(N8492) begin
      { mem[2115:2115] } <= { data_i[35:35] };
    end 
    if(N8491) begin
      { mem[2114:2114] } <= { data_i[34:34] };
    end 
    if(N8490) begin
      { mem[2113:2113] } <= { data_i[33:33] };
    end 
    if(N8489) begin
      { mem[2112:2112] } <= { data_i[32:32] };
    end 
    if(N8488) begin
      { mem[2111:2111] } <= { data_i[31:31] };
    end 
    if(N8487) begin
      { mem[2110:2110] } <= { data_i[30:30] };
    end 
    if(N8486) begin
      { mem[2109:2109] } <= { data_i[29:29] };
    end 
    if(N8485) begin
      { mem[2108:2108] } <= { data_i[28:28] };
    end 
    if(N8484) begin
      { mem[2107:2107] } <= { data_i[27:27] };
    end 
    if(N8483) begin
      { mem[2106:2106] } <= { data_i[26:26] };
    end 
    if(N8482) begin
      { mem[2105:2105] } <= { data_i[25:25] };
    end 
    if(N8481) begin
      { mem[2104:2104] } <= { data_i[24:24] };
    end 
    if(N8480) begin
      { mem[2103:2103] } <= { data_i[23:23] };
    end 
    if(N8479) begin
      { mem[2102:2102] } <= { data_i[22:22] };
    end 
    if(N8478) begin
      { mem[2101:2101] } <= { data_i[21:21] };
    end 
    if(N8477) begin
      { mem[2100:2100] } <= { data_i[20:20] };
    end 
    if(N8476) begin
      { mem[2099:2099] } <= { data_i[19:19] };
    end 
    if(N8475) begin
      { mem[2098:2098] } <= { data_i[18:18] };
    end 
    if(N8474) begin
      { mem[2097:2097] } <= { data_i[17:17] };
    end 
    if(N8473) begin
      { mem[2096:2096] } <= { data_i[16:16] };
    end 
    if(N8472) begin
      { mem[2095:2095] } <= { data_i[15:15] };
    end 
    if(N8471) begin
      { mem[2094:2094] } <= { data_i[14:14] };
    end 
    if(N8470) begin
      { mem[2093:2093] } <= { data_i[13:13] };
    end 
    if(N8469) begin
      { mem[2092:2092] } <= { data_i[12:12] };
    end 
    if(N8468) begin
      { mem[2091:2091] } <= { data_i[11:11] };
    end 
    if(N8467) begin
      { mem[2090:2090] } <= { data_i[10:10] };
    end 
    if(N8466) begin
      { mem[2089:2089] } <= { data_i[9:9] };
    end 
    if(N8465) begin
      { mem[2088:2088] } <= { data_i[8:8] };
    end 
    if(N8464) begin
      { mem[2087:2087] } <= { data_i[7:7] };
    end 
    if(N8463) begin
      { mem[2086:2086] } <= { data_i[6:6] };
    end 
    if(N8462) begin
      { mem[2085:2085] } <= { data_i[5:5] };
    end 
    if(N8461) begin
      { mem[2084:2084] } <= { data_i[4:4] };
    end 
    if(N8460) begin
      { mem[2083:2083] } <= { data_i[3:3] };
    end 
    if(N8459) begin
      { mem[2082:2082] } <= { data_i[2:2] };
    end 
    if(N8458) begin
      { mem[2081:2081] } <= { data_i[1:1] };
    end 
    if(N8457) begin
      { mem[2080:2080] } <= { data_i[0:0] };
    end 
    if(N8456) begin
      { mem[2079:2079] } <= { data_i[79:79] };
    end 
    if(N8455) begin
      { mem[2078:2078] } <= { data_i[78:78] };
    end 
    if(N8454) begin
      { mem[2077:2077] } <= { data_i[77:77] };
    end 
    if(N8453) begin
      { mem[2076:2076] } <= { data_i[76:76] };
    end 
    if(N8452) begin
      { mem[2075:2075] } <= { data_i[75:75] };
    end 
    if(N8451) begin
      { mem[2074:2074] } <= { data_i[74:74] };
    end 
    if(N8450) begin
      { mem[2073:2073] } <= { data_i[73:73] };
    end 
    if(N8449) begin
      { mem[2072:2072] } <= { data_i[72:72] };
    end 
    if(N8448) begin
      { mem[2071:2071] } <= { data_i[71:71] };
    end 
    if(N8447) begin
      { mem[2070:2070] } <= { data_i[70:70] };
    end 
    if(N8446) begin
      { mem[2069:2069] } <= { data_i[69:69] };
    end 
    if(N8445) begin
      { mem[2068:2068] } <= { data_i[68:68] };
    end 
    if(N8444) begin
      { mem[2067:2067] } <= { data_i[67:67] };
    end 
    if(N8443) begin
      { mem[2066:2066] } <= { data_i[66:66] };
    end 
    if(N8442) begin
      { mem[2065:2065] } <= { data_i[65:65] };
    end 
    if(N8441) begin
      { mem[2064:2064] } <= { data_i[64:64] };
    end 
    if(N8440) begin
      { mem[2063:2063] } <= { data_i[63:63] };
    end 
    if(N8439) begin
      { mem[2062:2062] } <= { data_i[62:62] };
    end 
    if(N8438) begin
      { mem[2061:2061] } <= { data_i[61:61] };
    end 
    if(N8437) begin
      { mem[2060:2060] } <= { data_i[60:60] };
    end 
    if(N8436) begin
      { mem[2059:2059] } <= { data_i[59:59] };
    end 
    if(N8435) begin
      { mem[2058:2058] } <= { data_i[58:58] };
    end 
    if(N8434) begin
      { mem[2057:2057] } <= { data_i[57:57] };
    end 
    if(N8433) begin
      { mem[2056:2056] } <= { data_i[56:56] };
    end 
    if(N8432) begin
      { mem[2055:2055] } <= { data_i[55:55] };
    end 
    if(N8431) begin
      { mem[2054:2054] } <= { data_i[54:54] };
    end 
    if(N8430) begin
      { mem[2053:2053] } <= { data_i[53:53] };
    end 
    if(N8429) begin
      { mem[2052:2052] } <= { data_i[52:52] };
    end 
    if(N8428) begin
      { mem[2051:2051] } <= { data_i[51:51] };
    end 
    if(N8427) begin
      { mem[2050:2050] } <= { data_i[50:50] };
    end 
    if(N8426) begin
      { mem[2049:2049] } <= { data_i[49:49] };
    end 
    if(N8425) begin
      { mem[2048:2048] } <= { data_i[48:48] };
    end 
    if(N8424) begin
      { mem[2047:2047] } <= { data_i[47:47] };
    end 
    if(N8423) begin
      { mem[2046:2046] } <= { data_i[46:46] };
    end 
    if(N8422) begin
      { mem[2045:2045] } <= { data_i[45:45] };
    end 
    if(N8421) begin
      { mem[2044:2044] } <= { data_i[44:44] };
    end 
    if(N8420) begin
      { mem[2043:2043] } <= { data_i[43:43] };
    end 
    if(N8419) begin
      { mem[2042:2042] } <= { data_i[42:42] };
    end 
    if(N8418) begin
      { mem[2041:2041] } <= { data_i[41:41] };
    end 
    if(N8417) begin
      { mem[2040:2040] } <= { data_i[40:40] };
    end 
    if(N8416) begin
      { mem[2039:2039] } <= { data_i[39:39] };
    end 
    if(N8415) begin
      { mem[2038:2038] } <= { data_i[38:38] };
    end 
    if(N8414) begin
      { mem[2037:2037] } <= { data_i[37:37] };
    end 
    if(N8413) begin
      { mem[2036:2036] } <= { data_i[36:36] };
    end 
    if(N8412) begin
      { mem[2035:2035] } <= { data_i[35:35] };
    end 
    if(N8411) begin
      { mem[2034:2034] } <= { data_i[34:34] };
    end 
    if(N8410) begin
      { mem[2033:2033] } <= { data_i[33:33] };
    end 
    if(N8409) begin
      { mem[2032:2032] } <= { data_i[32:32] };
    end 
    if(N8408) begin
      { mem[2031:2031] } <= { data_i[31:31] };
    end 
    if(N8407) begin
      { mem[2030:2030] } <= { data_i[30:30] };
    end 
    if(N8406) begin
      { mem[2029:2029] } <= { data_i[29:29] };
    end 
    if(N8405) begin
      { mem[2028:2028] } <= { data_i[28:28] };
    end 
    if(N8404) begin
      { mem[2027:2027] } <= { data_i[27:27] };
    end 
    if(N8403) begin
      { mem[2026:2026] } <= { data_i[26:26] };
    end 
    if(N8402) begin
      { mem[2025:2025] } <= { data_i[25:25] };
    end 
    if(N8401) begin
      { mem[2024:2024] } <= { data_i[24:24] };
    end 
    if(N8400) begin
      { mem[2023:2023] } <= { data_i[23:23] };
    end 
    if(N8399) begin
      { mem[2022:2022] } <= { data_i[22:22] };
    end 
    if(N8398) begin
      { mem[2021:2021] } <= { data_i[21:21] };
    end 
    if(N8397) begin
      { mem[2020:2020] } <= { data_i[20:20] };
    end 
    if(N8396) begin
      { mem[2019:2019] } <= { data_i[19:19] };
    end 
    if(N8395) begin
      { mem[2018:2018] } <= { data_i[18:18] };
    end 
    if(N8394) begin
      { mem[2017:2017] } <= { data_i[17:17] };
    end 
    if(N8393) begin
      { mem[2016:2016] } <= { data_i[16:16] };
    end 
    if(N8392) begin
      { mem[2015:2015] } <= { data_i[15:15] };
    end 
    if(N8391) begin
      { mem[2014:2014] } <= { data_i[14:14] };
    end 
    if(N8390) begin
      { mem[2013:2013] } <= { data_i[13:13] };
    end 
    if(N8389) begin
      { mem[2012:2012] } <= { data_i[12:12] };
    end 
    if(N8388) begin
      { mem[2011:2011] } <= { data_i[11:11] };
    end 
    if(N8387) begin
      { mem[2010:2010] } <= { data_i[10:10] };
    end 
    if(N8386) begin
      { mem[2009:2009] } <= { data_i[9:9] };
    end 
    if(N8385) begin
      { mem[2008:2008] } <= { data_i[8:8] };
    end 
    if(N8384) begin
      { mem[2007:2007] } <= { data_i[7:7] };
    end 
    if(N8383) begin
      { mem[2006:2006] } <= { data_i[6:6] };
    end 
    if(N8382) begin
      { mem[2005:2005] } <= { data_i[5:5] };
    end 
    if(N8381) begin
      { mem[2004:2004] } <= { data_i[4:4] };
    end 
    if(N8380) begin
      { mem[2003:2003] } <= { data_i[3:3] };
    end 
    if(N8379) begin
      { mem[2002:2002] } <= { data_i[2:2] };
    end 
    if(N8378) begin
      { mem[2001:2001] } <= { data_i[1:1] };
    end 
    if(N8377) begin
      { mem[2000:2000] } <= { data_i[0:0] };
    end 
    if(N8376) begin
      { mem[1999:1999] } <= { data_i[79:79] };
    end 
    if(N8375) begin
      { mem[1998:1998] } <= { data_i[78:78] };
    end 
    if(N8374) begin
      { mem[1997:1997] } <= { data_i[77:77] };
    end 
    if(N8373) begin
      { mem[1996:1996] } <= { data_i[76:76] };
    end 
    if(N8372) begin
      { mem[1995:1995] } <= { data_i[75:75] };
    end 
    if(N8371) begin
      { mem[1994:1994] } <= { data_i[74:74] };
    end 
    if(N8370) begin
      { mem[1993:1993] } <= { data_i[73:73] };
    end 
    if(N8369) begin
      { mem[1992:1992] } <= { data_i[72:72] };
    end 
    if(N8368) begin
      { mem[1991:1991] } <= { data_i[71:71] };
    end 
    if(N8367) begin
      { mem[1990:1990] } <= { data_i[70:70] };
    end 
    if(N8366) begin
      { mem[1989:1989] } <= { data_i[69:69] };
    end 
    if(N8365) begin
      { mem[1988:1988] } <= { data_i[68:68] };
    end 
    if(N8364) begin
      { mem[1987:1987] } <= { data_i[67:67] };
    end 
    if(N8363) begin
      { mem[1986:1986] } <= { data_i[66:66] };
    end 
    if(N8362) begin
      { mem[1985:1985] } <= { data_i[65:65] };
    end 
    if(N8361) begin
      { mem[1984:1984] } <= { data_i[64:64] };
    end 
    if(N8360) begin
      { mem[1983:1983] } <= { data_i[63:63] };
    end 
    if(N8359) begin
      { mem[1982:1982] } <= { data_i[62:62] };
    end 
    if(N8358) begin
      { mem[1981:1981] } <= { data_i[61:61] };
    end 
    if(N8357) begin
      { mem[1980:1980] } <= { data_i[60:60] };
    end 
    if(N8356) begin
      { mem[1979:1979] } <= { data_i[59:59] };
    end 
    if(N8355) begin
      { mem[1978:1978] } <= { data_i[58:58] };
    end 
    if(N8354) begin
      { mem[1977:1977] } <= { data_i[57:57] };
    end 
    if(N8353) begin
      { mem[1976:1976] } <= { data_i[56:56] };
    end 
    if(N8352) begin
      { mem[1975:1975] } <= { data_i[55:55] };
    end 
    if(N8351) begin
      { mem[1974:1974] } <= { data_i[54:54] };
    end 
    if(N8350) begin
      { mem[1973:1973] } <= { data_i[53:53] };
    end 
    if(N8349) begin
      { mem[1972:1972] } <= { data_i[52:52] };
    end 
    if(N8348) begin
      { mem[1971:1971] } <= { data_i[51:51] };
    end 
    if(N8347) begin
      { mem[1970:1970] } <= { data_i[50:50] };
    end 
    if(N8346) begin
      { mem[1969:1969] } <= { data_i[49:49] };
    end 
    if(N8345) begin
      { mem[1968:1968] } <= { data_i[48:48] };
    end 
    if(N8344) begin
      { mem[1967:1967] } <= { data_i[47:47] };
    end 
    if(N8343) begin
      { mem[1966:1966] } <= { data_i[46:46] };
    end 
    if(N8342) begin
      { mem[1965:1965] } <= { data_i[45:45] };
    end 
    if(N8341) begin
      { mem[1964:1964] } <= { data_i[44:44] };
    end 
    if(N8340) begin
      { mem[1963:1963] } <= { data_i[43:43] };
    end 
    if(N8339) begin
      { mem[1962:1962] } <= { data_i[42:42] };
    end 
    if(N8338) begin
      { mem[1961:1961] } <= { data_i[41:41] };
    end 
    if(N8337) begin
      { mem[1960:1960] } <= { data_i[40:40] };
    end 
    if(N8336) begin
      { mem[1959:1959] } <= { data_i[39:39] };
    end 
    if(N8335) begin
      { mem[1958:1958] } <= { data_i[38:38] };
    end 
    if(N8334) begin
      { mem[1957:1957] } <= { data_i[37:37] };
    end 
    if(N8333) begin
      { mem[1956:1956] } <= { data_i[36:36] };
    end 
    if(N8332) begin
      { mem[1955:1955] } <= { data_i[35:35] };
    end 
    if(N8331) begin
      { mem[1954:1954] } <= { data_i[34:34] };
    end 
    if(N8330) begin
      { mem[1953:1953] } <= { data_i[33:33] };
    end 
    if(N8329) begin
      { mem[1952:1952] } <= { data_i[32:32] };
    end 
    if(N8328) begin
      { mem[1951:1951] } <= { data_i[31:31] };
    end 
    if(N8327) begin
      { mem[1950:1950] } <= { data_i[30:30] };
    end 
    if(N8326) begin
      { mem[1949:1949] } <= { data_i[29:29] };
    end 
    if(N8325) begin
      { mem[1948:1948] } <= { data_i[28:28] };
    end 
    if(N8324) begin
      { mem[1947:1947] } <= { data_i[27:27] };
    end 
    if(N8323) begin
      { mem[1946:1946] } <= { data_i[26:26] };
    end 
    if(N8322) begin
      { mem[1945:1945] } <= { data_i[25:25] };
    end 
    if(N8321) begin
      { mem[1944:1944] } <= { data_i[24:24] };
    end 
    if(N8320) begin
      { mem[1943:1943] } <= { data_i[23:23] };
    end 
    if(N8319) begin
      { mem[1942:1942] } <= { data_i[22:22] };
    end 
    if(N8318) begin
      { mem[1941:1941] } <= { data_i[21:21] };
    end 
    if(N8317) begin
      { mem[1940:1940] } <= { data_i[20:20] };
    end 
    if(N8316) begin
      { mem[1939:1939] } <= { data_i[19:19] };
    end 
    if(N8315) begin
      { mem[1938:1938] } <= { data_i[18:18] };
    end 
    if(N8314) begin
      { mem[1937:1937] } <= { data_i[17:17] };
    end 
    if(N8313) begin
      { mem[1936:1936] } <= { data_i[16:16] };
    end 
    if(N8312) begin
      { mem[1935:1935] } <= { data_i[15:15] };
    end 
    if(N8311) begin
      { mem[1934:1934] } <= { data_i[14:14] };
    end 
    if(N8310) begin
      { mem[1933:1933] } <= { data_i[13:13] };
    end 
    if(N8309) begin
      { mem[1932:1932] } <= { data_i[12:12] };
    end 
    if(N8308) begin
      { mem[1931:1931] } <= { data_i[11:11] };
    end 
    if(N8307) begin
      { mem[1930:1930] } <= { data_i[10:10] };
    end 
    if(N8306) begin
      { mem[1929:1929] } <= { data_i[9:9] };
    end 
    if(N8305) begin
      { mem[1928:1928] } <= { data_i[8:8] };
    end 
    if(N8304) begin
      { mem[1927:1927] } <= { data_i[7:7] };
    end 
    if(N8303) begin
      { mem[1926:1926] } <= { data_i[6:6] };
    end 
    if(N8302) begin
      { mem[1925:1925] } <= { data_i[5:5] };
    end 
    if(N8301) begin
      { mem[1924:1924] } <= { data_i[4:4] };
    end 
    if(N8300) begin
      { mem[1923:1923] } <= { data_i[3:3] };
    end 
    if(N8299) begin
      { mem[1922:1922] } <= { data_i[2:2] };
    end 
    if(N8298) begin
      { mem[1921:1921] } <= { data_i[1:1] };
    end 
    if(N8297) begin
      { mem[1920:1920] } <= { data_i[0:0] };
    end 
    if(N8296) begin
      { mem[1919:1919] } <= { data_i[79:79] };
    end 
    if(N8295) begin
      { mem[1918:1918] } <= { data_i[78:78] };
    end 
    if(N8294) begin
      { mem[1917:1917] } <= { data_i[77:77] };
    end 
    if(N8293) begin
      { mem[1916:1916] } <= { data_i[76:76] };
    end 
    if(N8292) begin
      { mem[1915:1915] } <= { data_i[75:75] };
    end 
    if(N8291) begin
      { mem[1914:1914] } <= { data_i[74:74] };
    end 
    if(N8290) begin
      { mem[1913:1913] } <= { data_i[73:73] };
    end 
    if(N8289) begin
      { mem[1912:1912] } <= { data_i[72:72] };
    end 
    if(N8288) begin
      { mem[1911:1911] } <= { data_i[71:71] };
    end 
    if(N8287) begin
      { mem[1910:1910] } <= { data_i[70:70] };
    end 
    if(N8286) begin
      { mem[1909:1909] } <= { data_i[69:69] };
    end 
    if(N8285) begin
      { mem[1908:1908] } <= { data_i[68:68] };
    end 
    if(N8284) begin
      { mem[1907:1907] } <= { data_i[67:67] };
    end 
    if(N8283) begin
      { mem[1906:1906] } <= { data_i[66:66] };
    end 
    if(N8282) begin
      { mem[1905:1905] } <= { data_i[65:65] };
    end 
    if(N8281) begin
      { mem[1904:1904] } <= { data_i[64:64] };
    end 
    if(N8280) begin
      { mem[1903:1903] } <= { data_i[63:63] };
    end 
    if(N8279) begin
      { mem[1902:1902] } <= { data_i[62:62] };
    end 
    if(N8278) begin
      { mem[1901:1901] } <= { data_i[61:61] };
    end 
    if(N8277) begin
      { mem[1900:1900] } <= { data_i[60:60] };
    end 
    if(N8276) begin
      { mem[1899:1899] } <= { data_i[59:59] };
    end 
    if(N8275) begin
      { mem[1898:1898] } <= { data_i[58:58] };
    end 
    if(N8274) begin
      { mem[1897:1897] } <= { data_i[57:57] };
    end 
    if(N8273) begin
      { mem[1896:1896] } <= { data_i[56:56] };
    end 
    if(N8272) begin
      { mem[1895:1895] } <= { data_i[55:55] };
    end 
    if(N8271) begin
      { mem[1894:1894] } <= { data_i[54:54] };
    end 
    if(N8270) begin
      { mem[1893:1893] } <= { data_i[53:53] };
    end 
    if(N8269) begin
      { mem[1892:1892] } <= { data_i[52:52] };
    end 
    if(N8268) begin
      { mem[1891:1891] } <= { data_i[51:51] };
    end 
    if(N8267) begin
      { mem[1890:1890] } <= { data_i[50:50] };
    end 
    if(N8266) begin
      { mem[1889:1889] } <= { data_i[49:49] };
    end 
    if(N8265) begin
      { mem[1888:1888] } <= { data_i[48:48] };
    end 
    if(N8264) begin
      { mem[1887:1887] } <= { data_i[47:47] };
    end 
    if(N8263) begin
      { mem[1886:1886] } <= { data_i[46:46] };
    end 
    if(N8262) begin
      { mem[1885:1885] } <= { data_i[45:45] };
    end 
    if(N8261) begin
      { mem[1884:1884] } <= { data_i[44:44] };
    end 
    if(N8260) begin
      { mem[1883:1883] } <= { data_i[43:43] };
    end 
    if(N8259) begin
      { mem[1882:1882] } <= { data_i[42:42] };
    end 
    if(N8258) begin
      { mem[1881:1881] } <= { data_i[41:41] };
    end 
    if(N8257) begin
      { mem[1880:1880] } <= { data_i[40:40] };
    end 
    if(N8256) begin
      { mem[1879:1879] } <= { data_i[39:39] };
    end 
    if(N8255) begin
      { mem[1878:1878] } <= { data_i[38:38] };
    end 
    if(N8254) begin
      { mem[1877:1877] } <= { data_i[37:37] };
    end 
    if(N8253) begin
      { mem[1876:1876] } <= { data_i[36:36] };
    end 
    if(N8252) begin
      { mem[1875:1875] } <= { data_i[35:35] };
    end 
    if(N8251) begin
      { mem[1874:1874] } <= { data_i[34:34] };
    end 
    if(N8250) begin
      { mem[1873:1873] } <= { data_i[33:33] };
    end 
    if(N8249) begin
      { mem[1872:1872] } <= { data_i[32:32] };
    end 
    if(N8248) begin
      { mem[1871:1871] } <= { data_i[31:31] };
    end 
    if(N8247) begin
      { mem[1870:1870] } <= { data_i[30:30] };
    end 
    if(N8246) begin
      { mem[1869:1869] } <= { data_i[29:29] };
    end 
    if(N8245) begin
      { mem[1868:1868] } <= { data_i[28:28] };
    end 
    if(N8244) begin
      { mem[1867:1867] } <= { data_i[27:27] };
    end 
    if(N8243) begin
      { mem[1866:1866] } <= { data_i[26:26] };
    end 
    if(N8242) begin
      { mem[1865:1865] } <= { data_i[25:25] };
    end 
    if(N8241) begin
      { mem[1864:1864] } <= { data_i[24:24] };
    end 
    if(N8240) begin
      { mem[1863:1863] } <= { data_i[23:23] };
    end 
    if(N8239) begin
      { mem[1862:1862] } <= { data_i[22:22] };
    end 
    if(N8238) begin
      { mem[1861:1861] } <= { data_i[21:21] };
    end 
    if(N8237) begin
      { mem[1860:1860] } <= { data_i[20:20] };
    end 
    if(N8236) begin
      { mem[1859:1859] } <= { data_i[19:19] };
    end 
    if(N8235) begin
      { mem[1858:1858] } <= { data_i[18:18] };
    end 
    if(N8234) begin
      { mem[1857:1857] } <= { data_i[17:17] };
    end 
    if(N8233) begin
      { mem[1856:1856] } <= { data_i[16:16] };
    end 
    if(N8232) begin
      { mem[1855:1855] } <= { data_i[15:15] };
    end 
    if(N8231) begin
      { mem[1854:1854] } <= { data_i[14:14] };
    end 
    if(N8230) begin
      { mem[1853:1853] } <= { data_i[13:13] };
    end 
    if(N8229) begin
      { mem[1852:1852] } <= { data_i[12:12] };
    end 
    if(N8228) begin
      { mem[1851:1851] } <= { data_i[11:11] };
    end 
    if(N8227) begin
      { mem[1850:1850] } <= { data_i[10:10] };
    end 
    if(N8226) begin
      { mem[1849:1849] } <= { data_i[9:9] };
    end 
    if(N8225) begin
      { mem[1848:1848] } <= { data_i[8:8] };
    end 
    if(N8224) begin
      { mem[1847:1847] } <= { data_i[7:7] };
    end 
    if(N8223) begin
      { mem[1846:1846] } <= { data_i[6:6] };
    end 
    if(N8222) begin
      { mem[1845:1845] } <= { data_i[5:5] };
    end 
    if(N8221) begin
      { mem[1844:1844] } <= { data_i[4:4] };
    end 
    if(N8220) begin
      { mem[1843:1843] } <= { data_i[3:3] };
    end 
    if(N8219) begin
      { mem[1842:1842] } <= { data_i[2:2] };
    end 
    if(N8218) begin
      { mem[1841:1841] } <= { data_i[1:1] };
    end 
    if(N8217) begin
      { mem[1840:1840] } <= { data_i[0:0] };
    end 
    if(N8216) begin
      { mem[1839:1839] } <= { data_i[79:79] };
    end 
    if(N8215) begin
      { mem[1838:1838] } <= { data_i[78:78] };
    end 
    if(N8214) begin
      { mem[1837:1837] } <= { data_i[77:77] };
    end 
    if(N8213) begin
      { mem[1836:1836] } <= { data_i[76:76] };
    end 
    if(N8212) begin
      { mem[1835:1835] } <= { data_i[75:75] };
    end 
    if(N8211) begin
      { mem[1834:1834] } <= { data_i[74:74] };
    end 
    if(N8210) begin
      { mem[1833:1833] } <= { data_i[73:73] };
    end 
    if(N8209) begin
      { mem[1832:1832] } <= { data_i[72:72] };
    end 
    if(N8208) begin
      { mem[1831:1831] } <= { data_i[71:71] };
    end 
    if(N8207) begin
      { mem[1830:1830] } <= { data_i[70:70] };
    end 
    if(N8206) begin
      { mem[1829:1829] } <= { data_i[69:69] };
    end 
    if(N8205) begin
      { mem[1828:1828] } <= { data_i[68:68] };
    end 
    if(N8204) begin
      { mem[1827:1827] } <= { data_i[67:67] };
    end 
    if(N8203) begin
      { mem[1826:1826] } <= { data_i[66:66] };
    end 
    if(N8202) begin
      { mem[1825:1825] } <= { data_i[65:65] };
    end 
    if(N8201) begin
      { mem[1824:1824] } <= { data_i[64:64] };
    end 
    if(N8200) begin
      { mem[1823:1823] } <= { data_i[63:63] };
    end 
    if(N8199) begin
      { mem[1822:1822] } <= { data_i[62:62] };
    end 
    if(N8198) begin
      { mem[1821:1821] } <= { data_i[61:61] };
    end 
    if(N8197) begin
      { mem[1820:1820] } <= { data_i[60:60] };
    end 
    if(N8196) begin
      { mem[1819:1819] } <= { data_i[59:59] };
    end 
    if(N8195) begin
      { mem[1818:1818] } <= { data_i[58:58] };
    end 
    if(N8194) begin
      { mem[1817:1817] } <= { data_i[57:57] };
    end 
    if(N8193) begin
      { mem[1816:1816] } <= { data_i[56:56] };
    end 
    if(N8192) begin
      { mem[1815:1815] } <= { data_i[55:55] };
    end 
    if(N8191) begin
      { mem[1814:1814] } <= { data_i[54:54] };
    end 
    if(N8190) begin
      { mem[1813:1813] } <= { data_i[53:53] };
    end 
    if(N8189) begin
      { mem[1812:1812] } <= { data_i[52:52] };
    end 
    if(N8188) begin
      { mem[1811:1811] } <= { data_i[51:51] };
    end 
    if(N8187) begin
      { mem[1810:1810] } <= { data_i[50:50] };
    end 
    if(N8186) begin
      { mem[1809:1809] } <= { data_i[49:49] };
    end 
    if(N8185) begin
      { mem[1808:1808] } <= { data_i[48:48] };
    end 
    if(N8184) begin
      { mem[1807:1807] } <= { data_i[47:47] };
    end 
    if(N8183) begin
      { mem[1806:1806] } <= { data_i[46:46] };
    end 
    if(N8182) begin
      { mem[1805:1805] } <= { data_i[45:45] };
    end 
    if(N8181) begin
      { mem[1804:1804] } <= { data_i[44:44] };
    end 
    if(N8180) begin
      { mem[1803:1803] } <= { data_i[43:43] };
    end 
    if(N8179) begin
      { mem[1802:1802] } <= { data_i[42:42] };
    end 
    if(N8178) begin
      { mem[1801:1801] } <= { data_i[41:41] };
    end 
    if(N8177) begin
      { mem[1800:1800] } <= { data_i[40:40] };
    end 
    if(N8176) begin
      { mem[1799:1799] } <= { data_i[39:39] };
    end 
    if(N8175) begin
      { mem[1798:1798] } <= { data_i[38:38] };
    end 
    if(N8174) begin
      { mem[1797:1797] } <= { data_i[37:37] };
    end 
    if(N8173) begin
      { mem[1796:1796] } <= { data_i[36:36] };
    end 
    if(N8172) begin
      { mem[1795:1795] } <= { data_i[35:35] };
    end 
    if(N8171) begin
      { mem[1794:1794] } <= { data_i[34:34] };
    end 
    if(N8170) begin
      { mem[1793:1793] } <= { data_i[33:33] };
    end 
    if(N8169) begin
      { mem[1792:1792] } <= { data_i[32:32] };
    end 
    if(N8168) begin
      { mem[1791:1791] } <= { data_i[31:31] };
    end 
    if(N8167) begin
      { mem[1790:1790] } <= { data_i[30:30] };
    end 
    if(N8166) begin
      { mem[1789:1789] } <= { data_i[29:29] };
    end 
    if(N8165) begin
      { mem[1788:1788] } <= { data_i[28:28] };
    end 
    if(N8164) begin
      { mem[1787:1787] } <= { data_i[27:27] };
    end 
    if(N8163) begin
      { mem[1786:1786] } <= { data_i[26:26] };
    end 
    if(N8162) begin
      { mem[1785:1785] } <= { data_i[25:25] };
    end 
    if(N8161) begin
      { mem[1784:1784] } <= { data_i[24:24] };
    end 
    if(N8160) begin
      { mem[1783:1783] } <= { data_i[23:23] };
    end 
    if(N8159) begin
      { mem[1782:1782] } <= { data_i[22:22] };
    end 
    if(N8158) begin
      { mem[1781:1781] } <= { data_i[21:21] };
    end 
    if(N8157) begin
      { mem[1780:1780] } <= { data_i[20:20] };
    end 
    if(N8156) begin
      { mem[1779:1779] } <= { data_i[19:19] };
    end 
    if(N8155) begin
      { mem[1778:1778] } <= { data_i[18:18] };
    end 
    if(N8154) begin
      { mem[1777:1777] } <= { data_i[17:17] };
    end 
    if(N8153) begin
      { mem[1776:1776] } <= { data_i[16:16] };
    end 
    if(N8152) begin
      { mem[1775:1775] } <= { data_i[15:15] };
    end 
    if(N8151) begin
      { mem[1774:1774] } <= { data_i[14:14] };
    end 
    if(N8150) begin
      { mem[1773:1773] } <= { data_i[13:13] };
    end 
    if(N8149) begin
      { mem[1772:1772] } <= { data_i[12:12] };
    end 
    if(N8148) begin
      { mem[1771:1771] } <= { data_i[11:11] };
    end 
    if(N8147) begin
      { mem[1770:1770] } <= { data_i[10:10] };
    end 
    if(N8146) begin
      { mem[1769:1769] } <= { data_i[9:9] };
    end 
    if(N8145) begin
      { mem[1768:1768] } <= { data_i[8:8] };
    end 
    if(N8144) begin
      { mem[1767:1767] } <= { data_i[7:7] };
    end 
    if(N8143) begin
      { mem[1766:1766] } <= { data_i[6:6] };
    end 
    if(N8142) begin
      { mem[1765:1765] } <= { data_i[5:5] };
    end 
    if(N8141) begin
      { mem[1764:1764] } <= { data_i[4:4] };
    end 
    if(N8140) begin
      { mem[1763:1763] } <= { data_i[3:3] };
    end 
    if(N8139) begin
      { mem[1762:1762] } <= { data_i[2:2] };
    end 
    if(N8138) begin
      { mem[1761:1761] } <= { data_i[1:1] };
    end 
    if(N8137) begin
      { mem[1760:1760] } <= { data_i[0:0] };
    end 
    if(N8136) begin
      { mem[1759:1759] } <= { data_i[79:79] };
    end 
    if(N8135) begin
      { mem[1758:1758] } <= { data_i[78:78] };
    end 
    if(N8134) begin
      { mem[1757:1757] } <= { data_i[77:77] };
    end 
    if(N8133) begin
      { mem[1756:1756] } <= { data_i[76:76] };
    end 
    if(N8132) begin
      { mem[1755:1755] } <= { data_i[75:75] };
    end 
    if(N8131) begin
      { mem[1754:1754] } <= { data_i[74:74] };
    end 
    if(N8130) begin
      { mem[1753:1753] } <= { data_i[73:73] };
    end 
    if(N8129) begin
      { mem[1752:1752] } <= { data_i[72:72] };
    end 
    if(N8128) begin
      { mem[1751:1751] } <= { data_i[71:71] };
    end 
    if(N8127) begin
      { mem[1750:1750] } <= { data_i[70:70] };
    end 
    if(N8126) begin
      { mem[1749:1749] } <= { data_i[69:69] };
    end 
    if(N8125) begin
      { mem[1748:1748] } <= { data_i[68:68] };
    end 
    if(N8124) begin
      { mem[1747:1747] } <= { data_i[67:67] };
    end 
    if(N8123) begin
      { mem[1746:1746] } <= { data_i[66:66] };
    end 
    if(N8122) begin
      { mem[1745:1745] } <= { data_i[65:65] };
    end 
    if(N8121) begin
      { mem[1744:1744] } <= { data_i[64:64] };
    end 
    if(N8120) begin
      { mem[1743:1743] } <= { data_i[63:63] };
    end 
    if(N8119) begin
      { mem[1742:1742] } <= { data_i[62:62] };
    end 
    if(N8118) begin
      { mem[1741:1741] } <= { data_i[61:61] };
    end 
    if(N8117) begin
      { mem[1740:1740] } <= { data_i[60:60] };
    end 
    if(N8116) begin
      { mem[1739:1739] } <= { data_i[59:59] };
    end 
    if(N8115) begin
      { mem[1738:1738] } <= { data_i[58:58] };
    end 
    if(N8114) begin
      { mem[1737:1737] } <= { data_i[57:57] };
    end 
    if(N8113) begin
      { mem[1736:1736] } <= { data_i[56:56] };
    end 
    if(N8112) begin
      { mem[1735:1735] } <= { data_i[55:55] };
    end 
    if(N8111) begin
      { mem[1734:1734] } <= { data_i[54:54] };
    end 
    if(N8110) begin
      { mem[1733:1733] } <= { data_i[53:53] };
    end 
    if(N8109) begin
      { mem[1732:1732] } <= { data_i[52:52] };
    end 
    if(N8108) begin
      { mem[1731:1731] } <= { data_i[51:51] };
    end 
    if(N8107) begin
      { mem[1730:1730] } <= { data_i[50:50] };
    end 
    if(N8106) begin
      { mem[1729:1729] } <= { data_i[49:49] };
    end 
    if(N8105) begin
      { mem[1728:1728] } <= { data_i[48:48] };
    end 
    if(N8104) begin
      { mem[1727:1727] } <= { data_i[47:47] };
    end 
    if(N8103) begin
      { mem[1726:1726] } <= { data_i[46:46] };
    end 
    if(N8102) begin
      { mem[1725:1725] } <= { data_i[45:45] };
    end 
    if(N8101) begin
      { mem[1724:1724] } <= { data_i[44:44] };
    end 
    if(N8100) begin
      { mem[1723:1723] } <= { data_i[43:43] };
    end 
    if(N8099) begin
      { mem[1722:1722] } <= { data_i[42:42] };
    end 
    if(N8098) begin
      { mem[1721:1721] } <= { data_i[41:41] };
    end 
    if(N8097) begin
      { mem[1720:1720] } <= { data_i[40:40] };
    end 
    if(N8096) begin
      { mem[1719:1719] } <= { data_i[39:39] };
    end 
    if(N8095) begin
      { mem[1718:1718] } <= { data_i[38:38] };
    end 
    if(N8094) begin
      { mem[1717:1717] } <= { data_i[37:37] };
    end 
    if(N8093) begin
      { mem[1716:1716] } <= { data_i[36:36] };
    end 
    if(N8092) begin
      { mem[1715:1715] } <= { data_i[35:35] };
    end 
    if(N8091) begin
      { mem[1714:1714] } <= { data_i[34:34] };
    end 
    if(N8090) begin
      { mem[1713:1713] } <= { data_i[33:33] };
    end 
    if(N8089) begin
      { mem[1712:1712] } <= { data_i[32:32] };
    end 
    if(N8088) begin
      { mem[1711:1711] } <= { data_i[31:31] };
    end 
    if(N8087) begin
      { mem[1710:1710] } <= { data_i[30:30] };
    end 
    if(N8086) begin
      { mem[1709:1709] } <= { data_i[29:29] };
    end 
    if(N8085) begin
      { mem[1708:1708] } <= { data_i[28:28] };
    end 
    if(N8084) begin
      { mem[1707:1707] } <= { data_i[27:27] };
    end 
    if(N8083) begin
      { mem[1706:1706] } <= { data_i[26:26] };
    end 
    if(N8082) begin
      { mem[1705:1705] } <= { data_i[25:25] };
    end 
    if(N8081) begin
      { mem[1704:1704] } <= { data_i[24:24] };
    end 
    if(N8080) begin
      { mem[1703:1703] } <= { data_i[23:23] };
    end 
    if(N8079) begin
      { mem[1702:1702] } <= { data_i[22:22] };
    end 
    if(N8078) begin
      { mem[1701:1701] } <= { data_i[21:21] };
    end 
    if(N8077) begin
      { mem[1700:1700] } <= { data_i[20:20] };
    end 
    if(N8076) begin
      { mem[1699:1699] } <= { data_i[19:19] };
    end 
    if(N8075) begin
      { mem[1698:1698] } <= { data_i[18:18] };
    end 
    if(N8074) begin
      { mem[1697:1697] } <= { data_i[17:17] };
    end 
    if(N8073) begin
      { mem[1696:1696] } <= { data_i[16:16] };
    end 
    if(N8072) begin
      { mem[1695:1695] } <= { data_i[15:15] };
    end 
    if(N8071) begin
      { mem[1694:1694] } <= { data_i[14:14] };
    end 
    if(N8070) begin
      { mem[1693:1693] } <= { data_i[13:13] };
    end 
    if(N8069) begin
      { mem[1692:1692] } <= { data_i[12:12] };
    end 
    if(N8068) begin
      { mem[1691:1691] } <= { data_i[11:11] };
    end 
    if(N8067) begin
      { mem[1690:1690] } <= { data_i[10:10] };
    end 
    if(N8066) begin
      { mem[1689:1689] } <= { data_i[9:9] };
    end 
    if(N8065) begin
      { mem[1688:1688] } <= { data_i[8:8] };
    end 
    if(N8064) begin
      { mem[1687:1687] } <= { data_i[7:7] };
    end 
    if(N8063) begin
      { mem[1686:1686] } <= { data_i[6:6] };
    end 
    if(N8062) begin
      { mem[1685:1685] } <= { data_i[5:5] };
    end 
    if(N8061) begin
      { mem[1684:1684] } <= { data_i[4:4] };
    end 
    if(N8060) begin
      { mem[1683:1683] } <= { data_i[3:3] };
    end 
    if(N8059) begin
      { mem[1682:1682] } <= { data_i[2:2] };
    end 
    if(N8058) begin
      { mem[1681:1681] } <= { data_i[1:1] };
    end 
    if(N8057) begin
      { mem[1680:1680] } <= { data_i[0:0] };
    end 
    if(N8056) begin
      { mem[1679:1679] } <= { data_i[79:79] };
    end 
    if(N8055) begin
      { mem[1678:1678] } <= { data_i[78:78] };
    end 
    if(N8054) begin
      { mem[1677:1677] } <= { data_i[77:77] };
    end 
    if(N8053) begin
      { mem[1676:1676] } <= { data_i[76:76] };
    end 
    if(N8052) begin
      { mem[1675:1675] } <= { data_i[75:75] };
    end 
    if(N8051) begin
      { mem[1674:1674] } <= { data_i[74:74] };
    end 
    if(N8050) begin
      { mem[1673:1673] } <= { data_i[73:73] };
    end 
    if(N8049) begin
      { mem[1672:1672] } <= { data_i[72:72] };
    end 
    if(N8048) begin
      { mem[1671:1671] } <= { data_i[71:71] };
    end 
    if(N8047) begin
      { mem[1670:1670] } <= { data_i[70:70] };
    end 
    if(N8046) begin
      { mem[1669:1669] } <= { data_i[69:69] };
    end 
    if(N8045) begin
      { mem[1668:1668] } <= { data_i[68:68] };
    end 
    if(N8044) begin
      { mem[1667:1667] } <= { data_i[67:67] };
    end 
    if(N8043) begin
      { mem[1666:1666] } <= { data_i[66:66] };
    end 
    if(N8042) begin
      { mem[1665:1665] } <= { data_i[65:65] };
    end 
    if(N8041) begin
      { mem[1664:1664] } <= { data_i[64:64] };
    end 
    if(N8040) begin
      { mem[1663:1663] } <= { data_i[63:63] };
    end 
    if(N8039) begin
      { mem[1662:1662] } <= { data_i[62:62] };
    end 
    if(N8038) begin
      { mem[1661:1661] } <= { data_i[61:61] };
    end 
    if(N8037) begin
      { mem[1660:1660] } <= { data_i[60:60] };
    end 
    if(N8036) begin
      { mem[1659:1659] } <= { data_i[59:59] };
    end 
    if(N8035) begin
      { mem[1658:1658] } <= { data_i[58:58] };
    end 
    if(N8034) begin
      { mem[1657:1657] } <= { data_i[57:57] };
    end 
    if(N8033) begin
      { mem[1656:1656] } <= { data_i[56:56] };
    end 
    if(N8032) begin
      { mem[1655:1655] } <= { data_i[55:55] };
    end 
    if(N8031) begin
      { mem[1654:1654] } <= { data_i[54:54] };
    end 
    if(N8030) begin
      { mem[1653:1653] } <= { data_i[53:53] };
    end 
    if(N8029) begin
      { mem[1652:1652] } <= { data_i[52:52] };
    end 
    if(N8028) begin
      { mem[1651:1651] } <= { data_i[51:51] };
    end 
    if(N8027) begin
      { mem[1650:1650] } <= { data_i[50:50] };
    end 
    if(N8026) begin
      { mem[1649:1649] } <= { data_i[49:49] };
    end 
    if(N8025) begin
      { mem[1648:1648] } <= { data_i[48:48] };
    end 
    if(N8024) begin
      { mem[1647:1647] } <= { data_i[47:47] };
    end 
    if(N8023) begin
      { mem[1646:1646] } <= { data_i[46:46] };
    end 
    if(N8022) begin
      { mem[1645:1645] } <= { data_i[45:45] };
    end 
    if(N8021) begin
      { mem[1644:1644] } <= { data_i[44:44] };
    end 
    if(N8020) begin
      { mem[1643:1643] } <= { data_i[43:43] };
    end 
    if(N8019) begin
      { mem[1642:1642] } <= { data_i[42:42] };
    end 
    if(N8018) begin
      { mem[1641:1641] } <= { data_i[41:41] };
    end 
    if(N8017) begin
      { mem[1640:1640] } <= { data_i[40:40] };
    end 
    if(N8016) begin
      { mem[1639:1639] } <= { data_i[39:39] };
    end 
    if(N8015) begin
      { mem[1638:1638] } <= { data_i[38:38] };
    end 
    if(N8014) begin
      { mem[1637:1637] } <= { data_i[37:37] };
    end 
    if(N8013) begin
      { mem[1636:1636] } <= { data_i[36:36] };
    end 
    if(N8012) begin
      { mem[1635:1635] } <= { data_i[35:35] };
    end 
    if(N8011) begin
      { mem[1634:1634] } <= { data_i[34:34] };
    end 
    if(N8010) begin
      { mem[1633:1633] } <= { data_i[33:33] };
    end 
    if(N8009) begin
      { mem[1632:1632] } <= { data_i[32:32] };
    end 
    if(N8008) begin
      { mem[1631:1631] } <= { data_i[31:31] };
    end 
    if(N8007) begin
      { mem[1630:1630] } <= { data_i[30:30] };
    end 
    if(N8006) begin
      { mem[1629:1629] } <= { data_i[29:29] };
    end 
    if(N8005) begin
      { mem[1628:1628] } <= { data_i[28:28] };
    end 
    if(N8004) begin
      { mem[1627:1627] } <= { data_i[27:27] };
    end 
    if(N8003) begin
      { mem[1626:1626] } <= { data_i[26:26] };
    end 
    if(N8002) begin
      { mem[1625:1625] } <= { data_i[25:25] };
    end 
    if(N8001) begin
      { mem[1624:1624] } <= { data_i[24:24] };
    end 
    if(N8000) begin
      { mem[1623:1623] } <= { data_i[23:23] };
    end 
    if(N7999) begin
      { mem[1622:1622] } <= { data_i[22:22] };
    end 
    if(N7998) begin
      { mem[1621:1621] } <= { data_i[21:21] };
    end 
    if(N7997) begin
      { mem[1620:1620] } <= { data_i[20:20] };
    end 
    if(N7996) begin
      { mem[1619:1619] } <= { data_i[19:19] };
    end 
    if(N7995) begin
      { mem[1618:1618] } <= { data_i[18:18] };
    end 
    if(N7994) begin
      { mem[1617:1617] } <= { data_i[17:17] };
    end 
    if(N7993) begin
      { mem[1616:1616] } <= { data_i[16:16] };
    end 
    if(N7992) begin
      { mem[1615:1615] } <= { data_i[15:15] };
    end 
    if(N7991) begin
      { mem[1614:1614] } <= { data_i[14:14] };
    end 
    if(N7990) begin
      { mem[1613:1613] } <= { data_i[13:13] };
    end 
    if(N7989) begin
      { mem[1612:1612] } <= { data_i[12:12] };
    end 
    if(N7988) begin
      { mem[1611:1611] } <= { data_i[11:11] };
    end 
    if(N7987) begin
      { mem[1610:1610] } <= { data_i[10:10] };
    end 
    if(N7986) begin
      { mem[1609:1609] } <= { data_i[9:9] };
    end 
    if(N7985) begin
      { mem[1608:1608] } <= { data_i[8:8] };
    end 
    if(N7984) begin
      { mem[1607:1607] } <= { data_i[7:7] };
    end 
    if(N7983) begin
      { mem[1606:1606] } <= { data_i[6:6] };
    end 
    if(N7982) begin
      { mem[1605:1605] } <= { data_i[5:5] };
    end 
    if(N7981) begin
      { mem[1604:1604] } <= { data_i[4:4] };
    end 
    if(N7980) begin
      { mem[1603:1603] } <= { data_i[3:3] };
    end 
    if(N7979) begin
      { mem[1602:1602] } <= { data_i[2:2] };
    end 
    if(N7978) begin
      { mem[1601:1601] } <= { data_i[1:1] };
    end 
    if(N7977) begin
      { mem[1600:1600] } <= { data_i[0:0] };
    end 
    if(N7976) begin
      { mem[1599:1599] } <= { data_i[79:79] };
    end 
    if(N7975) begin
      { mem[1598:1598] } <= { data_i[78:78] };
    end 
    if(N7974) begin
      { mem[1597:1597] } <= { data_i[77:77] };
    end 
    if(N7973) begin
      { mem[1596:1596] } <= { data_i[76:76] };
    end 
    if(N7972) begin
      { mem[1595:1595] } <= { data_i[75:75] };
    end 
    if(N7971) begin
      { mem[1594:1594] } <= { data_i[74:74] };
    end 
    if(N7970) begin
      { mem[1593:1593] } <= { data_i[73:73] };
    end 
    if(N7969) begin
      { mem[1592:1592] } <= { data_i[72:72] };
    end 
    if(N7968) begin
      { mem[1591:1591] } <= { data_i[71:71] };
    end 
    if(N7967) begin
      { mem[1590:1590] } <= { data_i[70:70] };
    end 
    if(N7966) begin
      { mem[1589:1589] } <= { data_i[69:69] };
    end 
    if(N7965) begin
      { mem[1588:1588] } <= { data_i[68:68] };
    end 
    if(N7964) begin
      { mem[1587:1587] } <= { data_i[67:67] };
    end 
    if(N7963) begin
      { mem[1586:1586] } <= { data_i[66:66] };
    end 
    if(N7962) begin
      { mem[1585:1585] } <= { data_i[65:65] };
    end 
    if(N7961) begin
      { mem[1584:1584] } <= { data_i[64:64] };
    end 
    if(N7960) begin
      { mem[1583:1583] } <= { data_i[63:63] };
    end 
    if(N7959) begin
      { mem[1582:1582] } <= { data_i[62:62] };
    end 
    if(N7958) begin
      { mem[1581:1581] } <= { data_i[61:61] };
    end 
    if(N7957) begin
      { mem[1580:1580] } <= { data_i[60:60] };
    end 
    if(N7956) begin
      { mem[1579:1579] } <= { data_i[59:59] };
    end 
    if(N7955) begin
      { mem[1578:1578] } <= { data_i[58:58] };
    end 
    if(N7954) begin
      { mem[1577:1577] } <= { data_i[57:57] };
    end 
    if(N7953) begin
      { mem[1576:1576] } <= { data_i[56:56] };
    end 
    if(N7952) begin
      { mem[1575:1575] } <= { data_i[55:55] };
    end 
    if(N7951) begin
      { mem[1574:1574] } <= { data_i[54:54] };
    end 
    if(N7950) begin
      { mem[1573:1573] } <= { data_i[53:53] };
    end 
    if(N7949) begin
      { mem[1572:1572] } <= { data_i[52:52] };
    end 
    if(N7948) begin
      { mem[1571:1571] } <= { data_i[51:51] };
    end 
    if(N7947) begin
      { mem[1570:1570] } <= { data_i[50:50] };
    end 
    if(N7946) begin
      { mem[1569:1569] } <= { data_i[49:49] };
    end 
    if(N7945) begin
      { mem[1568:1568] } <= { data_i[48:48] };
    end 
    if(N7944) begin
      { mem[1567:1567] } <= { data_i[47:47] };
    end 
    if(N7943) begin
      { mem[1566:1566] } <= { data_i[46:46] };
    end 
    if(N7942) begin
      { mem[1565:1565] } <= { data_i[45:45] };
    end 
    if(N7941) begin
      { mem[1564:1564] } <= { data_i[44:44] };
    end 
    if(N7940) begin
      { mem[1563:1563] } <= { data_i[43:43] };
    end 
    if(N7939) begin
      { mem[1562:1562] } <= { data_i[42:42] };
    end 
    if(N7938) begin
      { mem[1561:1561] } <= { data_i[41:41] };
    end 
    if(N7937) begin
      { mem[1560:1560] } <= { data_i[40:40] };
    end 
    if(N7936) begin
      { mem[1559:1559] } <= { data_i[39:39] };
    end 
    if(N7935) begin
      { mem[1558:1558] } <= { data_i[38:38] };
    end 
    if(N7934) begin
      { mem[1557:1557] } <= { data_i[37:37] };
    end 
    if(N7933) begin
      { mem[1556:1556] } <= { data_i[36:36] };
    end 
    if(N7932) begin
      { mem[1555:1555] } <= { data_i[35:35] };
    end 
    if(N7931) begin
      { mem[1554:1554] } <= { data_i[34:34] };
    end 
    if(N7930) begin
      { mem[1553:1553] } <= { data_i[33:33] };
    end 
    if(N7929) begin
      { mem[1552:1552] } <= { data_i[32:32] };
    end 
    if(N7928) begin
      { mem[1551:1551] } <= { data_i[31:31] };
    end 
    if(N7927) begin
      { mem[1550:1550] } <= { data_i[30:30] };
    end 
    if(N7926) begin
      { mem[1549:1549] } <= { data_i[29:29] };
    end 
    if(N7925) begin
      { mem[1548:1548] } <= { data_i[28:28] };
    end 
    if(N7924) begin
      { mem[1547:1547] } <= { data_i[27:27] };
    end 
    if(N7923) begin
      { mem[1546:1546] } <= { data_i[26:26] };
    end 
    if(N7922) begin
      { mem[1545:1545] } <= { data_i[25:25] };
    end 
    if(N7921) begin
      { mem[1544:1544] } <= { data_i[24:24] };
    end 
    if(N7920) begin
      { mem[1543:1543] } <= { data_i[23:23] };
    end 
    if(N7919) begin
      { mem[1542:1542] } <= { data_i[22:22] };
    end 
    if(N7918) begin
      { mem[1541:1541] } <= { data_i[21:21] };
    end 
    if(N7917) begin
      { mem[1540:1540] } <= { data_i[20:20] };
    end 
    if(N7916) begin
      { mem[1539:1539] } <= { data_i[19:19] };
    end 
    if(N7915) begin
      { mem[1538:1538] } <= { data_i[18:18] };
    end 
    if(N7914) begin
      { mem[1537:1537] } <= { data_i[17:17] };
    end 
    if(N7913) begin
      { mem[1536:1536] } <= { data_i[16:16] };
    end 
    if(N7912) begin
      { mem[1535:1535] } <= { data_i[15:15] };
    end 
    if(N7911) begin
      { mem[1534:1534] } <= { data_i[14:14] };
    end 
    if(N7910) begin
      { mem[1533:1533] } <= { data_i[13:13] };
    end 
    if(N7909) begin
      { mem[1532:1532] } <= { data_i[12:12] };
    end 
    if(N7908) begin
      { mem[1531:1531] } <= { data_i[11:11] };
    end 
    if(N7907) begin
      { mem[1530:1530] } <= { data_i[10:10] };
    end 
    if(N7906) begin
      { mem[1529:1529] } <= { data_i[9:9] };
    end 
    if(N7905) begin
      { mem[1528:1528] } <= { data_i[8:8] };
    end 
    if(N7904) begin
      { mem[1527:1527] } <= { data_i[7:7] };
    end 
    if(N7903) begin
      { mem[1526:1526] } <= { data_i[6:6] };
    end 
    if(N7902) begin
      { mem[1525:1525] } <= { data_i[5:5] };
    end 
    if(N7901) begin
      { mem[1524:1524] } <= { data_i[4:4] };
    end 
    if(N7900) begin
      { mem[1523:1523] } <= { data_i[3:3] };
    end 
    if(N7899) begin
      { mem[1522:1522] } <= { data_i[2:2] };
    end 
    if(N7898) begin
      { mem[1521:1521] } <= { data_i[1:1] };
    end 
    if(N7897) begin
      { mem[1520:1520] } <= { data_i[0:0] };
    end 
    if(N7896) begin
      { mem[1519:1519] } <= { data_i[79:79] };
    end 
    if(N7895) begin
      { mem[1518:1518] } <= { data_i[78:78] };
    end 
    if(N7894) begin
      { mem[1517:1517] } <= { data_i[77:77] };
    end 
    if(N7893) begin
      { mem[1516:1516] } <= { data_i[76:76] };
    end 
    if(N7892) begin
      { mem[1515:1515] } <= { data_i[75:75] };
    end 
    if(N7891) begin
      { mem[1514:1514] } <= { data_i[74:74] };
    end 
    if(N7890) begin
      { mem[1513:1513] } <= { data_i[73:73] };
    end 
    if(N7889) begin
      { mem[1512:1512] } <= { data_i[72:72] };
    end 
    if(N7888) begin
      { mem[1511:1511] } <= { data_i[71:71] };
    end 
    if(N7887) begin
      { mem[1510:1510] } <= { data_i[70:70] };
    end 
    if(N7886) begin
      { mem[1509:1509] } <= { data_i[69:69] };
    end 
    if(N7885) begin
      { mem[1508:1508] } <= { data_i[68:68] };
    end 
    if(N7884) begin
      { mem[1507:1507] } <= { data_i[67:67] };
    end 
    if(N7883) begin
      { mem[1506:1506] } <= { data_i[66:66] };
    end 
    if(N7882) begin
      { mem[1505:1505] } <= { data_i[65:65] };
    end 
    if(N7881) begin
      { mem[1504:1504] } <= { data_i[64:64] };
    end 
    if(N7880) begin
      { mem[1503:1503] } <= { data_i[63:63] };
    end 
    if(N7879) begin
      { mem[1502:1502] } <= { data_i[62:62] };
    end 
    if(N7878) begin
      { mem[1501:1501] } <= { data_i[61:61] };
    end 
    if(N7877) begin
      { mem[1500:1500] } <= { data_i[60:60] };
    end 
    if(N7876) begin
      { mem[1499:1499] } <= { data_i[59:59] };
    end 
    if(N7875) begin
      { mem[1498:1498] } <= { data_i[58:58] };
    end 
    if(N7874) begin
      { mem[1497:1497] } <= { data_i[57:57] };
    end 
    if(N7873) begin
      { mem[1496:1496] } <= { data_i[56:56] };
    end 
    if(N7872) begin
      { mem[1495:1495] } <= { data_i[55:55] };
    end 
    if(N7871) begin
      { mem[1494:1494] } <= { data_i[54:54] };
    end 
    if(N7870) begin
      { mem[1493:1493] } <= { data_i[53:53] };
    end 
    if(N7869) begin
      { mem[1492:1492] } <= { data_i[52:52] };
    end 
    if(N7868) begin
      { mem[1491:1491] } <= { data_i[51:51] };
    end 
    if(N7867) begin
      { mem[1490:1490] } <= { data_i[50:50] };
    end 
    if(N7866) begin
      { mem[1489:1489] } <= { data_i[49:49] };
    end 
    if(N7865) begin
      { mem[1488:1488] } <= { data_i[48:48] };
    end 
    if(N7864) begin
      { mem[1487:1487] } <= { data_i[47:47] };
    end 
    if(N7863) begin
      { mem[1486:1486] } <= { data_i[46:46] };
    end 
    if(N7862) begin
      { mem[1485:1485] } <= { data_i[45:45] };
    end 
    if(N7861) begin
      { mem[1484:1484] } <= { data_i[44:44] };
    end 
    if(N7860) begin
      { mem[1483:1483] } <= { data_i[43:43] };
    end 
    if(N7859) begin
      { mem[1482:1482] } <= { data_i[42:42] };
    end 
    if(N7858) begin
      { mem[1481:1481] } <= { data_i[41:41] };
    end 
    if(N7857) begin
      { mem[1480:1480] } <= { data_i[40:40] };
    end 
    if(N7856) begin
      { mem[1479:1479] } <= { data_i[39:39] };
    end 
    if(N7855) begin
      { mem[1478:1478] } <= { data_i[38:38] };
    end 
    if(N7854) begin
      { mem[1477:1477] } <= { data_i[37:37] };
    end 
    if(N7853) begin
      { mem[1476:1476] } <= { data_i[36:36] };
    end 
    if(N7852) begin
      { mem[1475:1475] } <= { data_i[35:35] };
    end 
    if(N7851) begin
      { mem[1474:1474] } <= { data_i[34:34] };
    end 
    if(N7850) begin
      { mem[1473:1473] } <= { data_i[33:33] };
    end 
    if(N7849) begin
      { mem[1472:1472] } <= { data_i[32:32] };
    end 
    if(N7848) begin
      { mem[1471:1471] } <= { data_i[31:31] };
    end 
    if(N7847) begin
      { mem[1470:1470] } <= { data_i[30:30] };
    end 
    if(N7846) begin
      { mem[1469:1469] } <= { data_i[29:29] };
    end 
    if(N7845) begin
      { mem[1468:1468] } <= { data_i[28:28] };
    end 
    if(N7844) begin
      { mem[1467:1467] } <= { data_i[27:27] };
    end 
    if(N7843) begin
      { mem[1466:1466] } <= { data_i[26:26] };
    end 
    if(N7842) begin
      { mem[1465:1465] } <= { data_i[25:25] };
    end 
    if(N7841) begin
      { mem[1464:1464] } <= { data_i[24:24] };
    end 
    if(N7840) begin
      { mem[1463:1463] } <= { data_i[23:23] };
    end 
    if(N7839) begin
      { mem[1462:1462] } <= { data_i[22:22] };
    end 
    if(N7838) begin
      { mem[1461:1461] } <= { data_i[21:21] };
    end 
    if(N7837) begin
      { mem[1460:1460] } <= { data_i[20:20] };
    end 
    if(N7836) begin
      { mem[1459:1459] } <= { data_i[19:19] };
    end 
    if(N7835) begin
      { mem[1458:1458] } <= { data_i[18:18] };
    end 
    if(N7834) begin
      { mem[1457:1457] } <= { data_i[17:17] };
    end 
    if(N7833) begin
      { mem[1456:1456] } <= { data_i[16:16] };
    end 
    if(N7832) begin
      { mem[1455:1455] } <= { data_i[15:15] };
    end 
    if(N7831) begin
      { mem[1454:1454] } <= { data_i[14:14] };
    end 
    if(N7830) begin
      { mem[1453:1453] } <= { data_i[13:13] };
    end 
    if(N7829) begin
      { mem[1452:1452] } <= { data_i[12:12] };
    end 
    if(N7828) begin
      { mem[1451:1451] } <= { data_i[11:11] };
    end 
    if(N7827) begin
      { mem[1450:1450] } <= { data_i[10:10] };
    end 
    if(N7826) begin
      { mem[1449:1449] } <= { data_i[9:9] };
    end 
    if(N7825) begin
      { mem[1448:1448] } <= { data_i[8:8] };
    end 
    if(N7824) begin
      { mem[1447:1447] } <= { data_i[7:7] };
    end 
    if(N7823) begin
      { mem[1446:1446] } <= { data_i[6:6] };
    end 
    if(N7822) begin
      { mem[1445:1445] } <= { data_i[5:5] };
    end 
    if(N7821) begin
      { mem[1444:1444] } <= { data_i[4:4] };
    end 
    if(N7820) begin
      { mem[1443:1443] } <= { data_i[3:3] };
    end 
    if(N7819) begin
      { mem[1442:1442] } <= { data_i[2:2] };
    end 
    if(N7818) begin
      { mem[1441:1441] } <= { data_i[1:1] };
    end 
    if(N7817) begin
      { mem[1440:1440] } <= { data_i[0:0] };
    end 
    if(N7816) begin
      { mem[1439:1439] } <= { data_i[79:79] };
    end 
    if(N7815) begin
      { mem[1438:1438] } <= { data_i[78:78] };
    end 
    if(N7814) begin
      { mem[1437:1437] } <= { data_i[77:77] };
    end 
    if(N7813) begin
      { mem[1436:1436] } <= { data_i[76:76] };
    end 
    if(N7812) begin
      { mem[1435:1435] } <= { data_i[75:75] };
    end 
    if(N7811) begin
      { mem[1434:1434] } <= { data_i[74:74] };
    end 
    if(N7810) begin
      { mem[1433:1433] } <= { data_i[73:73] };
    end 
    if(N7809) begin
      { mem[1432:1432] } <= { data_i[72:72] };
    end 
    if(N7808) begin
      { mem[1431:1431] } <= { data_i[71:71] };
    end 
    if(N7807) begin
      { mem[1430:1430] } <= { data_i[70:70] };
    end 
    if(N7806) begin
      { mem[1429:1429] } <= { data_i[69:69] };
    end 
    if(N7805) begin
      { mem[1428:1428] } <= { data_i[68:68] };
    end 
    if(N7804) begin
      { mem[1427:1427] } <= { data_i[67:67] };
    end 
    if(N7803) begin
      { mem[1426:1426] } <= { data_i[66:66] };
    end 
    if(N7802) begin
      { mem[1425:1425] } <= { data_i[65:65] };
    end 
    if(N7801) begin
      { mem[1424:1424] } <= { data_i[64:64] };
    end 
    if(N7800) begin
      { mem[1423:1423] } <= { data_i[63:63] };
    end 
    if(N7799) begin
      { mem[1422:1422] } <= { data_i[62:62] };
    end 
    if(N7798) begin
      { mem[1421:1421] } <= { data_i[61:61] };
    end 
    if(N7797) begin
      { mem[1420:1420] } <= { data_i[60:60] };
    end 
    if(N7796) begin
      { mem[1419:1419] } <= { data_i[59:59] };
    end 
    if(N7795) begin
      { mem[1418:1418] } <= { data_i[58:58] };
    end 
    if(N7794) begin
      { mem[1417:1417] } <= { data_i[57:57] };
    end 
    if(N7793) begin
      { mem[1416:1416] } <= { data_i[56:56] };
    end 
    if(N7792) begin
      { mem[1415:1415] } <= { data_i[55:55] };
    end 
    if(N7791) begin
      { mem[1414:1414] } <= { data_i[54:54] };
    end 
    if(N7790) begin
      { mem[1413:1413] } <= { data_i[53:53] };
    end 
    if(N7789) begin
      { mem[1412:1412] } <= { data_i[52:52] };
    end 
    if(N7788) begin
      { mem[1411:1411] } <= { data_i[51:51] };
    end 
    if(N7787) begin
      { mem[1410:1410] } <= { data_i[50:50] };
    end 
    if(N7786) begin
      { mem[1409:1409] } <= { data_i[49:49] };
    end 
    if(N7785) begin
      { mem[1408:1408] } <= { data_i[48:48] };
    end 
    if(N7784) begin
      { mem[1407:1407] } <= { data_i[47:47] };
    end 
    if(N7783) begin
      { mem[1406:1406] } <= { data_i[46:46] };
    end 
    if(N7782) begin
      { mem[1405:1405] } <= { data_i[45:45] };
    end 
    if(N7781) begin
      { mem[1404:1404] } <= { data_i[44:44] };
    end 
    if(N7780) begin
      { mem[1403:1403] } <= { data_i[43:43] };
    end 
    if(N7779) begin
      { mem[1402:1402] } <= { data_i[42:42] };
    end 
    if(N7778) begin
      { mem[1401:1401] } <= { data_i[41:41] };
    end 
    if(N7777) begin
      { mem[1400:1400] } <= { data_i[40:40] };
    end 
    if(N7776) begin
      { mem[1399:1399] } <= { data_i[39:39] };
    end 
    if(N7775) begin
      { mem[1398:1398] } <= { data_i[38:38] };
    end 
    if(N7774) begin
      { mem[1397:1397] } <= { data_i[37:37] };
    end 
    if(N7773) begin
      { mem[1396:1396] } <= { data_i[36:36] };
    end 
    if(N7772) begin
      { mem[1395:1395] } <= { data_i[35:35] };
    end 
    if(N7771) begin
      { mem[1394:1394] } <= { data_i[34:34] };
    end 
    if(N7770) begin
      { mem[1393:1393] } <= { data_i[33:33] };
    end 
    if(N7769) begin
      { mem[1392:1392] } <= { data_i[32:32] };
    end 
    if(N7768) begin
      { mem[1391:1391] } <= { data_i[31:31] };
    end 
    if(N7767) begin
      { mem[1390:1390] } <= { data_i[30:30] };
    end 
    if(N7766) begin
      { mem[1389:1389] } <= { data_i[29:29] };
    end 
    if(N7765) begin
      { mem[1388:1388] } <= { data_i[28:28] };
    end 
    if(N7764) begin
      { mem[1387:1387] } <= { data_i[27:27] };
    end 
    if(N7763) begin
      { mem[1386:1386] } <= { data_i[26:26] };
    end 
    if(N7762) begin
      { mem[1385:1385] } <= { data_i[25:25] };
    end 
    if(N7761) begin
      { mem[1384:1384] } <= { data_i[24:24] };
    end 
    if(N7760) begin
      { mem[1383:1383] } <= { data_i[23:23] };
    end 
    if(N7759) begin
      { mem[1382:1382] } <= { data_i[22:22] };
    end 
    if(N7758) begin
      { mem[1381:1381] } <= { data_i[21:21] };
    end 
    if(N7757) begin
      { mem[1380:1380] } <= { data_i[20:20] };
    end 
    if(N7756) begin
      { mem[1379:1379] } <= { data_i[19:19] };
    end 
    if(N7755) begin
      { mem[1378:1378] } <= { data_i[18:18] };
    end 
    if(N7754) begin
      { mem[1377:1377] } <= { data_i[17:17] };
    end 
    if(N7753) begin
      { mem[1376:1376] } <= { data_i[16:16] };
    end 
    if(N7752) begin
      { mem[1375:1375] } <= { data_i[15:15] };
    end 
    if(N7751) begin
      { mem[1374:1374] } <= { data_i[14:14] };
    end 
    if(N7750) begin
      { mem[1373:1373] } <= { data_i[13:13] };
    end 
    if(N7749) begin
      { mem[1372:1372] } <= { data_i[12:12] };
    end 
    if(N7748) begin
      { mem[1371:1371] } <= { data_i[11:11] };
    end 
    if(N7747) begin
      { mem[1370:1370] } <= { data_i[10:10] };
    end 
    if(N7746) begin
      { mem[1369:1369] } <= { data_i[9:9] };
    end 
    if(N7745) begin
      { mem[1368:1368] } <= { data_i[8:8] };
    end 
    if(N7744) begin
      { mem[1367:1367] } <= { data_i[7:7] };
    end 
    if(N7743) begin
      { mem[1366:1366] } <= { data_i[6:6] };
    end 
    if(N7742) begin
      { mem[1365:1365] } <= { data_i[5:5] };
    end 
    if(N7741) begin
      { mem[1364:1364] } <= { data_i[4:4] };
    end 
    if(N7740) begin
      { mem[1363:1363] } <= { data_i[3:3] };
    end 
    if(N7739) begin
      { mem[1362:1362] } <= { data_i[2:2] };
    end 
    if(N7738) begin
      { mem[1361:1361] } <= { data_i[1:1] };
    end 
    if(N7737) begin
      { mem[1360:1360] } <= { data_i[0:0] };
    end 
    if(N7736) begin
      { mem[1359:1359] } <= { data_i[79:79] };
    end 
    if(N7735) begin
      { mem[1358:1358] } <= { data_i[78:78] };
    end 
    if(N7734) begin
      { mem[1357:1357] } <= { data_i[77:77] };
    end 
    if(N7733) begin
      { mem[1356:1356] } <= { data_i[76:76] };
    end 
    if(N7732) begin
      { mem[1355:1355] } <= { data_i[75:75] };
    end 
    if(N7731) begin
      { mem[1354:1354] } <= { data_i[74:74] };
    end 
    if(N7730) begin
      { mem[1353:1353] } <= { data_i[73:73] };
    end 
    if(N7729) begin
      { mem[1352:1352] } <= { data_i[72:72] };
    end 
    if(N7728) begin
      { mem[1351:1351] } <= { data_i[71:71] };
    end 
    if(N7727) begin
      { mem[1350:1350] } <= { data_i[70:70] };
    end 
    if(N7726) begin
      { mem[1349:1349] } <= { data_i[69:69] };
    end 
    if(N7725) begin
      { mem[1348:1348] } <= { data_i[68:68] };
    end 
    if(N7724) begin
      { mem[1347:1347] } <= { data_i[67:67] };
    end 
    if(N7723) begin
      { mem[1346:1346] } <= { data_i[66:66] };
    end 
    if(N7722) begin
      { mem[1345:1345] } <= { data_i[65:65] };
    end 
    if(N7721) begin
      { mem[1344:1344] } <= { data_i[64:64] };
    end 
    if(N7720) begin
      { mem[1343:1343] } <= { data_i[63:63] };
    end 
    if(N7719) begin
      { mem[1342:1342] } <= { data_i[62:62] };
    end 
    if(N7718) begin
      { mem[1341:1341] } <= { data_i[61:61] };
    end 
    if(N7717) begin
      { mem[1340:1340] } <= { data_i[60:60] };
    end 
    if(N7716) begin
      { mem[1339:1339] } <= { data_i[59:59] };
    end 
    if(N7715) begin
      { mem[1338:1338] } <= { data_i[58:58] };
    end 
    if(N7714) begin
      { mem[1337:1337] } <= { data_i[57:57] };
    end 
    if(N7713) begin
      { mem[1336:1336] } <= { data_i[56:56] };
    end 
    if(N7712) begin
      { mem[1335:1335] } <= { data_i[55:55] };
    end 
    if(N7711) begin
      { mem[1334:1334] } <= { data_i[54:54] };
    end 
    if(N7710) begin
      { mem[1333:1333] } <= { data_i[53:53] };
    end 
    if(N7709) begin
      { mem[1332:1332] } <= { data_i[52:52] };
    end 
    if(N7708) begin
      { mem[1331:1331] } <= { data_i[51:51] };
    end 
    if(N7707) begin
      { mem[1330:1330] } <= { data_i[50:50] };
    end 
    if(N7706) begin
      { mem[1329:1329] } <= { data_i[49:49] };
    end 
    if(N7705) begin
      { mem[1328:1328] } <= { data_i[48:48] };
    end 
    if(N7704) begin
      { mem[1327:1327] } <= { data_i[47:47] };
    end 
    if(N7703) begin
      { mem[1326:1326] } <= { data_i[46:46] };
    end 
    if(N7702) begin
      { mem[1325:1325] } <= { data_i[45:45] };
    end 
    if(N7701) begin
      { mem[1324:1324] } <= { data_i[44:44] };
    end 
    if(N7700) begin
      { mem[1323:1323] } <= { data_i[43:43] };
    end 
    if(N7699) begin
      { mem[1322:1322] } <= { data_i[42:42] };
    end 
    if(N7698) begin
      { mem[1321:1321] } <= { data_i[41:41] };
    end 
    if(N7697) begin
      { mem[1320:1320] } <= { data_i[40:40] };
    end 
    if(N7696) begin
      { mem[1319:1319] } <= { data_i[39:39] };
    end 
    if(N7695) begin
      { mem[1318:1318] } <= { data_i[38:38] };
    end 
    if(N7694) begin
      { mem[1317:1317] } <= { data_i[37:37] };
    end 
    if(N7693) begin
      { mem[1316:1316] } <= { data_i[36:36] };
    end 
    if(N7692) begin
      { mem[1315:1315] } <= { data_i[35:35] };
    end 
    if(N7691) begin
      { mem[1314:1314] } <= { data_i[34:34] };
    end 
    if(N7690) begin
      { mem[1313:1313] } <= { data_i[33:33] };
    end 
    if(N7689) begin
      { mem[1312:1312] } <= { data_i[32:32] };
    end 
    if(N7688) begin
      { mem[1311:1311] } <= { data_i[31:31] };
    end 
    if(N7687) begin
      { mem[1310:1310] } <= { data_i[30:30] };
    end 
    if(N7686) begin
      { mem[1309:1309] } <= { data_i[29:29] };
    end 
    if(N7685) begin
      { mem[1308:1308] } <= { data_i[28:28] };
    end 
    if(N7684) begin
      { mem[1307:1307] } <= { data_i[27:27] };
    end 
    if(N7683) begin
      { mem[1306:1306] } <= { data_i[26:26] };
    end 
    if(N7682) begin
      { mem[1305:1305] } <= { data_i[25:25] };
    end 
    if(N7681) begin
      { mem[1304:1304] } <= { data_i[24:24] };
    end 
    if(N7680) begin
      { mem[1303:1303] } <= { data_i[23:23] };
    end 
    if(N7679) begin
      { mem[1302:1302] } <= { data_i[22:22] };
    end 
    if(N7678) begin
      { mem[1301:1301] } <= { data_i[21:21] };
    end 
    if(N7677) begin
      { mem[1300:1300] } <= { data_i[20:20] };
    end 
    if(N7676) begin
      { mem[1299:1299] } <= { data_i[19:19] };
    end 
    if(N7675) begin
      { mem[1298:1298] } <= { data_i[18:18] };
    end 
    if(N7674) begin
      { mem[1297:1297] } <= { data_i[17:17] };
    end 
    if(N7673) begin
      { mem[1296:1296] } <= { data_i[16:16] };
    end 
    if(N7672) begin
      { mem[1295:1295] } <= { data_i[15:15] };
    end 
    if(N7671) begin
      { mem[1294:1294] } <= { data_i[14:14] };
    end 
    if(N7670) begin
      { mem[1293:1293] } <= { data_i[13:13] };
    end 
    if(N7669) begin
      { mem[1292:1292] } <= { data_i[12:12] };
    end 
    if(N7668) begin
      { mem[1291:1291] } <= { data_i[11:11] };
    end 
    if(N7667) begin
      { mem[1290:1290] } <= { data_i[10:10] };
    end 
    if(N7666) begin
      { mem[1289:1289] } <= { data_i[9:9] };
    end 
    if(N7665) begin
      { mem[1288:1288] } <= { data_i[8:8] };
    end 
    if(N7664) begin
      { mem[1287:1287] } <= { data_i[7:7] };
    end 
    if(N7663) begin
      { mem[1286:1286] } <= { data_i[6:6] };
    end 
    if(N7662) begin
      { mem[1285:1285] } <= { data_i[5:5] };
    end 
    if(N7661) begin
      { mem[1284:1284] } <= { data_i[4:4] };
    end 
    if(N7660) begin
      { mem[1283:1283] } <= { data_i[3:3] };
    end 
    if(N7659) begin
      { mem[1282:1282] } <= { data_i[2:2] };
    end 
    if(N7658) begin
      { mem[1281:1281] } <= { data_i[1:1] };
    end 
    if(N7657) begin
      { mem[1280:1280] } <= { data_i[0:0] };
    end 
    if(N7656) begin
      { mem[1279:1279] } <= { data_i[79:79] };
    end 
    if(N7655) begin
      { mem[1278:1278] } <= { data_i[78:78] };
    end 
    if(N7654) begin
      { mem[1277:1277] } <= { data_i[77:77] };
    end 
    if(N7653) begin
      { mem[1276:1276] } <= { data_i[76:76] };
    end 
    if(N7652) begin
      { mem[1275:1275] } <= { data_i[75:75] };
    end 
    if(N7651) begin
      { mem[1274:1274] } <= { data_i[74:74] };
    end 
    if(N7650) begin
      { mem[1273:1273] } <= { data_i[73:73] };
    end 
    if(N7649) begin
      { mem[1272:1272] } <= { data_i[72:72] };
    end 
    if(N7648) begin
      { mem[1271:1271] } <= { data_i[71:71] };
    end 
    if(N7647) begin
      { mem[1270:1270] } <= { data_i[70:70] };
    end 
    if(N7646) begin
      { mem[1269:1269] } <= { data_i[69:69] };
    end 
    if(N7645) begin
      { mem[1268:1268] } <= { data_i[68:68] };
    end 
    if(N7644) begin
      { mem[1267:1267] } <= { data_i[67:67] };
    end 
    if(N7643) begin
      { mem[1266:1266] } <= { data_i[66:66] };
    end 
    if(N7642) begin
      { mem[1265:1265] } <= { data_i[65:65] };
    end 
    if(N7641) begin
      { mem[1264:1264] } <= { data_i[64:64] };
    end 
    if(N7640) begin
      { mem[1263:1263] } <= { data_i[63:63] };
    end 
    if(N7639) begin
      { mem[1262:1262] } <= { data_i[62:62] };
    end 
    if(N7638) begin
      { mem[1261:1261] } <= { data_i[61:61] };
    end 
    if(N7637) begin
      { mem[1260:1260] } <= { data_i[60:60] };
    end 
    if(N7636) begin
      { mem[1259:1259] } <= { data_i[59:59] };
    end 
    if(N7635) begin
      { mem[1258:1258] } <= { data_i[58:58] };
    end 
    if(N7634) begin
      { mem[1257:1257] } <= { data_i[57:57] };
    end 
    if(N7633) begin
      { mem[1256:1256] } <= { data_i[56:56] };
    end 
    if(N7632) begin
      { mem[1255:1255] } <= { data_i[55:55] };
    end 
    if(N7631) begin
      { mem[1254:1254] } <= { data_i[54:54] };
    end 
    if(N7630) begin
      { mem[1253:1253] } <= { data_i[53:53] };
    end 
    if(N7629) begin
      { mem[1252:1252] } <= { data_i[52:52] };
    end 
    if(N7628) begin
      { mem[1251:1251] } <= { data_i[51:51] };
    end 
    if(N7627) begin
      { mem[1250:1250] } <= { data_i[50:50] };
    end 
    if(N7626) begin
      { mem[1249:1249] } <= { data_i[49:49] };
    end 
    if(N7625) begin
      { mem[1248:1248] } <= { data_i[48:48] };
    end 
    if(N7624) begin
      { mem[1247:1247] } <= { data_i[47:47] };
    end 
    if(N7623) begin
      { mem[1246:1246] } <= { data_i[46:46] };
    end 
    if(N7622) begin
      { mem[1245:1245] } <= { data_i[45:45] };
    end 
    if(N7621) begin
      { mem[1244:1244] } <= { data_i[44:44] };
    end 
    if(N7620) begin
      { mem[1243:1243] } <= { data_i[43:43] };
    end 
    if(N7619) begin
      { mem[1242:1242] } <= { data_i[42:42] };
    end 
    if(N7618) begin
      { mem[1241:1241] } <= { data_i[41:41] };
    end 
    if(N7617) begin
      { mem[1240:1240] } <= { data_i[40:40] };
    end 
    if(N7616) begin
      { mem[1239:1239] } <= { data_i[39:39] };
    end 
    if(N7615) begin
      { mem[1238:1238] } <= { data_i[38:38] };
    end 
    if(N7614) begin
      { mem[1237:1237] } <= { data_i[37:37] };
    end 
    if(N7613) begin
      { mem[1236:1236] } <= { data_i[36:36] };
    end 
    if(N7612) begin
      { mem[1235:1235] } <= { data_i[35:35] };
    end 
    if(N7611) begin
      { mem[1234:1234] } <= { data_i[34:34] };
    end 
    if(N7610) begin
      { mem[1233:1233] } <= { data_i[33:33] };
    end 
    if(N7609) begin
      { mem[1232:1232] } <= { data_i[32:32] };
    end 
    if(N7608) begin
      { mem[1231:1231] } <= { data_i[31:31] };
    end 
    if(N7607) begin
      { mem[1230:1230] } <= { data_i[30:30] };
    end 
    if(N7606) begin
      { mem[1229:1229] } <= { data_i[29:29] };
    end 
    if(N7605) begin
      { mem[1228:1228] } <= { data_i[28:28] };
    end 
    if(N7604) begin
      { mem[1227:1227] } <= { data_i[27:27] };
    end 
    if(N7603) begin
      { mem[1226:1226] } <= { data_i[26:26] };
    end 
    if(N7602) begin
      { mem[1225:1225] } <= { data_i[25:25] };
    end 
    if(N7601) begin
      { mem[1224:1224] } <= { data_i[24:24] };
    end 
    if(N7600) begin
      { mem[1223:1223] } <= { data_i[23:23] };
    end 
    if(N7599) begin
      { mem[1222:1222] } <= { data_i[22:22] };
    end 
    if(N7598) begin
      { mem[1221:1221] } <= { data_i[21:21] };
    end 
    if(N7597) begin
      { mem[1220:1220] } <= { data_i[20:20] };
    end 
    if(N7596) begin
      { mem[1219:1219] } <= { data_i[19:19] };
    end 
    if(N7595) begin
      { mem[1218:1218] } <= { data_i[18:18] };
    end 
    if(N7594) begin
      { mem[1217:1217] } <= { data_i[17:17] };
    end 
    if(N7593) begin
      { mem[1216:1216] } <= { data_i[16:16] };
    end 
    if(N7592) begin
      { mem[1215:1215] } <= { data_i[15:15] };
    end 
    if(N7591) begin
      { mem[1214:1214] } <= { data_i[14:14] };
    end 
    if(N7590) begin
      { mem[1213:1213] } <= { data_i[13:13] };
    end 
    if(N7589) begin
      { mem[1212:1212] } <= { data_i[12:12] };
    end 
    if(N7588) begin
      { mem[1211:1211] } <= { data_i[11:11] };
    end 
    if(N7587) begin
      { mem[1210:1210] } <= { data_i[10:10] };
    end 
    if(N7586) begin
      { mem[1209:1209] } <= { data_i[9:9] };
    end 
    if(N7585) begin
      { mem[1208:1208] } <= { data_i[8:8] };
    end 
    if(N7584) begin
      { mem[1207:1207] } <= { data_i[7:7] };
    end 
    if(N7583) begin
      { mem[1206:1206] } <= { data_i[6:6] };
    end 
    if(N7582) begin
      { mem[1205:1205] } <= { data_i[5:5] };
    end 
    if(N7581) begin
      { mem[1204:1204] } <= { data_i[4:4] };
    end 
    if(N7580) begin
      { mem[1203:1203] } <= { data_i[3:3] };
    end 
    if(N7579) begin
      { mem[1202:1202] } <= { data_i[2:2] };
    end 
    if(N7578) begin
      { mem[1201:1201] } <= { data_i[1:1] };
    end 
    if(N7577) begin
      { mem[1200:1200] } <= { data_i[0:0] };
    end 
    if(N7576) begin
      { mem[1199:1199] } <= { data_i[79:79] };
    end 
    if(N7575) begin
      { mem[1198:1198] } <= { data_i[78:78] };
    end 
    if(N7574) begin
      { mem[1197:1197] } <= { data_i[77:77] };
    end 
    if(N7573) begin
      { mem[1196:1196] } <= { data_i[76:76] };
    end 
    if(N7572) begin
      { mem[1195:1195] } <= { data_i[75:75] };
    end 
    if(N7571) begin
      { mem[1194:1194] } <= { data_i[74:74] };
    end 
    if(N7570) begin
      { mem[1193:1193] } <= { data_i[73:73] };
    end 
    if(N7569) begin
      { mem[1192:1192] } <= { data_i[72:72] };
    end 
    if(N7568) begin
      { mem[1191:1191] } <= { data_i[71:71] };
    end 
    if(N7567) begin
      { mem[1190:1190] } <= { data_i[70:70] };
    end 
    if(N7566) begin
      { mem[1189:1189] } <= { data_i[69:69] };
    end 
    if(N7565) begin
      { mem[1188:1188] } <= { data_i[68:68] };
    end 
    if(N7564) begin
      { mem[1187:1187] } <= { data_i[67:67] };
    end 
    if(N7563) begin
      { mem[1186:1186] } <= { data_i[66:66] };
    end 
    if(N7562) begin
      { mem[1185:1185] } <= { data_i[65:65] };
    end 
    if(N7561) begin
      { mem[1184:1184] } <= { data_i[64:64] };
    end 
    if(N7560) begin
      { mem[1183:1183] } <= { data_i[63:63] };
    end 
    if(N7559) begin
      { mem[1182:1182] } <= { data_i[62:62] };
    end 
    if(N7558) begin
      { mem[1181:1181] } <= { data_i[61:61] };
    end 
    if(N7557) begin
      { mem[1180:1180] } <= { data_i[60:60] };
    end 
    if(N7556) begin
      { mem[1179:1179] } <= { data_i[59:59] };
    end 
    if(N7555) begin
      { mem[1178:1178] } <= { data_i[58:58] };
    end 
    if(N7554) begin
      { mem[1177:1177] } <= { data_i[57:57] };
    end 
    if(N7553) begin
      { mem[1176:1176] } <= { data_i[56:56] };
    end 
    if(N7552) begin
      { mem[1175:1175] } <= { data_i[55:55] };
    end 
    if(N7551) begin
      { mem[1174:1174] } <= { data_i[54:54] };
    end 
    if(N7550) begin
      { mem[1173:1173] } <= { data_i[53:53] };
    end 
    if(N7549) begin
      { mem[1172:1172] } <= { data_i[52:52] };
    end 
    if(N7548) begin
      { mem[1171:1171] } <= { data_i[51:51] };
    end 
    if(N7547) begin
      { mem[1170:1170] } <= { data_i[50:50] };
    end 
    if(N7546) begin
      { mem[1169:1169] } <= { data_i[49:49] };
    end 
    if(N7545) begin
      { mem[1168:1168] } <= { data_i[48:48] };
    end 
    if(N7544) begin
      { mem[1167:1167] } <= { data_i[47:47] };
    end 
    if(N7543) begin
      { mem[1166:1166] } <= { data_i[46:46] };
    end 
    if(N7542) begin
      { mem[1165:1165] } <= { data_i[45:45] };
    end 
    if(N7541) begin
      { mem[1164:1164] } <= { data_i[44:44] };
    end 
    if(N7540) begin
      { mem[1163:1163] } <= { data_i[43:43] };
    end 
    if(N7539) begin
      { mem[1162:1162] } <= { data_i[42:42] };
    end 
    if(N7538) begin
      { mem[1161:1161] } <= { data_i[41:41] };
    end 
    if(N7537) begin
      { mem[1160:1160] } <= { data_i[40:40] };
    end 
    if(N7536) begin
      { mem[1159:1159] } <= { data_i[39:39] };
    end 
    if(N7535) begin
      { mem[1158:1158] } <= { data_i[38:38] };
    end 
    if(N7534) begin
      { mem[1157:1157] } <= { data_i[37:37] };
    end 
    if(N7533) begin
      { mem[1156:1156] } <= { data_i[36:36] };
    end 
    if(N7532) begin
      { mem[1155:1155] } <= { data_i[35:35] };
    end 
    if(N7531) begin
      { mem[1154:1154] } <= { data_i[34:34] };
    end 
    if(N7530) begin
      { mem[1153:1153] } <= { data_i[33:33] };
    end 
    if(N7529) begin
      { mem[1152:1152] } <= { data_i[32:32] };
    end 
    if(N7528) begin
      { mem[1151:1151] } <= { data_i[31:31] };
    end 
    if(N7527) begin
      { mem[1150:1150] } <= { data_i[30:30] };
    end 
    if(N7526) begin
      { mem[1149:1149] } <= { data_i[29:29] };
    end 
    if(N7525) begin
      { mem[1148:1148] } <= { data_i[28:28] };
    end 
    if(N7524) begin
      { mem[1147:1147] } <= { data_i[27:27] };
    end 
    if(N7523) begin
      { mem[1146:1146] } <= { data_i[26:26] };
    end 
    if(N7522) begin
      { mem[1145:1145] } <= { data_i[25:25] };
    end 
    if(N7521) begin
      { mem[1144:1144] } <= { data_i[24:24] };
    end 
    if(N7520) begin
      { mem[1143:1143] } <= { data_i[23:23] };
    end 
    if(N7519) begin
      { mem[1142:1142] } <= { data_i[22:22] };
    end 
    if(N7518) begin
      { mem[1141:1141] } <= { data_i[21:21] };
    end 
    if(N7517) begin
      { mem[1140:1140] } <= { data_i[20:20] };
    end 
    if(N7516) begin
      { mem[1139:1139] } <= { data_i[19:19] };
    end 
    if(N7515) begin
      { mem[1138:1138] } <= { data_i[18:18] };
    end 
    if(N7514) begin
      { mem[1137:1137] } <= { data_i[17:17] };
    end 
    if(N7513) begin
      { mem[1136:1136] } <= { data_i[16:16] };
    end 
    if(N7512) begin
      { mem[1135:1135] } <= { data_i[15:15] };
    end 
    if(N7511) begin
      { mem[1134:1134] } <= { data_i[14:14] };
    end 
    if(N7510) begin
      { mem[1133:1133] } <= { data_i[13:13] };
    end 
    if(N7509) begin
      { mem[1132:1132] } <= { data_i[12:12] };
    end 
    if(N7508) begin
      { mem[1131:1131] } <= { data_i[11:11] };
    end 
    if(N7507) begin
      { mem[1130:1130] } <= { data_i[10:10] };
    end 
    if(N7506) begin
      { mem[1129:1129] } <= { data_i[9:9] };
    end 
    if(N7505) begin
      { mem[1128:1128] } <= { data_i[8:8] };
    end 
    if(N7504) begin
      { mem[1127:1127] } <= { data_i[7:7] };
    end 
    if(N7503) begin
      { mem[1126:1126] } <= { data_i[6:6] };
    end 
    if(N7502) begin
      { mem[1125:1125] } <= { data_i[5:5] };
    end 
    if(N7501) begin
      { mem[1124:1124] } <= { data_i[4:4] };
    end 
    if(N7500) begin
      { mem[1123:1123] } <= { data_i[3:3] };
    end 
    if(N7499) begin
      { mem[1122:1122] } <= { data_i[2:2] };
    end 
    if(N7498) begin
      { mem[1121:1121] } <= { data_i[1:1] };
    end 
    if(N7497) begin
      { mem[1120:1120] } <= { data_i[0:0] };
    end 
    if(N7496) begin
      { mem[1119:1119] } <= { data_i[79:79] };
    end 
    if(N7495) begin
      { mem[1118:1118] } <= { data_i[78:78] };
    end 
    if(N7494) begin
      { mem[1117:1117] } <= { data_i[77:77] };
    end 
    if(N7493) begin
      { mem[1116:1116] } <= { data_i[76:76] };
    end 
    if(N7492) begin
      { mem[1115:1115] } <= { data_i[75:75] };
    end 
    if(N7491) begin
      { mem[1114:1114] } <= { data_i[74:74] };
    end 
    if(N7490) begin
      { mem[1113:1113] } <= { data_i[73:73] };
    end 
    if(N7489) begin
      { mem[1112:1112] } <= { data_i[72:72] };
    end 
    if(N7488) begin
      { mem[1111:1111] } <= { data_i[71:71] };
    end 
    if(N7487) begin
      { mem[1110:1110] } <= { data_i[70:70] };
    end 
    if(N7486) begin
      { mem[1109:1109] } <= { data_i[69:69] };
    end 
    if(N7485) begin
      { mem[1108:1108] } <= { data_i[68:68] };
    end 
    if(N7484) begin
      { mem[1107:1107] } <= { data_i[67:67] };
    end 
    if(N7483) begin
      { mem[1106:1106] } <= { data_i[66:66] };
    end 
    if(N7482) begin
      { mem[1105:1105] } <= { data_i[65:65] };
    end 
    if(N7481) begin
      { mem[1104:1104] } <= { data_i[64:64] };
    end 
    if(N7480) begin
      { mem[1103:1103] } <= { data_i[63:63] };
    end 
    if(N7479) begin
      { mem[1102:1102] } <= { data_i[62:62] };
    end 
    if(N7478) begin
      { mem[1101:1101] } <= { data_i[61:61] };
    end 
    if(N7477) begin
      { mem[1100:1100] } <= { data_i[60:60] };
    end 
    if(N7476) begin
      { mem[1099:1099] } <= { data_i[59:59] };
    end 
    if(N7475) begin
      { mem[1098:1098] } <= { data_i[58:58] };
    end 
    if(N7474) begin
      { mem[1097:1097] } <= { data_i[57:57] };
    end 
    if(N7473) begin
      { mem[1096:1096] } <= { data_i[56:56] };
    end 
    if(N7472) begin
      { mem[1095:1095] } <= { data_i[55:55] };
    end 
    if(N7471) begin
      { mem[1094:1094] } <= { data_i[54:54] };
    end 
    if(N7470) begin
      { mem[1093:1093] } <= { data_i[53:53] };
    end 
    if(N7469) begin
      { mem[1092:1092] } <= { data_i[52:52] };
    end 
    if(N7468) begin
      { mem[1091:1091] } <= { data_i[51:51] };
    end 
    if(N7467) begin
      { mem[1090:1090] } <= { data_i[50:50] };
    end 
    if(N7466) begin
      { mem[1089:1089] } <= { data_i[49:49] };
    end 
    if(N7465) begin
      { mem[1088:1088] } <= { data_i[48:48] };
    end 
    if(N7464) begin
      { mem[1087:1087] } <= { data_i[47:47] };
    end 
    if(N7463) begin
      { mem[1086:1086] } <= { data_i[46:46] };
    end 
    if(N7462) begin
      { mem[1085:1085] } <= { data_i[45:45] };
    end 
    if(N7461) begin
      { mem[1084:1084] } <= { data_i[44:44] };
    end 
    if(N7460) begin
      { mem[1083:1083] } <= { data_i[43:43] };
    end 
    if(N7459) begin
      { mem[1082:1082] } <= { data_i[42:42] };
    end 
    if(N7458) begin
      { mem[1081:1081] } <= { data_i[41:41] };
    end 
    if(N7457) begin
      { mem[1080:1080] } <= { data_i[40:40] };
    end 
    if(N7456) begin
      { mem[1079:1079] } <= { data_i[39:39] };
    end 
    if(N7455) begin
      { mem[1078:1078] } <= { data_i[38:38] };
    end 
    if(N7454) begin
      { mem[1077:1077] } <= { data_i[37:37] };
    end 
    if(N7453) begin
      { mem[1076:1076] } <= { data_i[36:36] };
    end 
    if(N7452) begin
      { mem[1075:1075] } <= { data_i[35:35] };
    end 
    if(N7451) begin
      { mem[1074:1074] } <= { data_i[34:34] };
    end 
    if(N7450) begin
      { mem[1073:1073] } <= { data_i[33:33] };
    end 
    if(N7449) begin
      { mem[1072:1072] } <= { data_i[32:32] };
    end 
    if(N7448) begin
      { mem[1071:1071] } <= { data_i[31:31] };
    end 
    if(N7447) begin
      { mem[1070:1070] } <= { data_i[30:30] };
    end 
    if(N7446) begin
      { mem[1069:1069] } <= { data_i[29:29] };
    end 
    if(N7445) begin
      { mem[1068:1068] } <= { data_i[28:28] };
    end 
    if(N7444) begin
      { mem[1067:1067] } <= { data_i[27:27] };
    end 
    if(N7443) begin
      { mem[1066:1066] } <= { data_i[26:26] };
    end 
    if(N7442) begin
      { mem[1065:1065] } <= { data_i[25:25] };
    end 
    if(N7441) begin
      { mem[1064:1064] } <= { data_i[24:24] };
    end 
    if(N7440) begin
      { mem[1063:1063] } <= { data_i[23:23] };
    end 
    if(N7439) begin
      { mem[1062:1062] } <= { data_i[22:22] };
    end 
    if(N7438) begin
      { mem[1061:1061] } <= { data_i[21:21] };
    end 
    if(N7437) begin
      { mem[1060:1060] } <= { data_i[20:20] };
    end 
    if(N7436) begin
      { mem[1059:1059] } <= { data_i[19:19] };
    end 
    if(N7435) begin
      { mem[1058:1058] } <= { data_i[18:18] };
    end 
    if(N7434) begin
      { mem[1057:1057] } <= { data_i[17:17] };
    end 
    if(N7433) begin
      { mem[1056:1056] } <= { data_i[16:16] };
    end 
    if(N7432) begin
      { mem[1055:1055] } <= { data_i[15:15] };
    end 
    if(N7431) begin
      { mem[1054:1054] } <= { data_i[14:14] };
    end 
    if(N7430) begin
      { mem[1053:1053] } <= { data_i[13:13] };
    end 
    if(N7429) begin
      { mem[1052:1052] } <= { data_i[12:12] };
    end 
    if(N7428) begin
      { mem[1051:1051] } <= { data_i[11:11] };
    end 
    if(N7427) begin
      { mem[1050:1050] } <= { data_i[10:10] };
    end 
    if(N7426) begin
      { mem[1049:1049] } <= { data_i[9:9] };
    end 
    if(N7425) begin
      { mem[1048:1048] } <= { data_i[8:8] };
    end 
    if(N7424) begin
      { mem[1047:1047] } <= { data_i[7:7] };
    end 
    if(N7423) begin
      { mem[1046:1046] } <= { data_i[6:6] };
    end 
    if(N7422) begin
      { mem[1045:1045] } <= { data_i[5:5] };
    end 
    if(N7421) begin
      { mem[1044:1044] } <= { data_i[4:4] };
    end 
    if(N7420) begin
      { mem[1043:1043] } <= { data_i[3:3] };
    end 
    if(N7419) begin
      { mem[1042:1042] } <= { data_i[2:2] };
    end 
    if(N7418) begin
      { mem[1041:1041] } <= { data_i[1:1] };
    end 
    if(N7417) begin
      { mem[1040:1040] } <= { data_i[0:0] };
    end 
    if(N7416) begin
      { mem[1039:1039] } <= { data_i[79:79] };
    end 
    if(N7415) begin
      { mem[1038:1038] } <= { data_i[78:78] };
    end 
    if(N7414) begin
      { mem[1037:1037] } <= { data_i[77:77] };
    end 
    if(N7413) begin
      { mem[1036:1036] } <= { data_i[76:76] };
    end 
    if(N7412) begin
      { mem[1035:1035] } <= { data_i[75:75] };
    end 
    if(N7411) begin
      { mem[1034:1034] } <= { data_i[74:74] };
    end 
    if(N7410) begin
      { mem[1033:1033] } <= { data_i[73:73] };
    end 
    if(N7409) begin
      { mem[1032:1032] } <= { data_i[72:72] };
    end 
    if(N7408) begin
      { mem[1031:1031] } <= { data_i[71:71] };
    end 
    if(N7407) begin
      { mem[1030:1030] } <= { data_i[70:70] };
    end 
    if(N7406) begin
      { mem[1029:1029] } <= { data_i[69:69] };
    end 
    if(N7405) begin
      { mem[1028:1028] } <= { data_i[68:68] };
    end 
    if(N7404) begin
      { mem[1027:1027] } <= { data_i[67:67] };
    end 
    if(N7403) begin
      { mem[1026:1026] } <= { data_i[66:66] };
    end 
    if(N7402) begin
      { mem[1025:1025] } <= { data_i[65:65] };
    end 
    if(N7401) begin
      { mem[1024:1024] } <= { data_i[64:64] };
    end 
    if(N7400) begin
      { mem[1023:1023] } <= { data_i[63:63] };
    end 
    if(N7399) begin
      { mem[1022:1022] } <= { data_i[62:62] };
    end 
    if(N7398) begin
      { mem[1021:1021] } <= { data_i[61:61] };
    end 
    if(N7397) begin
      { mem[1020:1020] } <= { data_i[60:60] };
    end 
    if(N7396) begin
      { mem[1019:1019] } <= { data_i[59:59] };
    end 
    if(N7395) begin
      { mem[1018:1018] } <= { data_i[58:58] };
    end 
    if(N7394) begin
      { mem[1017:1017] } <= { data_i[57:57] };
    end 
    if(N7393) begin
      { mem[1016:1016] } <= { data_i[56:56] };
    end 
    if(N7392) begin
      { mem[1015:1015] } <= { data_i[55:55] };
    end 
    if(N7391) begin
      { mem[1014:1014] } <= { data_i[54:54] };
    end 
    if(N7390) begin
      { mem[1013:1013] } <= { data_i[53:53] };
    end 
    if(N7389) begin
      { mem[1012:1012] } <= { data_i[52:52] };
    end 
    if(N7388) begin
      { mem[1011:1011] } <= { data_i[51:51] };
    end 
    if(N7387) begin
      { mem[1010:1010] } <= { data_i[50:50] };
    end 
    if(N7386) begin
      { mem[1009:1009] } <= { data_i[49:49] };
    end 
    if(N7385) begin
      { mem[1008:1008] } <= { data_i[48:48] };
    end 
    if(N7384) begin
      { mem[1007:1007] } <= { data_i[47:47] };
    end 
    if(N7383) begin
      { mem[1006:1006] } <= { data_i[46:46] };
    end 
    if(N7382) begin
      { mem[1005:1005] } <= { data_i[45:45] };
    end 
    if(N7381) begin
      { mem[1004:1004] } <= { data_i[44:44] };
    end 
    if(N7380) begin
      { mem[1003:1003] } <= { data_i[43:43] };
    end 
    if(N7379) begin
      { mem[1002:1002] } <= { data_i[42:42] };
    end 
    if(N7378) begin
      { mem[1001:1001] } <= { data_i[41:41] };
    end 
    if(N7377) begin
      { mem[1000:1000] } <= { data_i[40:40] };
    end 
    if(N7376) begin
      { mem[999:999] } <= { data_i[39:39] };
    end 
    if(N7375) begin
      { mem[998:998] } <= { data_i[38:38] };
    end 
    if(N7374) begin
      { mem[997:997] } <= { data_i[37:37] };
    end 
    if(N7373) begin
      { mem[996:996] } <= { data_i[36:36] };
    end 
    if(N7372) begin
      { mem[995:995] } <= { data_i[35:35] };
    end 
    if(N7371) begin
      { mem[994:994] } <= { data_i[34:34] };
    end 
    if(N7370) begin
      { mem[993:993] } <= { data_i[33:33] };
    end 
    if(N7369) begin
      { mem[992:992] } <= { data_i[32:32] };
    end 
    if(N7368) begin
      { mem[991:991] } <= { data_i[31:31] };
    end 
    if(N7367) begin
      { mem[990:990] } <= { data_i[30:30] };
    end 
    if(N7366) begin
      { mem[989:989] } <= { data_i[29:29] };
    end 
    if(N7365) begin
      { mem[988:988] } <= { data_i[28:28] };
    end 
    if(N7364) begin
      { mem[987:987] } <= { data_i[27:27] };
    end 
    if(N7363) begin
      { mem[986:986] } <= { data_i[26:26] };
    end 
    if(N7362) begin
      { mem[985:985] } <= { data_i[25:25] };
    end 
    if(N7361) begin
      { mem[984:984] } <= { data_i[24:24] };
    end 
    if(N7360) begin
      { mem[983:983] } <= { data_i[23:23] };
    end 
    if(N7359) begin
      { mem[982:982] } <= { data_i[22:22] };
    end 
    if(N7358) begin
      { mem[981:981] } <= { data_i[21:21] };
    end 
    if(N7357) begin
      { mem[980:980] } <= { data_i[20:20] };
    end 
    if(N7356) begin
      { mem[979:979] } <= { data_i[19:19] };
    end 
    if(N7355) begin
      { mem[978:978] } <= { data_i[18:18] };
    end 
    if(N7354) begin
      { mem[977:977] } <= { data_i[17:17] };
    end 
    if(N7353) begin
      { mem[976:976] } <= { data_i[16:16] };
    end 
    if(N7352) begin
      { mem[975:975] } <= { data_i[15:15] };
    end 
    if(N7351) begin
      { mem[974:974] } <= { data_i[14:14] };
    end 
    if(N7350) begin
      { mem[973:973] } <= { data_i[13:13] };
    end 
    if(N7349) begin
      { mem[972:972] } <= { data_i[12:12] };
    end 
    if(N7348) begin
      { mem[971:971] } <= { data_i[11:11] };
    end 
    if(N7347) begin
      { mem[970:970] } <= { data_i[10:10] };
    end 
    if(N7346) begin
      { mem[969:969] } <= { data_i[9:9] };
    end 
    if(N7345) begin
      { mem[968:968] } <= { data_i[8:8] };
    end 
    if(N7344) begin
      { mem[967:967] } <= { data_i[7:7] };
    end 
    if(N7343) begin
      { mem[966:966] } <= { data_i[6:6] };
    end 
    if(N7342) begin
      { mem[965:965] } <= { data_i[5:5] };
    end 
    if(N7341) begin
      { mem[964:964] } <= { data_i[4:4] };
    end 
    if(N7340) begin
      { mem[963:963] } <= { data_i[3:3] };
    end 
    if(N7339) begin
      { mem[962:962] } <= { data_i[2:2] };
    end 
    if(N7338) begin
      { mem[961:961] } <= { data_i[1:1] };
    end 
    if(N7337) begin
      { mem[960:960] } <= { data_i[0:0] };
    end 
    if(N7336) begin
      { mem[959:959] } <= { data_i[79:79] };
    end 
    if(N7335) begin
      { mem[958:958] } <= { data_i[78:78] };
    end 
    if(N7334) begin
      { mem[957:957] } <= { data_i[77:77] };
    end 
    if(N7333) begin
      { mem[956:956] } <= { data_i[76:76] };
    end 
    if(N7332) begin
      { mem[955:955] } <= { data_i[75:75] };
    end 
    if(N7331) begin
      { mem[954:954] } <= { data_i[74:74] };
    end 
    if(N7330) begin
      { mem[953:953] } <= { data_i[73:73] };
    end 
    if(N7329) begin
      { mem[952:952] } <= { data_i[72:72] };
    end 
    if(N7328) begin
      { mem[951:951] } <= { data_i[71:71] };
    end 
    if(N7327) begin
      { mem[950:950] } <= { data_i[70:70] };
    end 
    if(N7326) begin
      { mem[949:949] } <= { data_i[69:69] };
    end 
    if(N7325) begin
      { mem[948:948] } <= { data_i[68:68] };
    end 
    if(N7324) begin
      { mem[947:947] } <= { data_i[67:67] };
    end 
    if(N7323) begin
      { mem[946:946] } <= { data_i[66:66] };
    end 
    if(N7322) begin
      { mem[945:945] } <= { data_i[65:65] };
    end 
    if(N7321) begin
      { mem[944:944] } <= { data_i[64:64] };
    end 
    if(N7320) begin
      { mem[943:943] } <= { data_i[63:63] };
    end 
    if(N7319) begin
      { mem[942:942] } <= { data_i[62:62] };
    end 
    if(N7318) begin
      { mem[941:941] } <= { data_i[61:61] };
    end 
    if(N7317) begin
      { mem[940:940] } <= { data_i[60:60] };
    end 
    if(N7316) begin
      { mem[939:939] } <= { data_i[59:59] };
    end 
    if(N7315) begin
      { mem[938:938] } <= { data_i[58:58] };
    end 
    if(N7314) begin
      { mem[937:937] } <= { data_i[57:57] };
    end 
    if(N7313) begin
      { mem[936:936] } <= { data_i[56:56] };
    end 
    if(N7312) begin
      { mem[935:935] } <= { data_i[55:55] };
    end 
    if(N7311) begin
      { mem[934:934] } <= { data_i[54:54] };
    end 
    if(N7310) begin
      { mem[933:933] } <= { data_i[53:53] };
    end 
    if(N7309) begin
      { mem[932:932] } <= { data_i[52:52] };
    end 
    if(N7308) begin
      { mem[931:931] } <= { data_i[51:51] };
    end 
    if(N7307) begin
      { mem[930:930] } <= { data_i[50:50] };
    end 
    if(N7306) begin
      { mem[929:929] } <= { data_i[49:49] };
    end 
    if(N7305) begin
      { mem[928:928] } <= { data_i[48:48] };
    end 
    if(N7304) begin
      { mem[927:927] } <= { data_i[47:47] };
    end 
    if(N7303) begin
      { mem[926:926] } <= { data_i[46:46] };
    end 
    if(N7302) begin
      { mem[925:925] } <= { data_i[45:45] };
    end 
    if(N7301) begin
      { mem[924:924] } <= { data_i[44:44] };
    end 
    if(N7300) begin
      { mem[923:923] } <= { data_i[43:43] };
    end 
    if(N7299) begin
      { mem[922:922] } <= { data_i[42:42] };
    end 
    if(N7298) begin
      { mem[921:921] } <= { data_i[41:41] };
    end 
    if(N7297) begin
      { mem[920:920] } <= { data_i[40:40] };
    end 
    if(N7296) begin
      { mem[919:919] } <= { data_i[39:39] };
    end 
    if(N7295) begin
      { mem[918:918] } <= { data_i[38:38] };
    end 
    if(N7294) begin
      { mem[917:917] } <= { data_i[37:37] };
    end 
    if(N7293) begin
      { mem[916:916] } <= { data_i[36:36] };
    end 
    if(N7292) begin
      { mem[915:915] } <= { data_i[35:35] };
    end 
    if(N7291) begin
      { mem[914:914] } <= { data_i[34:34] };
    end 
    if(N7290) begin
      { mem[913:913] } <= { data_i[33:33] };
    end 
    if(N7289) begin
      { mem[912:912] } <= { data_i[32:32] };
    end 
    if(N7288) begin
      { mem[911:911] } <= { data_i[31:31] };
    end 
    if(N7287) begin
      { mem[910:910] } <= { data_i[30:30] };
    end 
    if(N7286) begin
      { mem[909:909] } <= { data_i[29:29] };
    end 
    if(N7285) begin
      { mem[908:908] } <= { data_i[28:28] };
    end 
    if(N7284) begin
      { mem[907:907] } <= { data_i[27:27] };
    end 
    if(N7283) begin
      { mem[906:906] } <= { data_i[26:26] };
    end 
    if(N7282) begin
      { mem[905:905] } <= { data_i[25:25] };
    end 
    if(N7281) begin
      { mem[904:904] } <= { data_i[24:24] };
    end 
    if(N7280) begin
      { mem[903:903] } <= { data_i[23:23] };
    end 
    if(N7279) begin
      { mem[902:902] } <= { data_i[22:22] };
    end 
    if(N7278) begin
      { mem[901:901] } <= { data_i[21:21] };
    end 
    if(N7277) begin
      { mem[900:900] } <= { data_i[20:20] };
    end 
    if(N7276) begin
      { mem[899:899] } <= { data_i[19:19] };
    end 
    if(N7275) begin
      { mem[898:898] } <= { data_i[18:18] };
    end 
    if(N7274) begin
      { mem[897:897] } <= { data_i[17:17] };
    end 
    if(N7273) begin
      { mem[896:896] } <= { data_i[16:16] };
    end 
    if(N7272) begin
      { mem[895:895] } <= { data_i[15:15] };
    end 
    if(N7271) begin
      { mem[894:894] } <= { data_i[14:14] };
    end 
    if(N7270) begin
      { mem[893:893] } <= { data_i[13:13] };
    end 
    if(N7269) begin
      { mem[892:892] } <= { data_i[12:12] };
    end 
    if(N7268) begin
      { mem[891:891] } <= { data_i[11:11] };
    end 
    if(N7267) begin
      { mem[890:890] } <= { data_i[10:10] };
    end 
    if(N7266) begin
      { mem[889:889] } <= { data_i[9:9] };
    end 
    if(N7265) begin
      { mem[888:888] } <= { data_i[8:8] };
    end 
    if(N7264) begin
      { mem[887:887] } <= { data_i[7:7] };
    end 
    if(N7263) begin
      { mem[886:886] } <= { data_i[6:6] };
    end 
    if(N7262) begin
      { mem[885:885] } <= { data_i[5:5] };
    end 
    if(N7261) begin
      { mem[884:884] } <= { data_i[4:4] };
    end 
    if(N7260) begin
      { mem[883:883] } <= { data_i[3:3] };
    end 
    if(N7259) begin
      { mem[882:882] } <= { data_i[2:2] };
    end 
    if(N7258) begin
      { mem[881:881] } <= { data_i[1:1] };
    end 
    if(N7257) begin
      { mem[880:880] } <= { data_i[0:0] };
    end 
    if(N7256) begin
      { mem[879:879] } <= { data_i[79:79] };
    end 
    if(N7255) begin
      { mem[878:878] } <= { data_i[78:78] };
    end 
    if(N7254) begin
      { mem[877:877] } <= { data_i[77:77] };
    end 
    if(N7253) begin
      { mem[876:876] } <= { data_i[76:76] };
    end 
    if(N7252) begin
      { mem[875:875] } <= { data_i[75:75] };
    end 
    if(N7251) begin
      { mem[874:874] } <= { data_i[74:74] };
    end 
    if(N7250) begin
      { mem[873:873] } <= { data_i[73:73] };
    end 
    if(N7249) begin
      { mem[872:872] } <= { data_i[72:72] };
    end 
    if(N7248) begin
      { mem[871:871] } <= { data_i[71:71] };
    end 
    if(N7247) begin
      { mem[870:870] } <= { data_i[70:70] };
    end 
    if(N7246) begin
      { mem[869:869] } <= { data_i[69:69] };
    end 
    if(N7245) begin
      { mem[868:868] } <= { data_i[68:68] };
    end 
    if(N7244) begin
      { mem[867:867] } <= { data_i[67:67] };
    end 
    if(N7243) begin
      { mem[866:866] } <= { data_i[66:66] };
    end 
    if(N7242) begin
      { mem[865:865] } <= { data_i[65:65] };
    end 
    if(N7241) begin
      { mem[864:864] } <= { data_i[64:64] };
    end 
    if(N7240) begin
      { mem[863:863] } <= { data_i[63:63] };
    end 
    if(N7239) begin
      { mem[862:862] } <= { data_i[62:62] };
    end 
    if(N7238) begin
      { mem[861:861] } <= { data_i[61:61] };
    end 
    if(N7237) begin
      { mem[860:860] } <= { data_i[60:60] };
    end 
    if(N7236) begin
      { mem[859:859] } <= { data_i[59:59] };
    end 
    if(N7235) begin
      { mem[858:858] } <= { data_i[58:58] };
    end 
    if(N7234) begin
      { mem[857:857] } <= { data_i[57:57] };
    end 
    if(N7233) begin
      { mem[856:856] } <= { data_i[56:56] };
    end 
    if(N7232) begin
      { mem[855:855] } <= { data_i[55:55] };
    end 
    if(N7231) begin
      { mem[854:854] } <= { data_i[54:54] };
    end 
    if(N7230) begin
      { mem[853:853] } <= { data_i[53:53] };
    end 
    if(N7229) begin
      { mem[852:852] } <= { data_i[52:52] };
    end 
    if(N7228) begin
      { mem[851:851] } <= { data_i[51:51] };
    end 
    if(N7227) begin
      { mem[850:850] } <= { data_i[50:50] };
    end 
    if(N7226) begin
      { mem[849:849] } <= { data_i[49:49] };
    end 
    if(N7225) begin
      { mem[848:848] } <= { data_i[48:48] };
    end 
    if(N7224) begin
      { mem[847:847] } <= { data_i[47:47] };
    end 
    if(N7223) begin
      { mem[846:846] } <= { data_i[46:46] };
    end 
    if(N7222) begin
      { mem[845:845] } <= { data_i[45:45] };
    end 
    if(N7221) begin
      { mem[844:844] } <= { data_i[44:44] };
    end 
    if(N7220) begin
      { mem[843:843] } <= { data_i[43:43] };
    end 
    if(N7219) begin
      { mem[842:842] } <= { data_i[42:42] };
    end 
    if(N7218) begin
      { mem[841:841] } <= { data_i[41:41] };
    end 
    if(N7217) begin
      { mem[840:840] } <= { data_i[40:40] };
    end 
    if(N7216) begin
      { mem[839:839] } <= { data_i[39:39] };
    end 
    if(N7215) begin
      { mem[838:838] } <= { data_i[38:38] };
    end 
    if(N7214) begin
      { mem[837:837] } <= { data_i[37:37] };
    end 
    if(N7213) begin
      { mem[836:836] } <= { data_i[36:36] };
    end 
    if(N7212) begin
      { mem[835:835] } <= { data_i[35:35] };
    end 
    if(N7211) begin
      { mem[834:834] } <= { data_i[34:34] };
    end 
    if(N7210) begin
      { mem[833:833] } <= { data_i[33:33] };
    end 
    if(N7209) begin
      { mem[832:832] } <= { data_i[32:32] };
    end 
    if(N7208) begin
      { mem[831:831] } <= { data_i[31:31] };
    end 
    if(N7207) begin
      { mem[830:830] } <= { data_i[30:30] };
    end 
    if(N7206) begin
      { mem[829:829] } <= { data_i[29:29] };
    end 
    if(N7205) begin
      { mem[828:828] } <= { data_i[28:28] };
    end 
    if(N7204) begin
      { mem[827:827] } <= { data_i[27:27] };
    end 
    if(N7203) begin
      { mem[826:826] } <= { data_i[26:26] };
    end 
    if(N7202) begin
      { mem[825:825] } <= { data_i[25:25] };
    end 
    if(N7201) begin
      { mem[824:824] } <= { data_i[24:24] };
    end 
    if(N7200) begin
      { mem[823:823] } <= { data_i[23:23] };
    end 
    if(N7199) begin
      { mem[822:822] } <= { data_i[22:22] };
    end 
    if(N7198) begin
      { mem[821:821] } <= { data_i[21:21] };
    end 
    if(N7197) begin
      { mem[820:820] } <= { data_i[20:20] };
    end 
    if(N7196) begin
      { mem[819:819] } <= { data_i[19:19] };
    end 
    if(N7195) begin
      { mem[818:818] } <= { data_i[18:18] };
    end 
    if(N7194) begin
      { mem[817:817] } <= { data_i[17:17] };
    end 
    if(N7193) begin
      { mem[816:816] } <= { data_i[16:16] };
    end 
    if(N7192) begin
      { mem[815:815] } <= { data_i[15:15] };
    end 
    if(N7191) begin
      { mem[814:814] } <= { data_i[14:14] };
    end 
    if(N7190) begin
      { mem[813:813] } <= { data_i[13:13] };
    end 
    if(N7189) begin
      { mem[812:812] } <= { data_i[12:12] };
    end 
    if(N7188) begin
      { mem[811:811] } <= { data_i[11:11] };
    end 
    if(N7187) begin
      { mem[810:810] } <= { data_i[10:10] };
    end 
    if(N7186) begin
      { mem[809:809] } <= { data_i[9:9] };
    end 
    if(N7185) begin
      { mem[808:808] } <= { data_i[8:8] };
    end 
    if(N7184) begin
      { mem[807:807] } <= { data_i[7:7] };
    end 
    if(N7183) begin
      { mem[806:806] } <= { data_i[6:6] };
    end 
    if(N7182) begin
      { mem[805:805] } <= { data_i[5:5] };
    end 
    if(N7181) begin
      { mem[804:804] } <= { data_i[4:4] };
    end 
    if(N7180) begin
      { mem[803:803] } <= { data_i[3:3] };
    end 
    if(N7179) begin
      { mem[802:802] } <= { data_i[2:2] };
    end 
    if(N7178) begin
      { mem[801:801] } <= { data_i[1:1] };
    end 
    if(N7177) begin
      { mem[800:800] } <= { data_i[0:0] };
    end 
    if(N7176) begin
      { mem[799:799] } <= { data_i[79:79] };
    end 
    if(N7175) begin
      { mem[798:798] } <= { data_i[78:78] };
    end 
    if(N7174) begin
      { mem[797:797] } <= { data_i[77:77] };
    end 
    if(N7173) begin
      { mem[796:796] } <= { data_i[76:76] };
    end 
    if(N7172) begin
      { mem[795:795] } <= { data_i[75:75] };
    end 
    if(N7171) begin
      { mem[794:794] } <= { data_i[74:74] };
    end 
    if(N7170) begin
      { mem[793:793] } <= { data_i[73:73] };
    end 
    if(N7169) begin
      { mem[792:792] } <= { data_i[72:72] };
    end 
    if(N7168) begin
      { mem[791:791] } <= { data_i[71:71] };
    end 
    if(N7167) begin
      { mem[790:790] } <= { data_i[70:70] };
    end 
    if(N7166) begin
      { mem[789:789] } <= { data_i[69:69] };
    end 
    if(N7165) begin
      { mem[788:788] } <= { data_i[68:68] };
    end 
    if(N7164) begin
      { mem[787:787] } <= { data_i[67:67] };
    end 
    if(N7163) begin
      { mem[786:786] } <= { data_i[66:66] };
    end 
    if(N7162) begin
      { mem[785:785] } <= { data_i[65:65] };
    end 
    if(N7161) begin
      { mem[784:784] } <= { data_i[64:64] };
    end 
    if(N7160) begin
      { mem[783:783] } <= { data_i[63:63] };
    end 
    if(N7159) begin
      { mem[782:782] } <= { data_i[62:62] };
    end 
    if(N7158) begin
      { mem[781:781] } <= { data_i[61:61] };
    end 
    if(N7157) begin
      { mem[780:780] } <= { data_i[60:60] };
    end 
    if(N7156) begin
      { mem[779:779] } <= { data_i[59:59] };
    end 
    if(N7155) begin
      { mem[778:778] } <= { data_i[58:58] };
    end 
    if(N7154) begin
      { mem[777:777] } <= { data_i[57:57] };
    end 
    if(N7153) begin
      { mem[776:776] } <= { data_i[56:56] };
    end 
    if(N7152) begin
      { mem[775:775] } <= { data_i[55:55] };
    end 
    if(N7151) begin
      { mem[774:774] } <= { data_i[54:54] };
    end 
    if(N7150) begin
      { mem[773:773] } <= { data_i[53:53] };
    end 
    if(N7149) begin
      { mem[772:772] } <= { data_i[52:52] };
    end 
    if(N7148) begin
      { mem[771:771] } <= { data_i[51:51] };
    end 
    if(N7147) begin
      { mem[770:770] } <= { data_i[50:50] };
    end 
    if(N7146) begin
      { mem[769:769] } <= { data_i[49:49] };
    end 
    if(N7145) begin
      { mem[768:768] } <= { data_i[48:48] };
    end 
    if(N7144) begin
      { mem[767:767] } <= { data_i[47:47] };
    end 
    if(N7143) begin
      { mem[766:766] } <= { data_i[46:46] };
    end 
    if(N7142) begin
      { mem[765:765] } <= { data_i[45:45] };
    end 
    if(N7141) begin
      { mem[764:764] } <= { data_i[44:44] };
    end 
    if(N7140) begin
      { mem[763:763] } <= { data_i[43:43] };
    end 
    if(N7139) begin
      { mem[762:762] } <= { data_i[42:42] };
    end 
    if(N7138) begin
      { mem[761:761] } <= { data_i[41:41] };
    end 
    if(N7137) begin
      { mem[760:760] } <= { data_i[40:40] };
    end 
    if(N7136) begin
      { mem[759:759] } <= { data_i[39:39] };
    end 
    if(N7135) begin
      { mem[758:758] } <= { data_i[38:38] };
    end 
    if(N7134) begin
      { mem[757:757] } <= { data_i[37:37] };
    end 
    if(N7133) begin
      { mem[756:756] } <= { data_i[36:36] };
    end 
    if(N7132) begin
      { mem[755:755] } <= { data_i[35:35] };
    end 
    if(N7131) begin
      { mem[754:754] } <= { data_i[34:34] };
    end 
    if(N7130) begin
      { mem[753:753] } <= { data_i[33:33] };
    end 
    if(N7129) begin
      { mem[752:752] } <= { data_i[32:32] };
    end 
    if(N7128) begin
      { mem[751:751] } <= { data_i[31:31] };
    end 
    if(N7127) begin
      { mem[750:750] } <= { data_i[30:30] };
    end 
    if(N7126) begin
      { mem[749:749] } <= { data_i[29:29] };
    end 
    if(N7125) begin
      { mem[748:748] } <= { data_i[28:28] };
    end 
    if(N7124) begin
      { mem[747:747] } <= { data_i[27:27] };
    end 
    if(N7123) begin
      { mem[746:746] } <= { data_i[26:26] };
    end 
    if(N7122) begin
      { mem[745:745] } <= { data_i[25:25] };
    end 
    if(N7121) begin
      { mem[744:744] } <= { data_i[24:24] };
    end 
    if(N7120) begin
      { mem[743:743] } <= { data_i[23:23] };
    end 
    if(N7119) begin
      { mem[742:742] } <= { data_i[22:22] };
    end 
    if(N7118) begin
      { mem[741:741] } <= { data_i[21:21] };
    end 
    if(N7117) begin
      { mem[740:740] } <= { data_i[20:20] };
    end 
    if(N7116) begin
      { mem[739:739] } <= { data_i[19:19] };
    end 
    if(N7115) begin
      { mem[738:738] } <= { data_i[18:18] };
    end 
    if(N7114) begin
      { mem[737:737] } <= { data_i[17:17] };
    end 
    if(N7113) begin
      { mem[736:736] } <= { data_i[16:16] };
    end 
    if(N7112) begin
      { mem[735:735] } <= { data_i[15:15] };
    end 
    if(N7111) begin
      { mem[734:734] } <= { data_i[14:14] };
    end 
    if(N7110) begin
      { mem[733:733] } <= { data_i[13:13] };
    end 
    if(N7109) begin
      { mem[732:732] } <= { data_i[12:12] };
    end 
    if(N7108) begin
      { mem[731:731] } <= { data_i[11:11] };
    end 
    if(N7107) begin
      { mem[730:730] } <= { data_i[10:10] };
    end 
    if(N7106) begin
      { mem[729:729] } <= { data_i[9:9] };
    end 
    if(N7105) begin
      { mem[728:728] } <= { data_i[8:8] };
    end 
    if(N7104) begin
      { mem[727:727] } <= { data_i[7:7] };
    end 
    if(N7103) begin
      { mem[726:726] } <= { data_i[6:6] };
    end 
    if(N7102) begin
      { mem[725:725] } <= { data_i[5:5] };
    end 
    if(N7101) begin
      { mem[724:724] } <= { data_i[4:4] };
    end 
    if(N7100) begin
      { mem[723:723] } <= { data_i[3:3] };
    end 
    if(N7099) begin
      { mem[722:722] } <= { data_i[2:2] };
    end 
    if(N7098) begin
      { mem[721:721] } <= { data_i[1:1] };
    end 
    if(N7097) begin
      { mem[720:720] } <= { data_i[0:0] };
    end 
    if(N7096) begin
      { mem[719:719] } <= { data_i[79:79] };
    end 
    if(N7095) begin
      { mem[718:718] } <= { data_i[78:78] };
    end 
    if(N7094) begin
      { mem[717:717] } <= { data_i[77:77] };
    end 
    if(N7093) begin
      { mem[716:716] } <= { data_i[76:76] };
    end 
    if(N7092) begin
      { mem[715:715] } <= { data_i[75:75] };
    end 
    if(N7091) begin
      { mem[714:714] } <= { data_i[74:74] };
    end 
    if(N7090) begin
      { mem[713:713] } <= { data_i[73:73] };
    end 
    if(N7089) begin
      { mem[712:712] } <= { data_i[72:72] };
    end 
    if(N7088) begin
      { mem[711:711] } <= { data_i[71:71] };
    end 
    if(N7087) begin
      { mem[710:710] } <= { data_i[70:70] };
    end 
    if(N7086) begin
      { mem[709:709] } <= { data_i[69:69] };
    end 
    if(N7085) begin
      { mem[708:708] } <= { data_i[68:68] };
    end 
    if(N7084) begin
      { mem[707:707] } <= { data_i[67:67] };
    end 
    if(N7083) begin
      { mem[706:706] } <= { data_i[66:66] };
    end 
    if(N7082) begin
      { mem[705:705] } <= { data_i[65:65] };
    end 
    if(N7081) begin
      { mem[704:704] } <= { data_i[64:64] };
    end 
    if(N7080) begin
      { mem[703:703] } <= { data_i[63:63] };
    end 
    if(N7079) begin
      { mem[702:702] } <= { data_i[62:62] };
    end 
    if(N7078) begin
      { mem[701:701] } <= { data_i[61:61] };
    end 
    if(N7077) begin
      { mem[700:700] } <= { data_i[60:60] };
    end 
    if(N7076) begin
      { mem[699:699] } <= { data_i[59:59] };
    end 
    if(N7075) begin
      { mem[698:698] } <= { data_i[58:58] };
    end 
    if(N7074) begin
      { mem[697:697] } <= { data_i[57:57] };
    end 
    if(N7073) begin
      { mem[696:696] } <= { data_i[56:56] };
    end 
    if(N7072) begin
      { mem[695:695] } <= { data_i[55:55] };
    end 
    if(N7071) begin
      { mem[694:694] } <= { data_i[54:54] };
    end 
    if(N7070) begin
      { mem[693:693] } <= { data_i[53:53] };
    end 
    if(N7069) begin
      { mem[692:692] } <= { data_i[52:52] };
    end 
    if(N7068) begin
      { mem[691:691] } <= { data_i[51:51] };
    end 
    if(N7067) begin
      { mem[690:690] } <= { data_i[50:50] };
    end 
    if(N7066) begin
      { mem[689:689] } <= { data_i[49:49] };
    end 
    if(N7065) begin
      { mem[688:688] } <= { data_i[48:48] };
    end 
    if(N7064) begin
      { mem[687:687] } <= { data_i[47:47] };
    end 
    if(N7063) begin
      { mem[686:686] } <= { data_i[46:46] };
    end 
    if(N7062) begin
      { mem[685:685] } <= { data_i[45:45] };
    end 
    if(N7061) begin
      { mem[684:684] } <= { data_i[44:44] };
    end 
    if(N7060) begin
      { mem[683:683] } <= { data_i[43:43] };
    end 
    if(N7059) begin
      { mem[682:682] } <= { data_i[42:42] };
    end 
    if(N7058) begin
      { mem[681:681] } <= { data_i[41:41] };
    end 
    if(N7057) begin
      { mem[680:680] } <= { data_i[40:40] };
    end 
    if(N7056) begin
      { mem[679:679] } <= { data_i[39:39] };
    end 
    if(N7055) begin
      { mem[678:678] } <= { data_i[38:38] };
    end 
    if(N7054) begin
      { mem[677:677] } <= { data_i[37:37] };
    end 
    if(N7053) begin
      { mem[676:676] } <= { data_i[36:36] };
    end 
    if(N7052) begin
      { mem[675:675] } <= { data_i[35:35] };
    end 
    if(N7051) begin
      { mem[674:674] } <= { data_i[34:34] };
    end 
    if(N7050) begin
      { mem[673:673] } <= { data_i[33:33] };
    end 
    if(N7049) begin
      { mem[672:672] } <= { data_i[32:32] };
    end 
    if(N7048) begin
      { mem[671:671] } <= { data_i[31:31] };
    end 
    if(N7047) begin
      { mem[670:670] } <= { data_i[30:30] };
    end 
    if(N7046) begin
      { mem[669:669] } <= { data_i[29:29] };
    end 
    if(N7045) begin
      { mem[668:668] } <= { data_i[28:28] };
    end 
    if(N7044) begin
      { mem[667:667] } <= { data_i[27:27] };
    end 
    if(N7043) begin
      { mem[666:666] } <= { data_i[26:26] };
    end 
    if(N7042) begin
      { mem[665:665] } <= { data_i[25:25] };
    end 
    if(N7041) begin
      { mem[664:664] } <= { data_i[24:24] };
    end 
    if(N7040) begin
      { mem[663:663] } <= { data_i[23:23] };
    end 
    if(N7039) begin
      { mem[662:662] } <= { data_i[22:22] };
    end 
    if(N7038) begin
      { mem[661:661] } <= { data_i[21:21] };
    end 
    if(N7037) begin
      { mem[660:660] } <= { data_i[20:20] };
    end 
    if(N7036) begin
      { mem[659:659] } <= { data_i[19:19] };
    end 
    if(N7035) begin
      { mem[658:658] } <= { data_i[18:18] };
    end 
    if(N7034) begin
      { mem[657:657] } <= { data_i[17:17] };
    end 
    if(N7033) begin
      { mem[656:656] } <= { data_i[16:16] };
    end 
    if(N7032) begin
      { mem[655:655] } <= { data_i[15:15] };
    end 
    if(N7031) begin
      { mem[654:654] } <= { data_i[14:14] };
    end 
    if(N7030) begin
      { mem[653:653] } <= { data_i[13:13] };
    end 
    if(N7029) begin
      { mem[652:652] } <= { data_i[12:12] };
    end 
    if(N7028) begin
      { mem[651:651] } <= { data_i[11:11] };
    end 
    if(N7027) begin
      { mem[650:650] } <= { data_i[10:10] };
    end 
    if(N7026) begin
      { mem[649:649] } <= { data_i[9:9] };
    end 
    if(N7025) begin
      { mem[648:648] } <= { data_i[8:8] };
    end 
    if(N7024) begin
      { mem[647:647] } <= { data_i[7:7] };
    end 
    if(N7023) begin
      { mem[646:646] } <= { data_i[6:6] };
    end 
    if(N7022) begin
      { mem[645:645] } <= { data_i[5:5] };
    end 
    if(N7021) begin
      { mem[644:644] } <= { data_i[4:4] };
    end 
    if(N7020) begin
      { mem[643:643] } <= { data_i[3:3] };
    end 
    if(N7019) begin
      { mem[642:642] } <= { data_i[2:2] };
    end 
    if(N7018) begin
      { mem[641:641] } <= { data_i[1:1] };
    end 
    if(N7017) begin
      { mem[640:640] } <= { data_i[0:0] };
    end 
    if(N7016) begin
      { mem[639:639] } <= { data_i[79:79] };
    end 
    if(N7015) begin
      { mem[638:638] } <= { data_i[78:78] };
    end 
    if(N7014) begin
      { mem[637:637] } <= { data_i[77:77] };
    end 
    if(N7013) begin
      { mem[636:636] } <= { data_i[76:76] };
    end 
    if(N7012) begin
      { mem[635:635] } <= { data_i[75:75] };
    end 
    if(N7011) begin
      { mem[634:634] } <= { data_i[74:74] };
    end 
    if(N7010) begin
      { mem[633:633] } <= { data_i[73:73] };
    end 
    if(N7009) begin
      { mem[632:632] } <= { data_i[72:72] };
    end 
    if(N7008) begin
      { mem[631:631] } <= { data_i[71:71] };
    end 
    if(N7007) begin
      { mem[630:630] } <= { data_i[70:70] };
    end 
    if(N7006) begin
      { mem[629:629] } <= { data_i[69:69] };
    end 
    if(N7005) begin
      { mem[628:628] } <= { data_i[68:68] };
    end 
    if(N7004) begin
      { mem[627:627] } <= { data_i[67:67] };
    end 
    if(N7003) begin
      { mem[626:626] } <= { data_i[66:66] };
    end 
    if(N7002) begin
      { mem[625:625] } <= { data_i[65:65] };
    end 
    if(N7001) begin
      { mem[624:624] } <= { data_i[64:64] };
    end 
    if(N7000) begin
      { mem[623:623] } <= { data_i[63:63] };
    end 
    if(N6999) begin
      { mem[622:622] } <= { data_i[62:62] };
    end 
    if(N6998) begin
      { mem[621:621] } <= { data_i[61:61] };
    end 
    if(N6997) begin
      { mem[620:620] } <= { data_i[60:60] };
    end 
    if(N6996) begin
      { mem[619:619] } <= { data_i[59:59] };
    end 
    if(N6995) begin
      { mem[618:618] } <= { data_i[58:58] };
    end 
    if(N6994) begin
      { mem[617:617] } <= { data_i[57:57] };
    end 
    if(N6993) begin
      { mem[616:616] } <= { data_i[56:56] };
    end 
    if(N6992) begin
      { mem[615:615] } <= { data_i[55:55] };
    end 
    if(N6991) begin
      { mem[614:614] } <= { data_i[54:54] };
    end 
    if(N6990) begin
      { mem[613:613] } <= { data_i[53:53] };
    end 
    if(N6989) begin
      { mem[612:612] } <= { data_i[52:52] };
    end 
    if(N6988) begin
      { mem[611:611] } <= { data_i[51:51] };
    end 
    if(N6987) begin
      { mem[610:610] } <= { data_i[50:50] };
    end 
    if(N6986) begin
      { mem[609:609] } <= { data_i[49:49] };
    end 
    if(N6985) begin
      { mem[608:608] } <= { data_i[48:48] };
    end 
    if(N6984) begin
      { mem[607:607] } <= { data_i[47:47] };
    end 
    if(N6983) begin
      { mem[606:606] } <= { data_i[46:46] };
    end 
    if(N6982) begin
      { mem[605:605] } <= { data_i[45:45] };
    end 
    if(N6981) begin
      { mem[604:604] } <= { data_i[44:44] };
    end 
    if(N6980) begin
      { mem[603:603] } <= { data_i[43:43] };
    end 
    if(N6979) begin
      { mem[602:602] } <= { data_i[42:42] };
    end 
    if(N6978) begin
      { mem[601:601] } <= { data_i[41:41] };
    end 
    if(N6977) begin
      { mem[600:600] } <= { data_i[40:40] };
    end 
    if(N6976) begin
      { mem[599:599] } <= { data_i[39:39] };
    end 
    if(N6975) begin
      { mem[598:598] } <= { data_i[38:38] };
    end 
    if(N6974) begin
      { mem[597:597] } <= { data_i[37:37] };
    end 
    if(N6973) begin
      { mem[596:596] } <= { data_i[36:36] };
    end 
    if(N6972) begin
      { mem[595:595] } <= { data_i[35:35] };
    end 
    if(N6971) begin
      { mem[594:594] } <= { data_i[34:34] };
    end 
    if(N6970) begin
      { mem[593:593] } <= { data_i[33:33] };
    end 
    if(N6969) begin
      { mem[592:592] } <= { data_i[32:32] };
    end 
    if(N6968) begin
      { mem[591:591] } <= { data_i[31:31] };
    end 
    if(N6967) begin
      { mem[590:590] } <= { data_i[30:30] };
    end 
    if(N6966) begin
      { mem[589:589] } <= { data_i[29:29] };
    end 
    if(N6965) begin
      { mem[588:588] } <= { data_i[28:28] };
    end 
    if(N6964) begin
      { mem[587:587] } <= { data_i[27:27] };
    end 
    if(N6963) begin
      { mem[586:586] } <= { data_i[26:26] };
    end 
    if(N6962) begin
      { mem[585:585] } <= { data_i[25:25] };
    end 
    if(N6961) begin
      { mem[584:584] } <= { data_i[24:24] };
    end 
    if(N6960) begin
      { mem[583:583] } <= { data_i[23:23] };
    end 
    if(N6959) begin
      { mem[582:582] } <= { data_i[22:22] };
    end 
    if(N6958) begin
      { mem[581:581] } <= { data_i[21:21] };
    end 
    if(N6957) begin
      { mem[580:580] } <= { data_i[20:20] };
    end 
    if(N6956) begin
      { mem[579:579] } <= { data_i[19:19] };
    end 
    if(N6955) begin
      { mem[578:578] } <= { data_i[18:18] };
    end 
    if(N6954) begin
      { mem[577:577] } <= { data_i[17:17] };
    end 
    if(N6953) begin
      { mem[576:576] } <= { data_i[16:16] };
    end 
    if(N6952) begin
      { mem[575:575] } <= { data_i[15:15] };
    end 
    if(N6951) begin
      { mem[574:574] } <= { data_i[14:14] };
    end 
    if(N6950) begin
      { mem[573:573] } <= { data_i[13:13] };
    end 
    if(N6949) begin
      { mem[572:572] } <= { data_i[12:12] };
    end 
    if(N6948) begin
      { mem[571:571] } <= { data_i[11:11] };
    end 
    if(N6947) begin
      { mem[570:570] } <= { data_i[10:10] };
    end 
    if(N6946) begin
      { mem[569:569] } <= { data_i[9:9] };
    end 
    if(N6945) begin
      { mem[568:568] } <= { data_i[8:8] };
    end 
    if(N6944) begin
      { mem[567:567] } <= { data_i[7:7] };
    end 
    if(N6943) begin
      { mem[566:566] } <= { data_i[6:6] };
    end 
    if(N6942) begin
      { mem[565:565] } <= { data_i[5:5] };
    end 
    if(N6941) begin
      { mem[564:564] } <= { data_i[4:4] };
    end 
    if(N6940) begin
      { mem[563:563] } <= { data_i[3:3] };
    end 
    if(N6939) begin
      { mem[562:562] } <= { data_i[2:2] };
    end 
    if(N6938) begin
      { mem[561:561] } <= { data_i[1:1] };
    end 
    if(N6937) begin
      { mem[560:560] } <= { data_i[0:0] };
    end 
    if(N6936) begin
      { mem[559:559] } <= { data_i[79:79] };
    end 
    if(N6935) begin
      { mem[558:558] } <= { data_i[78:78] };
    end 
    if(N6934) begin
      { mem[557:557] } <= { data_i[77:77] };
    end 
    if(N6933) begin
      { mem[556:556] } <= { data_i[76:76] };
    end 
    if(N6932) begin
      { mem[555:555] } <= { data_i[75:75] };
    end 
    if(N6931) begin
      { mem[554:554] } <= { data_i[74:74] };
    end 
    if(N6930) begin
      { mem[553:553] } <= { data_i[73:73] };
    end 
    if(N6929) begin
      { mem[552:552] } <= { data_i[72:72] };
    end 
    if(N6928) begin
      { mem[551:551] } <= { data_i[71:71] };
    end 
    if(N6927) begin
      { mem[550:550] } <= { data_i[70:70] };
    end 
    if(N6926) begin
      { mem[549:549] } <= { data_i[69:69] };
    end 
    if(N6925) begin
      { mem[548:548] } <= { data_i[68:68] };
    end 
    if(N6924) begin
      { mem[547:547] } <= { data_i[67:67] };
    end 
    if(N6923) begin
      { mem[546:546] } <= { data_i[66:66] };
    end 
    if(N6922) begin
      { mem[545:545] } <= { data_i[65:65] };
    end 
    if(N6921) begin
      { mem[544:544] } <= { data_i[64:64] };
    end 
    if(N6920) begin
      { mem[543:543] } <= { data_i[63:63] };
    end 
    if(N6919) begin
      { mem[542:542] } <= { data_i[62:62] };
    end 
    if(N6918) begin
      { mem[541:541] } <= { data_i[61:61] };
    end 
    if(N6917) begin
      { mem[540:540] } <= { data_i[60:60] };
    end 
    if(N6916) begin
      { mem[539:539] } <= { data_i[59:59] };
    end 
    if(N6915) begin
      { mem[538:538] } <= { data_i[58:58] };
    end 
    if(N6914) begin
      { mem[537:537] } <= { data_i[57:57] };
    end 
    if(N6913) begin
      { mem[536:536] } <= { data_i[56:56] };
    end 
    if(N6912) begin
      { mem[535:535] } <= { data_i[55:55] };
    end 
    if(N6911) begin
      { mem[534:534] } <= { data_i[54:54] };
    end 
    if(N6910) begin
      { mem[533:533] } <= { data_i[53:53] };
    end 
    if(N6909) begin
      { mem[532:532] } <= { data_i[52:52] };
    end 
    if(N6908) begin
      { mem[531:531] } <= { data_i[51:51] };
    end 
    if(N6907) begin
      { mem[530:530] } <= { data_i[50:50] };
    end 
    if(N6906) begin
      { mem[529:529] } <= { data_i[49:49] };
    end 
    if(N6905) begin
      { mem[528:528] } <= { data_i[48:48] };
    end 
    if(N6904) begin
      { mem[527:527] } <= { data_i[47:47] };
    end 
    if(N6903) begin
      { mem[526:526] } <= { data_i[46:46] };
    end 
    if(N6902) begin
      { mem[525:525] } <= { data_i[45:45] };
    end 
    if(N6901) begin
      { mem[524:524] } <= { data_i[44:44] };
    end 
    if(N6900) begin
      { mem[523:523] } <= { data_i[43:43] };
    end 
    if(N6899) begin
      { mem[522:522] } <= { data_i[42:42] };
    end 
    if(N6898) begin
      { mem[521:521] } <= { data_i[41:41] };
    end 
    if(N6897) begin
      { mem[520:520] } <= { data_i[40:40] };
    end 
    if(N6896) begin
      { mem[519:519] } <= { data_i[39:39] };
    end 
    if(N6895) begin
      { mem[518:518] } <= { data_i[38:38] };
    end 
    if(N6894) begin
      { mem[517:517] } <= { data_i[37:37] };
    end 
    if(N6893) begin
      { mem[516:516] } <= { data_i[36:36] };
    end 
    if(N6892) begin
      { mem[515:515] } <= { data_i[35:35] };
    end 
    if(N6891) begin
      { mem[514:514] } <= { data_i[34:34] };
    end 
    if(N6890) begin
      { mem[513:513] } <= { data_i[33:33] };
    end 
    if(N6889) begin
      { mem[512:512] } <= { data_i[32:32] };
    end 
    if(N6888) begin
      { mem[511:511] } <= { data_i[31:31] };
    end 
    if(N6887) begin
      { mem[510:510] } <= { data_i[30:30] };
    end 
    if(N6886) begin
      { mem[509:509] } <= { data_i[29:29] };
    end 
    if(N6885) begin
      { mem[508:508] } <= { data_i[28:28] };
    end 
    if(N6884) begin
      { mem[507:507] } <= { data_i[27:27] };
    end 
    if(N6883) begin
      { mem[506:506] } <= { data_i[26:26] };
    end 
    if(N6882) begin
      { mem[505:505] } <= { data_i[25:25] };
    end 
    if(N6881) begin
      { mem[504:504] } <= { data_i[24:24] };
    end 
    if(N6880) begin
      { mem[503:503] } <= { data_i[23:23] };
    end 
    if(N6879) begin
      { mem[502:502] } <= { data_i[22:22] };
    end 
    if(N6878) begin
      { mem[501:501] } <= { data_i[21:21] };
    end 
    if(N6877) begin
      { mem[500:500] } <= { data_i[20:20] };
    end 
    if(N6876) begin
      { mem[499:499] } <= { data_i[19:19] };
    end 
    if(N6875) begin
      { mem[498:498] } <= { data_i[18:18] };
    end 
    if(N6874) begin
      { mem[497:497] } <= { data_i[17:17] };
    end 
    if(N6873) begin
      { mem[496:496] } <= { data_i[16:16] };
    end 
    if(N6872) begin
      { mem[495:495] } <= { data_i[15:15] };
    end 
    if(N6871) begin
      { mem[494:494] } <= { data_i[14:14] };
    end 
    if(N6870) begin
      { mem[493:493] } <= { data_i[13:13] };
    end 
    if(N6869) begin
      { mem[492:492] } <= { data_i[12:12] };
    end 
    if(N6868) begin
      { mem[491:491] } <= { data_i[11:11] };
    end 
    if(N6867) begin
      { mem[490:490] } <= { data_i[10:10] };
    end 
    if(N6866) begin
      { mem[489:489] } <= { data_i[9:9] };
    end 
    if(N6865) begin
      { mem[488:488] } <= { data_i[8:8] };
    end 
    if(N6864) begin
      { mem[487:487] } <= { data_i[7:7] };
    end 
    if(N6863) begin
      { mem[486:486] } <= { data_i[6:6] };
    end 
    if(N6862) begin
      { mem[485:485] } <= { data_i[5:5] };
    end 
    if(N6861) begin
      { mem[484:484] } <= { data_i[4:4] };
    end 
    if(N6860) begin
      { mem[483:483] } <= { data_i[3:3] };
    end 
    if(N6859) begin
      { mem[482:482] } <= { data_i[2:2] };
    end 
    if(N6858) begin
      { mem[481:481] } <= { data_i[1:1] };
    end 
    if(N6857) begin
      { mem[480:480] } <= { data_i[0:0] };
    end 
    if(N6856) begin
      { mem[479:479] } <= { data_i[79:79] };
    end 
    if(N6855) begin
      { mem[478:478] } <= { data_i[78:78] };
    end 
    if(N6854) begin
      { mem[477:477] } <= { data_i[77:77] };
    end 
    if(N6853) begin
      { mem[476:476] } <= { data_i[76:76] };
    end 
    if(N6852) begin
      { mem[475:475] } <= { data_i[75:75] };
    end 
    if(N6851) begin
      { mem[474:474] } <= { data_i[74:74] };
    end 
    if(N6850) begin
      { mem[473:473] } <= { data_i[73:73] };
    end 
    if(N6849) begin
      { mem[472:472] } <= { data_i[72:72] };
    end 
    if(N6848) begin
      { mem[471:471] } <= { data_i[71:71] };
    end 
    if(N6847) begin
      { mem[470:470] } <= { data_i[70:70] };
    end 
    if(N6846) begin
      { mem[469:469] } <= { data_i[69:69] };
    end 
    if(N6845) begin
      { mem[468:468] } <= { data_i[68:68] };
    end 
    if(N6844) begin
      { mem[467:467] } <= { data_i[67:67] };
    end 
    if(N6843) begin
      { mem[466:466] } <= { data_i[66:66] };
    end 
    if(N6842) begin
      { mem[465:465] } <= { data_i[65:65] };
    end 
    if(N6841) begin
      { mem[464:464] } <= { data_i[64:64] };
    end 
    if(N6840) begin
      { mem[463:463] } <= { data_i[63:63] };
    end 
    if(N6839) begin
      { mem[462:462] } <= { data_i[62:62] };
    end 
    if(N6838) begin
      { mem[461:461] } <= { data_i[61:61] };
    end 
    if(N6837) begin
      { mem[460:460] } <= { data_i[60:60] };
    end 
    if(N6836) begin
      { mem[459:459] } <= { data_i[59:59] };
    end 
    if(N6835) begin
      { mem[458:458] } <= { data_i[58:58] };
    end 
    if(N6834) begin
      { mem[457:457] } <= { data_i[57:57] };
    end 
    if(N6833) begin
      { mem[456:456] } <= { data_i[56:56] };
    end 
    if(N6832) begin
      { mem[455:455] } <= { data_i[55:55] };
    end 
    if(N6831) begin
      { mem[454:454] } <= { data_i[54:54] };
    end 
    if(N6830) begin
      { mem[453:453] } <= { data_i[53:53] };
    end 
    if(N6829) begin
      { mem[452:452] } <= { data_i[52:52] };
    end 
    if(N6828) begin
      { mem[451:451] } <= { data_i[51:51] };
    end 
    if(N6827) begin
      { mem[450:450] } <= { data_i[50:50] };
    end 
    if(N6826) begin
      { mem[449:449] } <= { data_i[49:49] };
    end 
    if(N6825) begin
      { mem[448:448] } <= { data_i[48:48] };
    end 
    if(N6824) begin
      { mem[447:447] } <= { data_i[47:47] };
    end 
    if(N6823) begin
      { mem[446:446] } <= { data_i[46:46] };
    end 
    if(N6822) begin
      { mem[445:445] } <= { data_i[45:45] };
    end 
    if(N6821) begin
      { mem[444:444] } <= { data_i[44:44] };
    end 
    if(N6820) begin
      { mem[443:443] } <= { data_i[43:43] };
    end 
    if(N6819) begin
      { mem[442:442] } <= { data_i[42:42] };
    end 
    if(N6818) begin
      { mem[441:441] } <= { data_i[41:41] };
    end 
    if(N6817) begin
      { mem[440:440] } <= { data_i[40:40] };
    end 
    if(N6816) begin
      { mem[439:439] } <= { data_i[39:39] };
    end 
    if(N6815) begin
      { mem[438:438] } <= { data_i[38:38] };
    end 
    if(N6814) begin
      { mem[437:437] } <= { data_i[37:37] };
    end 
    if(N6813) begin
      { mem[436:436] } <= { data_i[36:36] };
    end 
    if(N6812) begin
      { mem[435:435] } <= { data_i[35:35] };
    end 
    if(N6811) begin
      { mem[434:434] } <= { data_i[34:34] };
    end 
    if(N6810) begin
      { mem[433:433] } <= { data_i[33:33] };
    end 
    if(N6809) begin
      { mem[432:432] } <= { data_i[32:32] };
    end 
    if(N6808) begin
      { mem[431:431] } <= { data_i[31:31] };
    end 
    if(N6807) begin
      { mem[430:430] } <= { data_i[30:30] };
    end 
    if(N6806) begin
      { mem[429:429] } <= { data_i[29:29] };
    end 
    if(N6805) begin
      { mem[428:428] } <= { data_i[28:28] };
    end 
    if(N6804) begin
      { mem[427:427] } <= { data_i[27:27] };
    end 
    if(N6803) begin
      { mem[426:426] } <= { data_i[26:26] };
    end 
    if(N6802) begin
      { mem[425:425] } <= { data_i[25:25] };
    end 
    if(N6801) begin
      { mem[424:424] } <= { data_i[24:24] };
    end 
    if(N6800) begin
      { mem[423:423] } <= { data_i[23:23] };
    end 
    if(N6799) begin
      { mem[422:422] } <= { data_i[22:22] };
    end 
    if(N6798) begin
      { mem[421:421] } <= { data_i[21:21] };
    end 
    if(N6797) begin
      { mem[420:420] } <= { data_i[20:20] };
    end 
    if(N6796) begin
      { mem[419:419] } <= { data_i[19:19] };
    end 
    if(N6795) begin
      { mem[418:418] } <= { data_i[18:18] };
    end 
    if(N6794) begin
      { mem[417:417] } <= { data_i[17:17] };
    end 
    if(N6793) begin
      { mem[416:416] } <= { data_i[16:16] };
    end 
    if(N6792) begin
      { mem[415:415] } <= { data_i[15:15] };
    end 
    if(N6791) begin
      { mem[414:414] } <= { data_i[14:14] };
    end 
    if(N6790) begin
      { mem[413:413] } <= { data_i[13:13] };
    end 
    if(N6789) begin
      { mem[412:412] } <= { data_i[12:12] };
    end 
    if(N6788) begin
      { mem[411:411] } <= { data_i[11:11] };
    end 
    if(N6787) begin
      { mem[410:410] } <= { data_i[10:10] };
    end 
    if(N6786) begin
      { mem[409:409] } <= { data_i[9:9] };
    end 
    if(N6785) begin
      { mem[408:408] } <= { data_i[8:8] };
    end 
    if(N6784) begin
      { mem[407:407] } <= { data_i[7:7] };
    end 
    if(N6783) begin
      { mem[406:406] } <= { data_i[6:6] };
    end 
    if(N6782) begin
      { mem[405:405] } <= { data_i[5:5] };
    end 
    if(N6781) begin
      { mem[404:404] } <= { data_i[4:4] };
    end 
    if(N6780) begin
      { mem[403:403] } <= { data_i[3:3] };
    end 
    if(N6779) begin
      { mem[402:402] } <= { data_i[2:2] };
    end 
    if(N6778) begin
      { mem[401:401] } <= { data_i[1:1] };
    end 
    if(N6777) begin
      { mem[400:400] } <= { data_i[0:0] };
    end 
    if(N6776) begin
      { mem[399:399] } <= { data_i[79:79] };
    end 
    if(N6775) begin
      { mem[398:398] } <= { data_i[78:78] };
    end 
    if(N6774) begin
      { mem[397:397] } <= { data_i[77:77] };
    end 
    if(N6773) begin
      { mem[396:396] } <= { data_i[76:76] };
    end 
    if(N6772) begin
      { mem[395:395] } <= { data_i[75:75] };
    end 
    if(N6771) begin
      { mem[394:394] } <= { data_i[74:74] };
    end 
    if(N6770) begin
      { mem[393:393] } <= { data_i[73:73] };
    end 
    if(N6769) begin
      { mem[392:392] } <= { data_i[72:72] };
    end 
    if(N6768) begin
      { mem[391:391] } <= { data_i[71:71] };
    end 
    if(N6767) begin
      { mem[390:390] } <= { data_i[70:70] };
    end 
    if(N6766) begin
      { mem[389:389] } <= { data_i[69:69] };
    end 
    if(N6765) begin
      { mem[388:388] } <= { data_i[68:68] };
    end 
    if(N6764) begin
      { mem[387:387] } <= { data_i[67:67] };
    end 
    if(N6763) begin
      { mem[386:386] } <= { data_i[66:66] };
    end 
    if(N6762) begin
      { mem[385:385] } <= { data_i[65:65] };
    end 
    if(N6761) begin
      { mem[384:384] } <= { data_i[64:64] };
    end 
    if(N6760) begin
      { mem[383:383] } <= { data_i[63:63] };
    end 
    if(N6759) begin
      { mem[382:382] } <= { data_i[62:62] };
    end 
    if(N6758) begin
      { mem[381:381] } <= { data_i[61:61] };
    end 
    if(N6757) begin
      { mem[380:380] } <= { data_i[60:60] };
    end 
    if(N6756) begin
      { mem[379:379] } <= { data_i[59:59] };
    end 
    if(N6755) begin
      { mem[378:378] } <= { data_i[58:58] };
    end 
    if(N6754) begin
      { mem[377:377] } <= { data_i[57:57] };
    end 
    if(N6753) begin
      { mem[376:376] } <= { data_i[56:56] };
    end 
    if(N6752) begin
      { mem[375:375] } <= { data_i[55:55] };
    end 
    if(N6751) begin
      { mem[374:374] } <= { data_i[54:54] };
    end 
    if(N6750) begin
      { mem[373:373] } <= { data_i[53:53] };
    end 
    if(N6749) begin
      { mem[372:372] } <= { data_i[52:52] };
    end 
    if(N6748) begin
      { mem[371:371] } <= { data_i[51:51] };
    end 
    if(N6747) begin
      { mem[370:370] } <= { data_i[50:50] };
    end 
    if(N6746) begin
      { mem[369:369] } <= { data_i[49:49] };
    end 
    if(N6745) begin
      { mem[368:368] } <= { data_i[48:48] };
    end 
    if(N6744) begin
      { mem[367:367] } <= { data_i[47:47] };
    end 
    if(N6743) begin
      { mem[366:366] } <= { data_i[46:46] };
    end 
    if(N6742) begin
      { mem[365:365] } <= { data_i[45:45] };
    end 
    if(N6741) begin
      { mem[364:364] } <= { data_i[44:44] };
    end 
    if(N6740) begin
      { mem[363:363] } <= { data_i[43:43] };
    end 
    if(N6739) begin
      { mem[362:362] } <= { data_i[42:42] };
    end 
    if(N6738) begin
      { mem[361:361] } <= { data_i[41:41] };
    end 
    if(N6737) begin
      { mem[360:360] } <= { data_i[40:40] };
    end 
    if(N6736) begin
      { mem[359:359] } <= { data_i[39:39] };
    end 
    if(N6735) begin
      { mem[358:358] } <= { data_i[38:38] };
    end 
    if(N6734) begin
      { mem[357:357] } <= { data_i[37:37] };
    end 
    if(N6733) begin
      { mem[356:356] } <= { data_i[36:36] };
    end 
    if(N6732) begin
      { mem[355:355] } <= { data_i[35:35] };
    end 
    if(N6731) begin
      { mem[354:354] } <= { data_i[34:34] };
    end 
    if(N6730) begin
      { mem[353:353] } <= { data_i[33:33] };
    end 
    if(N6729) begin
      { mem[352:352] } <= { data_i[32:32] };
    end 
    if(N6728) begin
      { mem[351:351] } <= { data_i[31:31] };
    end 
    if(N6727) begin
      { mem[350:350] } <= { data_i[30:30] };
    end 
    if(N6726) begin
      { mem[349:349] } <= { data_i[29:29] };
    end 
    if(N6725) begin
      { mem[348:348] } <= { data_i[28:28] };
    end 
    if(N6724) begin
      { mem[347:347] } <= { data_i[27:27] };
    end 
    if(N6723) begin
      { mem[346:346] } <= { data_i[26:26] };
    end 
    if(N6722) begin
      { mem[345:345] } <= { data_i[25:25] };
    end 
    if(N6721) begin
      { mem[344:344] } <= { data_i[24:24] };
    end 
    if(N6720) begin
      { mem[343:343] } <= { data_i[23:23] };
    end 
    if(N6719) begin
      { mem[342:342] } <= { data_i[22:22] };
    end 
    if(N6718) begin
      { mem[341:341] } <= { data_i[21:21] };
    end 
    if(N6717) begin
      { mem[340:340] } <= { data_i[20:20] };
    end 
    if(N6716) begin
      { mem[339:339] } <= { data_i[19:19] };
    end 
    if(N6715) begin
      { mem[338:338] } <= { data_i[18:18] };
    end 
    if(N6714) begin
      { mem[337:337] } <= { data_i[17:17] };
    end 
    if(N6713) begin
      { mem[336:336] } <= { data_i[16:16] };
    end 
    if(N6712) begin
      { mem[335:335] } <= { data_i[15:15] };
    end 
    if(N6711) begin
      { mem[334:334] } <= { data_i[14:14] };
    end 
    if(N6710) begin
      { mem[333:333] } <= { data_i[13:13] };
    end 
    if(N6709) begin
      { mem[332:332] } <= { data_i[12:12] };
    end 
    if(N6708) begin
      { mem[331:331] } <= { data_i[11:11] };
    end 
    if(N6707) begin
      { mem[330:330] } <= { data_i[10:10] };
    end 
    if(N6706) begin
      { mem[329:329] } <= { data_i[9:9] };
    end 
    if(N6705) begin
      { mem[328:328] } <= { data_i[8:8] };
    end 
    if(N6704) begin
      { mem[327:327] } <= { data_i[7:7] };
    end 
    if(N6703) begin
      { mem[326:326] } <= { data_i[6:6] };
    end 
    if(N6702) begin
      { mem[325:325] } <= { data_i[5:5] };
    end 
    if(N6701) begin
      { mem[324:324] } <= { data_i[4:4] };
    end 
    if(N6700) begin
      { mem[323:323] } <= { data_i[3:3] };
    end 
    if(N6699) begin
      { mem[322:322] } <= { data_i[2:2] };
    end 
    if(N6698) begin
      { mem[321:321] } <= { data_i[1:1] };
    end 
    if(N6697) begin
      { mem[320:320] } <= { data_i[0:0] };
    end 
    if(N6696) begin
      { mem[319:319] } <= { data_i[79:79] };
    end 
    if(N6695) begin
      { mem[318:318] } <= { data_i[78:78] };
    end 
    if(N6694) begin
      { mem[317:317] } <= { data_i[77:77] };
    end 
    if(N6693) begin
      { mem[316:316] } <= { data_i[76:76] };
    end 
    if(N6692) begin
      { mem[315:315] } <= { data_i[75:75] };
    end 
    if(N6691) begin
      { mem[314:314] } <= { data_i[74:74] };
    end 
    if(N6690) begin
      { mem[313:313] } <= { data_i[73:73] };
    end 
    if(N6689) begin
      { mem[312:312] } <= { data_i[72:72] };
    end 
    if(N6688) begin
      { mem[311:311] } <= { data_i[71:71] };
    end 
    if(N6687) begin
      { mem[310:310] } <= { data_i[70:70] };
    end 
    if(N6686) begin
      { mem[309:309] } <= { data_i[69:69] };
    end 
    if(N6685) begin
      { mem[308:308] } <= { data_i[68:68] };
    end 
    if(N6684) begin
      { mem[307:307] } <= { data_i[67:67] };
    end 
    if(N6683) begin
      { mem[306:306] } <= { data_i[66:66] };
    end 
    if(N6682) begin
      { mem[305:305] } <= { data_i[65:65] };
    end 
    if(N6681) begin
      { mem[304:304] } <= { data_i[64:64] };
    end 
    if(N6680) begin
      { mem[303:303] } <= { data_i[63:63] };
    end 
    if(N6679) begin
      { mem[302:302] } <= { data_i[62:62] };
    end 
    if(N6678) begin
      { mem[301:301] } <= { data_i[61:61] };
    end 
    if(N6677) begin
      { mem[300:300] } <= { data_i[60:60] };
    end 
    if(N6676) begin
      { mem[299:299] } <= { data_i[59:59] };
    end 
    if(N6675) begin
      { mem[298:298] } <= { data_i[58:58] };
    end 
    if(N6674) begin
      { mem[297:297] } <= { data_i[57:57] };
    end 
    if(N6673) begin
      { mem[296:296] } <= { data_i[56:56] };
    end 
    if(N6672) begin
      { mem[295:295] } <= { data_i[55:55] };
    end 
    if(N6671) begin
      { mem[294:294] } <= { data_i[54:54] };
    end 
    if(N6670) begin
      { mem[293:293] } <= { data_i[53:53] };
    end 
    if(N6669) begin
      { mem[292:292] } <= { data_i[52:52] };
    end 
    if(N6668) begin
      { mem[291:291] } <= { data_i[51:51] };
    end 
    if(N6667) begin
      { mem[290:290] } <= { data_i[50:50] };
    end 
    if(N6666) begin
      { mem[289:289] } <= { data_i[49:49] };
    end 
    if(N6665) begin
      { mem[288:288] } <= { data_i[48:48] };
    end 
    if(N6664) begin
      { mem[287:287] } <= { data_i[47:47] };
    end 
    if(N6663) begin
      { mem[286:286] } <= { data_i[46:46] };
    end 
    if(N6662) begin
      { mem[285:285] } <= { data_i[45:45] };
    end 
    if(N6661) begin
      { mem[284:284] } <= { data_i[44:44] };
    end 
    if(N6660) begin
      { mem[283:283] } <= { data_i[43:43] };
    end 
    if(N6659) begin
      { mem[282:282] } <= { data_i[42:42] };
    end 
    if(N6658) begin
      { mem[281:281] } <= { data_i[41:41] };
    end 
    if(N6657) begin
      { mem[280:280] } <= { data_i[40:40] };
    end 
    if(N6656) begin
      { mem[279:279] } <= { data_i[39:39] };
    end 
    if(N6655) begin
      { mem[278:278] } <= { data_i[38:38] };
    end 
    if(N6654) begin
      { mem[277:277] } <= { data_i[37:37] };
    end 
    if(N6653) begin
      { mem[276:276] } <= { data_i[36:36] };
    end 
    if(N6652) begin
      { mem[275:275] } <= { data_i[35:35] };
    end 
    if(N6651) begin
      { mem[274:274] } <= { data_i[34:34] };
    end 
    if(N6650) begin
      { mem[273:273] } <= { data_i[33:33] };
    end 
    if(N6649) begin
      { mem[272:272] } <= { data_i[32:32] };
    end 
    if(N6648) begin
      { mem[271:271] } <= { data_i[31:31] };
    end 
    if(N6647) begin
      { mem[270:270] } <= { data_i[30:30] };
    end 
    if(N6646) begin
      { mem[269:269] } <= { data_i[29:29] };
    end 
    if(N6645) begin
      { mem[268:268] } <= { data_i[28:28] };
    end 
    if(N6644) begin
      { mem[267:267] } <= { data_i[27:27] };
    end 
    if(N6643) begin
      { mem[266:266] } <= { data_i[26:26] };
    end 
    if(N6642) begin
      { mem[265:265] } <= { data_i[25:25] };
    end 
    if(N6641) begin
      { mem[264:264] } <= { data_i[24:24] };
    end 
    if(N6640) begin
      { mem[263:263] } <= { data_i[23:23] };
    end 
    if(N6639) begin
      { mem[262:262] } <= { data_i[22:22] };
    end 
    if(N6638) begin
      { mem[261:261] } <= { data_i[21:21] };
    end 
    if(N6637) begin
      { mem[260:260] } <= { data_i[20:20] };
    end 
    if(N6636) begin
      { mem[259:259] } <= { data_i[19:19] };
    end 
    if(N6635) begin
      { mem[258:258] } <= { data_i[18:18] };
    end 
    if(N6634) begin
      { mem[257:257] } <= { data_i[17:17] };
    end 
    if(N6633) begin
      { mem[256:256] } <= { data_i[16:16] };
    end 
    if(N6632) begin
      { mem[255:255] } <= { data_i[15:15] };
    end 
    if(N6631) begin
      { mem[254:254] } <= { data_i[14:14] };
    end 
    if(N6630) begin
      { mem[253:253] } <= { data_i[13:13] };
    end 
    if(N6629) begin
      { mem[252:252] } <= { data_i[12:12] };
    end 
    if(N6628) begin
      { mem[251:251] } <= { data_i[11:11] };
    end 
    if(N6627) begin
      { mem[250:250] } <= { data_i[10:10] };
    end 
    if(N6626) begin
      { mem[249:249] } <= { data_i[9:9] };
    end 
    if(N6625) begin
      { mem[248:248] } <= { data_i[8:8] };
    end 
    if(N6624) begin
      { mem[247:247] } <= { data_i[7:7] };
    end 
    if(N6623) begin
      { mem[246:246] } <= { data_i[6:6] };
    end 
    if(N6622) begin
      { mem[245:245] } <= { data_i[5:5] };
    end 
    if(N6621) begin
      { mem[244:244] } <= { data_i[4:4] };
    end 
    if(N6620) begin
      { mem[243:243] } <= { data_i[3:3] };
    end 
    if(N6619) begin
      { mem[242:242] } <= { data_i[2:2] };
    end 
    if(N6618) begin
      { mem[241:241] } <= { data_i[1:1] };
    end 
    if(N6617) begin
      { mem[240:240] } <= { data_i[0:0] };
    end 
    if(N6616) begin
      { mem[239:239] } <= { data_i[79:79] };
    end 
    if(N6615) begin
      { mem[238:238] } <= { data_i[78:78] };
    end 
    if(N6614) begin
      { mem[237:237] } <= { data_i[77:77] };
    end 
    if(N6613) begin
      { mem[236:236] } <= { data_i[76:76] };
    end 
    if(N6612) begin
      { mem[235:235] } <= { data_i[75:75] };
    end 
    if(N6611) begin
      { mem[234:234] } <= { data_i[74:74] };
    end 
    if(N6610) begin
      { mem[233:233] } <= { data_i[73:73] };
    end 
    if(N6609) begin
      { mem[232:232] } <= { data_i[72:72] };
    end 
    if(N6608) begin
      { mem[231:231] } <= { data_i[71:71] };
    end 
    if(N6607) begin
      { mem[230:230] } <= { data_i[70:70] };
    end 
    if(N6606) begin
      { mem[229:229] } <= { data_i[69:69] };
    end 
    if(N6605) begin
      { mem[228:228] } <= { data_i[68:68] };
    end 
    if(N6604) begin
      { mem[227:227] } <= { data_i[67:67] };
    end 
    if(N6603) begin
      { mem[226:226] } <= { data_i[66:66] };
    end 
    if(N6602) begin
      { mem[225:225] } <= { data_i[65:65] };
    end 
    if(N6601) begin
      { mem[224:224] } <= { data_i[64:64] };
    end 
    if(N6600) begin
      { mem[223:223] } <= { data_i[63:63] };
    end 
    if(N6599) begin
      { mem[222:222] } <= { data_i[62:62] };
    end 
    if(N6598) begin
      { mem[221:221] } <= { data_i[61:61] };
    end 
    if(N6597) begin
      { mem[220:220] } <= { data_i[60:60] };
    end 
    if(N6596) begin
      { mem[219:219] } <= { data_i[59:59] };
    end 
    if(N6595) begin
      { mem[218:218] } <= { data_i[58:58] };
    end 
    if(N6594) begin
      { mem[217:217] } <= { data_i[57:57] };
    end 
    if(N6593) begin
      { mem[216:216] } <= { data_i[56:56] };
    end 
    if(N6592) begin
      { mem[215:215] } <= { data_i[55:55] };
    end 
    if(N6591) begin
      { mem[214:214] } <= { data_i[54:54] };
    end 
    if(N6590) begin
      { mem[213:213] } <= { data_i[53:53] };
    end 
    if(N6589) begin
      { mem[212:212] } <= { data_i[52:52] };
    end 
    if(N6588) begin
      { mem[211:211] } <= { data_i[51:51] };
    end 
    if(N6587) begin
      { mem[210:210] } <= { data_i[50:50] };
    end 
    if(N6586) begin
      { mem[209:209] } <= { data_i[49:49] };
    end 
    if(N6585) begin
      { mem[208:208] } <= { data_i[48:48] };
    end 
    if(N6584) begin
      { mem[207:207] } <= { data_i[47:47] };
    end 
    if(N6583) begin
      { mem[206:206] } <= { data_i[46:46] };
    end 
    if(N6582) begin
      { mem[205:205] } <= { data_i[45:45] };
    end 
    if(N6581) begin
      { mem[204:204] } <= { data_i[44:44] };
    end 
    if(N6580) begin
      { mem[203:203] } <= { data_i[43:43] };
    end 
    if(N6579) begin
      { mem[202:202] } <= { data_i[42:42] };
    end 
    if(N6578) begin
      { mem[201:201] } <= { data_i[41:41] };
    end 
    if(N6577) begin
      { mem[200:200] } <= { data_i[40:40] };
    end 
    if(N6576) begin
      { mem[199:199] } <= { data_i[39:39] };
    end 
    if(N6575) begin
      { mem[198:198] } <= { data_i[38:38] };
    end 
    if(N6574) begin
      { mem[197:197] } <= { data_i[37:37] };
    end 
    if(N6573) begin
      { mem[196:196] } <= { data_i[36:36] };
    end 
    if(N6572) begin
      { mem[195:195] } <= { data_i[35:35] };
    end 
    if(N6571) begin
      { mem[194:194] } <= { data_i[34:34] };
    end 
    if(N6570) begin
      { mem[193:193] } <= { data_i[33:33] };
    end 
    if(N6569) begin
      { mem[192:192] } <= { data_i[32:32] };
    end 
    if(N6568) begin
      { mem[191:191] } <= { data_i[31:31] };
    end 
    if(N6567) begin
      { mem[190:190] } <= { data_i[30:30] };
    end 
    if(N6566) begin
      { mem[189:189] } <= { data_i[29:29] };
    end 
    if(N6565) begin
      { mem[188:188] } <= { data_i[28:28] };
    end 
    if(N6564) begin
      { mem[187:187] } <= { data_i[27:27] };
    end 
    if(N6563) begin
      { mem[186:186] } <= { data_i[26:26] };
    end 
    if(N6562) begin
      { mem[185:185] } <= { data_i[25:25] };
    end 
    if(N6561) begin
      { mem[184:184] } <= { data_i[24:24] };
    end 
    if(N6560) begin
      { mem[183:183] } <= { data_i[23:23] };
    end 
    if(N6559) begin
      { mem[182:182] } <= { data_i[22:22] };
    end 
    if(N6558) begin
      { mem[181:181] } <= { data_i[21:21] };
    end 
    if(N6557) begin
      { mem[180:180] } <= { data_i[20:20] };
    end 
    if(N6556) begin
      { mem[179:179] } <= { data_i[19:19] };
    end 
    if(N6555) begin
      { mem[178:178] } <= { data_i[18:18] };
    end 
    if(N6554) begin
      { mem[177:177] } <= { data_i[17:17] };
    end 
    if(N6553) begin
      { mem[176:176] } <= { data_i[16:16] };
    end 
    if(N6552) begin
      { mem[175:175] } <= { data_i[15:15] };
    end 
    if(N6551) begin
      { mem[174:174] } <= { data_i[14:14] };
    end 
    if(N6550) begin
      { mem[173:173] } <= { data_i[13:13] };
    end 
    if(N6549) begin
      { mem[172:172] } <= { data_i[12:12] };
    end 
    if(N6548) begin
      { mem[171:171] } <= { data_i[11:11] };
    end 
    if(N6547) begin
      { mem[170:170] } <= { data_i[10:10] };
    end 
    if(N6546) begin
      { mem[169:169] } <= { data_i[9:9] };
    end 
    if(N6545) begin
      { mem[168:168] } <= { data_i[8:8] };
    end 
    if(N6544) begin
      { mem[167:167] } <= { data_i[7:7] };
    end 
    if(N6543) begin
      { mem[166:166] } <= { data_i[6:6] };
    end 
    if(N6542) begin
      { mem[165:165] } <= { data_i[5:5] };
    end 
    if(N6541) begin
      { mem[164:164] } <= { data_i[4:4] };
    end 
    if(N6540) begin
      { mem[163:163] } <= { data_i[3:3] };
    end 
    if(N6539) begin
      { mem[162:162] } <= { data_i[2:2] };
    end 
    if(N6538) begin
      { mem[161:161] } <= { data_i[1:1] };
    end 
    if(N6537) begin
      { mem[160:160] } <= { data_i[0:0] };
    end 
    if(N6536) begin
      { mem[159:159] } <= { data_i[79:79] };
    end 
    if(N6535) begin
      { mem[158:158] } <= { data_i[78:78] };
    end 
    if(N6534) begin
      { mem[157:157] } <= { data_i[77:77] };
    end 
    if(N6533) begin
      { mem[156:156] } <= { data_i[76:76] };
    end 
    if(N6532) begin
      { mem[155:155] } <= { data_i[75:75] };
    end 
    if(N6531) begin
      { mem[154:154] } <= { data_i[74:74] };
    end 
    if(N6530) begin
      { mem[153:153] } <= { data_i[73:73] };
    end 
    if(N6529) begin
      { mem[152:152] } <= { data_i[72:72] };
    end 
    if(N6528) begin
      { mem[151:151] } <= { data_i[71:71] };
    end 
    if(N6527) begin
      { mem[150:150] } <= { data_i[70:70] };
    end 
    if(N6526) begin
      { mem[149:149] } <= { data_i[69:69] };
    end 
    if(N6525) begin
      { mem[148:148] } <= { data_i[68:68] };
    end 
    if(N6524) begin
      { mem[147:147] } <= { data_i[67:67] };
    end 
    if(N6523) begin
      { mem[146:146] } <= { data_i[66:66] };
    end 
    if(N6522) begin
      { mem[145:145] } <= { data_i[65:65] };
    end 
    if(N6521) begin
      { mem[144:144] } <= { data_i[64:64] };
    end 
    if(N6520) begin
      { mem[143:143] } <= { data_i[63:63] };
    end 
    if(N6519) begin
      { mem[142:142] } <= { data_i[62:62] };
    end 
    if(N6518) begin
      { mem[141:141] } <= { data_i[61:61] };
    end 
    if(N6517) begin
      { mem[140:140] } <= { data_i[60:60] };
    end 
    if(N6516) begin
      { mem[139:139] } <= { data_i[59:59] };
    end 
    if(N6515) begin
      { mem[138:138] } <= { data_i[58:58] };
    end 
    if(N6514) begin
      { mem[137:137] } <= { data_i[57:57] };
    end 
    if(N6513) begin
      { mem[136:136] } <= { data_i[56:56] };
    end 
    if(N6512) begin
      { mem[135:135] } <= { data_i[55:55] };
    end 
    if(N6511) begin
      { mem[134:134] } <= { data_i[54:54] };
    end 
    if(N6510) begin
      { mem[133:133] } <= { data_i[53:53] };
    end 
    if(N6509) begin
      { mem[132:132] } <= { data_i[52:52] };
    end 
    if(N6508) begin
      { mem[131:131] } <= { data_i[51:51] };
    end 
    if(N6507) begin
      { mem[130:130] } <= { data_i[50:50] };
    end 
    if(N6506) begin
      { mem[129:129] } <= { data_i[49:49] };
    end 
    if(N6505) begin
      { mem[128:128] } <= { data_i[48:48] };
    end 
    if(N6504) begin
      { mem[127:127] } <= { data_i[47:47] };
    end 
    if(N6503) begin
      { mem[126:126] } <= { data_i[46:46] };
    end 
    if(N6502) begin
      { mem[125:125] } <= { data_i[45:45] };
    end 
    if(N6501) begin
      { mem[124:124] } <= { data_i[44:44] };
    end 
    if(N6500) begin
      { mem[123:123] } <= { data_i[43:43] };
    end 
    if(N6499) begin
      { mem[122:122] } <= { data_i[42:42] };
    end 
    if(N6498) begin
      { mem[121:121] } <= { data_i[41:41] };
    end 
    if(N6497) begin
      { mem[120:120] } <= { data_i[40:40] };
    end 
    if(N6496) begin
      { mem[119:119] } <= { data_i[39:39] };
    end 
    if(N6495) begin
      { mem[118:118] } <= { data_i[38:38] };
    end 
    if(N6494) begin
      { mem[117:117] } <= { data_i[37:37] };
    end 
    if(N6493) begin
      { mem[116:116] } <= { data_i[36:36] };
    end 
    if(N6492) begin
      { mem[115:115] } <= { data_i[35:35] };
    end 
    if(N6491) begin
      { mem[114:114] } <= { data_i[34:34] };
    end 
    if(N6490) begin
      { mem[113:113] } <= { data_i[33:33] };
    end 
    if(N6489) begin
      { mem[112:112] } <= { data_i[32:32] };
    end 
    if(N6488) begin
      { mem[111:111] } <= { data_i[31:31] };
    end 
    if(N6487) begin
      { mem[110:110] } <= { data_i[30:30] };
    end 
    if(N6486) begin
      { mem[109:109] } <= { data_i[29:29] };
    end 
    if(N6485) begin
      { mem[108:108] } <= { data_i[28:28] };
    end 
    if(N6484) begin
      { mem[107:107] } <= { data_i[27:27] };
    end 
    if(N6483) begin
      { mem[106:106] } <= { data_i[26:26] };
    end 
    if(N6482) begin
      { mem[105:105] } <= { data_i[25:25] };
    end 
    if(N6481) begin
      { mem[104:104] } <= { data_i[24:24] };
    end 
    if(N6480) begin
      { mem[103:103] } <= { data_i[23:23] };
    end 
    if(N6479) begin
      { mem[102:102] } <= { data_i[22:22] };
    end 
    if(N6478) begin
      { mem[101:101] } <= { data_i[21:21] };
    end 
    if(N6477) begin
      { mem[100:100] } <= { data_i[20:20] };
    end 
    if(N6476) begin
      { mem[99:99] } <= { data_i[19:19] };
    end 
    if(N6475) begin
      { mem[98:98] } <= { data_i[18:18] };
    end 
    if(N6474) begin
      { mem[97:97] } <= { data_i[17:17] };
    end 
    if(N6473) begin
      { mem[96:96] } <= { data_i[16:16] };
    end 
    if(N6472) begin
      { mem[95:95] } <= { data_i[15:15] };
    end 
    if(N6471) begin
      { mem[94:94] } <= { data_i[14:14] };
    end 
    if(N6470) begin
      { mem[93:93] } <= { data_i[13:13] };
    end 
    if(N6469) begin
      { mem[92:92] } <= { data_i[12:12] };
    end 
    if(N6468) begin
      { mem[91:91] } <= { data_i[11:11] };
    end 
    if(N6467) begin
      { mem[90:90] } <= { data_i[10:10] };
    end 
    if(N6466) begin
      { mem[89:89] } <= { data_i[9:9] };
    end 
    if(N6465) begin
      { mem[88:88] } <= { data_i[8:8] };
    end 
    if(N6464) begin
      { mem[87:87] } <= { data_i[7:7] };
    end 
    if(N6463) begin
      { mem[86:86] } <= { data_i[6:6] };
    end 
    if(N6462) begin
      { mem[85:85] } <= { data_i[5:5] };
    end 
    if(N6461) begin
      { mem[84:84] } <= { data_i[4:4] };
    end 
    if(N6460) begin
      { mem[83:83] } <= { data_i[3:3] };
    end 
    if(N6459) begin
      { mem[82:82] } <= { data_i[2:2] };
    end 
    if(N6458) begin
      { mem[81:81] } <= { data_i[1:1] };
    end 
    if(N6457) begin
      { mem[80:80] } <= { data_i[0:0] };
    end 
    if(N6456) begin
      { mem[79:79] } <= { data_i[79:79] };
    end 
    if(N6455) begin
      { mem[78:78] } <= { data_i[78:78] };
    end 
    if(N6454) begin
      { mem[77:77] } <= { data_i[77:77] };
    end 
    if(N6453) begin
      { mem[76:76] } <= { data_i[76:76] };
    end 
    if(N6452) begin
      { mem[75:75] } <= { data_i[75:75] };
    end 
    if(N6451) begin
      { mem[74:74] } <= { data_i[74:74] };
    end 
    if(N6450) begin
      { mem[73:73] } <= { data_i[73:73] };
    end 
    if(N6449) begin
      { mem[72:72] } <= { data_i[72:72] };
    end 
    if(N6448) begin
      { mem[71:71] } <= { data_i[71:71] };
    end 
    if(N6447) begin
      { mem[70:70] } <= { data_i[70:70] };
    end 
    if(N6446) begin
      { mem[69:69] } <= { data_i[69:69] };
    end 
    if(N6445) begin
      { mem[68:68] } <= { data_i[68:68] };
    end 
    if(N6444) begin
      { mem[67:67] } <= { data_i[67:67] };
    end 
    if(N6443) begin
      { mem[66:66] } <= { data_i[66:66] };
    end 
    if(N6442) begin
      { mem[65:65] } <= { data_i[65:65] };
    end 
    if(N6441) begin
      { mem[64:64] } <= { data_i[64:64] };
    end 
    if(N6440) begin
      { mem[63:63] } <= { data_i[63:63] };
    end 
    if(N6439) begin
      { mem[62:62] } <= { data_i[62:62] };
    end 
    if(N6438) begin
      { mem[61:61] } <= { data_i[61:61] };
    end 
    if(N6437) begin
      { mem[60:60] } <= { data_i[60:60] };
    end 
    if(N6436) begin
      { mem[59:59] } <= { data_i[59:59] };
    end 
    if(N6435) begin
      { mem[58:58] } <= { data_i[58:58] };
    end 
    if(N6434) begin
      { mem[57:57] } <= { data_i[57:57] };
    end 
    if(N6433) begin
      { mem[56:56] } <= { data_i[56:56] };
    end 
    if(N6432) begin
      { mem[55:55] } <= { data_i[55:55] };
    end 
    if(N6431) begin
      { mem[54:54] } <= { data_i[54:54] };
    end 
    if(N6430) begin
      { mem[53:53] } <= { data_i[53:53] };
    end 
    if(N6429) begin
      { mem[52:52] } <= { data_i[52:52] };
    end 
    if(N6428) begin
      { mem[51:51] } <= { data_i[51:51] };
    end 
    if(N6427) begin
      { mem[50:50] } <= { data_i[50:50] };
    end 
    if(N6426) begin
      { mem[49:49] } <= { data_i[49:49] };
    end 
    if(N6425) begin
      { mem[48:48] } <= { data_i[48:48] };
    end 
    if(N6424) begin
      { mem[47:47] } <= { data_i[47:47] };
    end 
    if(N6423) begin
      { mem[46:46] } <= { data_i[46:46] };
    end 
    if(N6422) begin
      { mem[45:45] } <= { data_i[45:45] };
    end 
    if(N6421) begin
      { mem[44:44] } <= { data_i[44:44] };
    end 
    if(N6420) begin
      { mem[43:43] } <= { data_i[43:43] };
    end 
    if(N6419) begin
      { mem[42:42] } <= { data_i[42:42] };
    end 
    if(N6418) begin
      { mem[41:41] } <= { data_i[41:41] };
    end 
    if(N6417) begin
      { mem[40:40] } <= { data_i[40:40] };
    end 
    if(N6416) begin
      { mem[39:39] } <= { data_i[39:39] };
    end 
    if(N6415) begin
      { mem[38:38] } <= { data_i[38:38] };
    end 
    if(N6414) begin
      { mem[37:37] } <= { data_i[37:37] };
    end 
    if(N6413) begin
      { mem[36:36] } <= { data_i[36:36] };
    end 
    if(N6412) begin
      { mem[35:35] } <= { data_i[35:35] };
    end 
    if(N6411) begin
      { mem[34:34] } <= { data_i[34:34] };
    end 
    if(N6410) begin
      { mem[33:33] } <= { data_i[33:33] };
    end 
    if(N6409) begin
      { mem[32:32] } <= { data_i[32:32] };
    end 
    if(N6408) begin
      { mem[31:31] } <= { data_i[31:31] };
    end 
    if(N6407) begin
      { mem[30:30] } <= { data_i[30:30] };
    end 
    if(N6406) begin
      { mem[29:29] } <= { data_i[29:29] };
    end 
    if(N6405) begin
      { mem[28:28] } <= { data_i[28:28] };
    end 
    if(N6404) begin
      { mem[27:27] } <= { data_i[27:27] };
    end 
    if(N6403) begin
      { mem[26:26] } <= { data_i[26:26] };
    end 
    if(N6402) begin
      { mem[25:25] } <= { data_i[25:25] };
    end 
    if(N6401) begin
      { mem[24:24] } <= { data_i[24:24] };
    end 
    if(N6400) begin
      { mem[23:23] } <= { data_i[23:23] };
    end 
    if(N6399) begin
      { mem[22:22] } <= { data_i[22:22] };
    end 
    if(N6398) begin
      { mem[21:21] } <= { data_i[21:21] };
    end 
    if(N6397) begin
      { mem[20:20] } <= { data_i[20:20] };
    end 
    if(N6396) begin
      { mem[19:19] } <= { data_i[19:19] };
    end 
    if(N6395) begin
      { mem[18:18] } <= { data_i[18:18] };
    end 
    if(N6394) begin
      { mem[17:17] } <= { data_i[17:17] };
    end 
    if(N6393) begin
      { mem[16:16] } <= { data_i[16:16] };
    end 
    if(N6392) begin
      { mem[15:15] } <= { data_i[15:15] };
    end 
    if(N6391) begin
      { mem[14:14] } <= { data_i[14:14] };
    end 
    if(N6390) begin
      { mem[13:13] } <= { data_i[13:13] };
    end 
    if(N6389) begin
      { mem[12:12] } <= { data_i[12:12] };
    end 
    if(N6388) begin
      { mem[11:11] } <= { data_i[11:11] };
    end 
    if(N6387) begin
      { mem[10:10] } <= { data_i[10:10] };
    end 
    if(N6386) begin
      { mem[9:9] } <= { data_i[9:9] };
    end 
    if(N6385) begin
      { mem[8:8] } <= { data_i[8:8] };
    end 
    if(N6384) begin
      { mem[7:7] } <= { data_i[7:7] };
    end 
    if(N6383) begin
      { mem[6:6] } <= { data_i[6:6] };
    end 
    if(N6382) begin
      { mem[5:5] } <= { data_i[5:5] };
    end 
    if(N6381) begin
      { mem[4:4] } <= { data_i[4:4] };
    end 
    if(N6380) begin
      { mem[3:3] } <= { data_i[3:3] };
    end 
    if(N6379) begin
      { mem[2:2] } <= { data_i[2:2] };
    end 
    if(N6378) begin
      { mem[1:1] } <= { data_i[1:1] };
    end 
    if(N6377) begin
      { mem[0:0] } <= { data_i[0:0] };
    end 
  end


endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p80_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [79:0] data_i;
  input [5:0] addr_i;
  input [79:0] w_mask_i;
  output [79:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [79:0] data_o;

  bsg_mem_1rw_sync_mask_write_bit_synth_width_p80_els_p64_latch_last_read_p1
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_dff_en_width_p8_harden_p0_strength_p0
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [7:0] data_i;
  output [7:0] data_o;
  input clk_i;
  input en_i;
  reg [7:0] data_o;

  always @(posedge clk_i) begin
    if(en_i) begin
      { data_o[7:0] } <= { data_i[7:0] };
    end 
  end


endmodule



module bsg_dff_en_bypass_width_p8
(
  clk_i,
  en_i,
  data_i,
  data_o
);

  input [7:0] data_i;
  output [7:0] data_o;
  input clk_i;
  input en_i;
  wire [7:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_en_width_p8_harden_p0_strength_p0
  dff
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .en_i(en_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_mem_1rw_sync_synth_width_p8_els_p256_latch_last_read_p1
(
  clk_i,
  v_i,
  reset_i,
  data_i,
  addr_i,
  w_i,
  data_o
);

  input [7:0] data_i;
  input [7:0] addr_i;
  output [7:0] data_o;
  input clk_i;
  input v_i;
  input reset_i;
  input w_i;
  wire [7:0] data_o,data_out;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,read_en,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
  N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,
  N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,
  N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,
  N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,
  N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,
  N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,
  N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,
  N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,
  N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,
  N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,
  N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,
  N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,
  N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,
  N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,
  N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,
  N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,
  N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,
  N532,llr_read_en_r,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,
  N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,
  N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,
  N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,
  N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,
  N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,
  N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,
  N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,
  N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,
  N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,
  N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,
  N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,
  N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,
  N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
  N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,
  N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,
  N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,
  N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,
  N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,
  N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,
  N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,
  N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,
  N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,
  N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,
  N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,
  N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,
  N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,
  N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,
  N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,
  N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,
  N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,
  N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,
  N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,
  N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,
  N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,
  N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,
  N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095;
  reg [7:0] addr_r;
  reg [2047:0] mem;
  assign data_out[7] = (N277)? mem[7] : 
                       (N279)? mem[15] : 
                       (N281)? mem[23] : 
                       (N283)? mem[31] : 
                       (N285)? mem[39] : 
                       (N287)? mem[47] : 
                       (N289)? mem[55] : 
                       (N291)? mem[63] : 
                       (N293)? mem[71] : 
                       (N295)? mem[79] : 
                       (N297)? mem[87] : 
                       (N299)? mem[95] : 
                       (N301)? mem[103] : 
                       (N303)? mem[111] : 
                       (N305)? mem[119] : 
                       (N307)? mem[127] : 
                       (N309)? mem[135] : 
                       (N311)? mem[143] : 
                       (N313)? mem[151] : 
                       (N315)? mem[159] : 
                       (N317)? mem[167] : 
                       (N319)? mem[175] : 
                       (N321)? mem[183] : 
                       (N323)? mem[191] : 
                       (N325)? mem[199] : 
                       (N327)? mem[207] : 
                       (N329)? mem[215] : 
                       (N331)? mem[223] : 
                       (N333)? mem[231] : 
                       (N335)? mem[239] : 
                       (N337)? mem[247] : 
                       (N339)? mem[255] : 
                       (N341)? mem[263] : 
                       (N343)? mem[271] : 
                       (N345)? mem[279] : 
                       (N347)? mem[287] : 
                       (N349)? mem[295] : 
                       (N351)? mem[303] : 
                       (N353)? mem[311] : 
                       (N355)? mem[319] : 
                       (N357)? mem[327] : 
                       (N359)? mem[335] : 
                       (N361)? mem[343] : 
                       (N363)? mem[351] : 
                       (N365)? mem[359] : 
                       (N367)? mem[367] : 
                       (N369)? mem[375] : 
                       (N371)? mem[383] : 
                       (N373)? mem[391] : 
                       (N375)? mem[399] : 
                       (N377)? mem[407] : 
                       (N379)? mem[415] : 
                       (N381)? mem[423] : 
                       (N383)? mem[431] : 
                       (N385)? mem[439] : 
                       (N387)? mem[447] : 
                       (N389)? mem[455] : 
                       (N391)? mem[463] : 
                       (N393)? mem[471] : 
                       (N395)? mem[479] : 
                       (N397)? mem[487] : 
                       (N399)? mem[495] : 
                       (N401)? mem[503] : 
                       (N403)? mem[511] : 
                       (N405)? mem[519] : 
                       (N407)? mem[527] : 
                       (N409)? mem[535] : 
                       (N411)? mem[543] : 
                       (N413)? mem[551] : 
                       (N415)? mem[559] : 
                       (N417)? mem[567] : 
                       (N419)? mem[575] : 
                       (N421)? mem[583] : 
                       (N423)? mem[591] : 
                       (N425)? mem[599] : 
                       (N427)? mem[607] : 
                       (N429)? mem[615] : 
                       (N431)? mem[623] : 
                       (N433)? mem[631] : 
                       (N435)? mem[639] : 
                       (N437)? mem[647] : 
                       (N439)? mem[655] : 
                       (N441)? mem[663] : 
                       (N443)? mem[671] : 
                       (N445)? mem[679] : 
                       (N447)? mem[687] : 
                       (N449)? mem[695] : 
                       (N451)? mem[703] : 
                       (N453)? mem[711] : 
                       (N455)? mem[719] : 
                       (N457)? mem[727] : 
                       (N459)? mem[735] : 
                       (N461)? mem[743] : 
                       (N463)? mem[751] : 
                       (N465)? mem[759] : 
                       (N467)? mem[767] : 
                       (N469)? mem[775] : 
                       (N471)? mem[783] : 
                       (N473)? mem[791] : 
                       (N475)? mem[799] : 
                       (N477)? mem[807] : 
                       (N479)? mem[815] : 
                       (N481)? mem[823] : 
                       (N483)? mem[831] : 
                       (N485)? mem[839] : 
                       (N487)? mem[847] : 
                       (N489)? mem[855] : 
                       (N491)? mem[863] : 
                       (N493)? mem[871] : 
                       (N495)? mem[879] : 
                       (N497)? mem[887] : 
                       (N499)? mem[895] : 
                       (N501)? mem[903] : 
                       (N503)? mem[911] : 
                       (N505)? mem[919] : 
                       (N507)? mem[927] : 
                       (N509)? mem[935] : 
                       (N511)? mem[943] : 
                       (N513)? mem[951] : 
                       (N515)? mem[959] : 
                       (N517)? mem[967] : 
                       (N519)? mem[975] : 
                       (N521)? mem[983] : 
                       (N523)? mem[991] : 
                       (N525)? mem[999] : 
                       (N527)? mem[1007] : 
                       (N529)? mem[1015] : 
                       (N531)? mem[1023] : 
                       (N278)? mem[1031] : 
                       (N280)? mem[1039] : 
                       (N282)? mem[1047] : 
                       (N284)? mem[1055] : 
                       (N286)? mem[1063] : 
                       (N288)? mem[1071] : 
                       (N290)? mem[1079] : 
                       (N292)? mem[1087] : 
                       (N294)? mem[1095] : 
                       (N296)? mem[1103] : 
                       (N298)? mem[1111] : 
                       (N300)? mem[1119] : 
                       (N302)? mem[1127] : 
                       (N304)? mem[1135] : 
                       (N306)? mem[1143] : 
                       (N308)? mem[1151] : 
                       (N310)? mem[1159] : 
                       (N312)? mem[1167] : 
                       (N314)? mem[1175] : 
                       (N316)? mem[1183] : 
                       (N318)? mem[1191] : 
                       (N320)? mem[1199] : 
                       (N322)? mem[1207] : 
                       (N324)? mem[1215] : 
                       (N326)? mem[1223] : 
                       (N328)? mem[1231] : 
                       (N330)? mem[1239] : 
                       (N332)? mem[1247] : 
                       (N334)? mem[1255] : 
                       (N336)? mem[1263] : 
                       (N338)? mem[1271] : 
                       (N340)? mem[1279] : 
                       (N342)? mem[1287] : 
                       (N344)? mem[1295] : 
                       (N346)? mem[1303] : 
                       (N348)? mem[1311] : 
                       (N350)? mem[1319] : 
                       (N352)? mem[1327] : 
                       (N354)? mem[1335] : 
                       (N356)? mem[1343] : 
                       (N358)? mem[1351] : 
                       (N360)? mem[1359] : 
                       (N362)? mem[1367] : 
                       (N364)? mem[1375] : 
                       (N366)? mem[1383] : 
                       (N368)? mem[1391] : 
                       (N370)? mem[1399] : 
                       (N372)? mem[1407] : 
                       (N374)? mem[1415] : 
                       (N376)? mem[1423] : 
                       (N378)? mem[1431] : 
                       (N380)? mem[1439] : 
                       (N382)? mem[1447] : 
                       (N384)? mem[1455] : 
                       (N386)? mem[1463] : 
                       (N388)? mem[1471] : 
                       (N390)? mem[1479] : 
                       (N392)? mem[1487] : 
                       (N394)? mem[1495] : 
                       (N396)? mem[1503] : 
                       (N398)? mem[1511] : 
                       (N400)? mem[1519] : 
                       (N402)? mem[1527] : 
                       (N404)? mem[1535] : 
                       (N406)? mem[1543] : 
                       (N408)? mem[1551] : 
                       (N410)? mem[1559] : 
                       (N412)? mem[1567] : 
                       (N414)? mem[1575] : 
                       (N416)? mem[1583] : 
                       (N418)? mem[1591] : 
                       (N420)? mem[1599] : 
                       (N422)? mem[1607] : 
                       (N424)? mem[1615] : 
                       (N426)? mem[1623] : 
                       (N428)? mem[1631] : 
                       (N430)? mem[1639] : 
                       (N432)? mem[1647] : 
                       (N434)? mem[1655] : 
                       (N436)? mem[1663] : 
                       (N438)? mem[1671] : 
                       (N440)? mem[1679] : 
                       (N442)? mem[1687] : 
                       (N444)? mem[1695] : 
                       (N446)? mem[1703] : 
                       (N448)? mem[1711] : 
                       (N450)? mem[1719] : 
                       (N452)? mem[1727] : 
                       (N454)? mem[1735] : 
                       (N456)? mem[1743] : 
                       (N458)? mem[1751] : 
                       (N460)? mem[1759] : 
                       (N462)? mem[1767] : 
                       (N464)? mem[1775] : 
                       (N466)? mem[1783] : 
                       (N468)? mem[1791] : 
                       (N470)? mem[1799] : 
                       (N472)? mem[1807] : 
                       (N474)? mem[1815] : 
                       (N476)? mem[1823] : 
                       (N478)? mem[1831] : 
                       (N480)? mem[1839] : 
                       (N482)? mem[1847] : 
                       (N484)? mem[1855] : 
                       (N486)? mem[1863] : 
                       (N488)? mem[1871] : 
                       (N490)? mem[1879] : 
                       (N492)? mem[1887] : 
                       (N494)? mem[1895] : 
                       (N496)? mem[1903] : 
                       (N498)? mem[1911] : 
                       (N500)? mem[1919] : 
                       (N502)? mem[1927] : 
                       (N504)? mem[1935] : 
                       (N506)? mem[1943] : 
                       (N508)? mem[1951] : 
                       (N510)? mem[1959] : 
                       (N512)? mem[1967] : 
                       (N514)? mem[1975] : 
                       (N516)? mem[1983] : 
                       (N518)? mem[1991] : 
                       (N520)? mem[1999] : 
                       (N522)? mem[2007] : 
                       (N524)? mem[2015] : 
                       (N526)? mem[2023] : 
                       (N528)? mem[2031] : 
                       (N530)? mem[2039] : 
                       (N532)? mem[2047] : 1'b0;
  assign data_out[6] = (N277)? mem[6] : 
                       (N279)? mem[14] : 
                       (N281)? mem[22] : 
                       (N283)? mem[30] : 
                       (N285)? mem[38] : 
                       (N287)? mem[46] : 
                       (N289)? mem[54] : 
                       (N291)? mem[62] : 
                       (N293)? mem[70] : 
                       (N295)? mem[78] : 
                       (N297)? mem[86] : 
                       (N299)? mem[94] : 
                       (N301)? mem[102] : 
                       (N303)? mem[110] : 
                       (N305)? mem[118] : 
                       (N307)? mem[126] : 
                       (N309)? mem[134] : 
                       (N311)? mem[142] : 
                       (N313)? mem[150] : 
                       (N315)? mem[158] : 
                       (N317)? mem[166] : 
                       (N319)? mem[174] : 
                       (N321)? mem[182] : 
                       (N323)? mem[190] : 
                       (N325)? mem[198] : 
                       (N327)? mem[206] : 
                       (N329)? mem[214] : 
                       (N331)? mem[222] : 
                       (N333)? mem[230] : 
                       (N335)? mem[238] : 
                       (N337)? mem[246] : 
                       (N339)? mem[254] : 
                       (N341)? mem[262] : 
                       (N343)? mem[270] : 
                       (N345)? mem[278] : 
                       (N347)? mem[286] : 
                       (N349)? mem[294] : 
                       (N351)? mem[302] : 
                       (N353)? mem[310] : 
                       (N355)? mem[318] : 
                       (N357)? mem[326] : 
                       (N359)? mem[334] : 
                       (N361)? mem[342] : 
                       (N363)? mem[350] : 
                       (N365)? mem[358] : 
                       (N367)? mem[366] : 
                       (N369)? mem[374] : 
                       (N371)? mem[382] : 
                       (N373)? mem[390] : 
                       (N375)? mem[398] : 
                       (N377)? mem[406] : 
                       (N379)? mem[414] : 
                       (N381)? mem[422] : 
                       (N383)? mem[430] : 
                       (N385)? mem[438] : 
                       (N387)? mem[446] : 
                       (N389)? mem[454] : 
                       (N391)? mem[462] : 
                       (N393)? mem[470] : 
                       (N395)? mem[478] : 
                       (N397)? mem[486] : 
                       (N399)? mem[494] : 
                       (N401)? mem[502] : 
                       (N403)? mem[510] : 
                       (N405)? mem[518] : 
                       (N407)? mem[526] : 
                       (N409)? mem[534] : 
                       (N411)? mem[542] : 
                       (N413)? mem[550] : 
                       (N415)? mem[558] : 
                       (N417)? mem[566] : 
                       (N419)? mem[574] : 
                       (N421)? mem[582] : 
                       (N423)? mem[590] : 
                       (N425)? mem[598] : 
                       (N427)? mem[606] : 
                       (N429)? mem[614] : 
                       (N431)? mem[622] : 
                       (N433)? mem[630] : 
                       (N435)? mem[638] : 
                       (N437)? mem[646] : 
                       (N439)? mem[654] : 
                       (N441)? mem[662] : 
                       (N443)? mem[670] : 
                       (N445)? mem[678] : 
                       (N447)? mem[686] : 
                       (N449)? mem[694] : 
                       (N451)? mem[702] : 
                       (N453)? mem[710] : 
                       (N455)? mem[718] : 
                       (N457)? mem[726] : 
                       (N459)? mem[734] : 
                       (N461)? mem[742] : 
                       (N463)? mem[750] : 
                       (N465)? mem[758] : 
                       (N467)? mem[766] : 
                       (N469)? mem[774] : 
                       (N471)? mem[782] : 
                       (N473)? mem[790] : 
                       (N475)? mem[798] : 
                       (N477)? mem[806] : 
                       (N479)? mem[814] : 
                       (N481)? mem[822] : 
                       (N483)? mem[830] : 
                       (N485)? mem[838] : 
                       (N487)? mem[846] : 
                       (N489)? mem[854] : 
                       (N491)? mem[862] : 
                       (N493)? mem[870] : 
                       (N495)? mem[878] : 
                       (N497)? mem[886] : 
                       (N499)? mem[894] : 
                       (N501)? mem[902] : 
                       (N503)? mem[910] : 
                       (N505)? mem[918] : 
                       (N507)? mem[926] : 
                       (N509)? mem[934] : 
                       (N511)? mem[942] : 
                       (N513)? mem[950] : 
                       (N515)? mem[958] : 
                       (N517)? mem[966] : 
                       (N519)? mem[974] : 
                       (N521)? mem[982] : 
                       (N523)? mem[990] : 
                       (N525)? mem[998] : 
                       (N527)? mem[1006] : 
                       (N529)? mem[1014] : 
                       (N531)? mem[1022] : 
                       (N278)? mem[1030] : 
                       (N280)? mem[1038] : 
                       (N282)? mem[1046] : 
                       (N284)? mem[1054] : 
                       (N286)? mem[1062] : 
                       (N288)? mem[1070] : 
                       (N290)? mem[1078] : 
                       (N292)? mem[1086] : 
                       (N294)? mem[1094] : 
                       (N296)? mem[1102] : 
                       (N298)? mem[1110] : 
                       (N300)? mem[1118] : 
                       (N302)? mem[1126] : 
                       (N304)? mem[1134] : 
                       (N306)? mem[1142] : 
                       (N308)? mem[1150] : 
                       (N310)? mem[1158] : 
                       (N312)? mem[1166] : 
                       (N314)? mem[1174] : 
                       (N316)? mem[1182] : 
                       (N318)? mem[1190] : 
                       (N320)? mem[1198] : 
                       (N322)? mem[1206] : 
                       (N324)? mem[1214] : 
                       (N326)? mem[1222] : 
                       (N328)? mem[1230] : 
                       (N330)? mem[1238] : 
                       (N332)? mem[1246] : 
                       (N334)? mem[1254] : 
                       (N336)? mem[1262] : 
                       (N338)? mem[1270] : 
                       (N340)? mem[1278] : 
                       (N342)? mem[1286] : 
                       (N344)? mem[1294] : 
                       (N346)? mem[1302] : 
                       (N348)? mem[1310] : 
                       (N350)? mem[1318] : 
                       (N352)? mem[1326] : 
                       (N354)? mem[1334] : 
                       (N356)? mem[1342] : 
                       (N358)? mem[1350] : 
                       (N360)? mem[1358] : 
                       (N362)? mem[1366] : 
                       (N364)? mem[1374] : 
                       (N366)? mem[1382] : 
                       (N368)? mem[1390] : 
                       (N370)? mem[1398] : 
                       (N372)? mem[1406] : 
                       (N374)? mem[1414] : 
                       (N376)? mem[1422] : 
                       (N378)? mem[1430] : 
                       (N380)? mem[1438] : 
                       (N382)? mem[1446] : 
                       (N384)? mem[1454] : 
                       (N386)? mem[1462] : 
                       (N388)? mem[1470] : 
                       (N390)? mem[1478] : 
                       (N392)? mem[1486] : 
                       (N394)? mem[1494] : 
                       (N396)? mem[1502] : 
                       (N398)? mem[1510] : 
                       (N400)? mem[1518] : 
                       (N402)? mem[1526] : 
                       (N404)? mem[1534] : 
                       (N406)? mem[1542] : 
                       (N408)? mem[1550] : 
                       (N410)? mem[1558] : 
                       (N412)? mem[1566] : 
                       (N414)? mem[1574] : 
                       (N416)? mem[1582] : 
                       (N418)? mem[1590] : 
                       (N420)? mem[1598] : 
                       (N422)? mem[1606] : 
                       (N424)? mem[1614] : 
                       (N426)? mem[1622] : 
                       (N428)? mem[1630] : 
                       (N430)? mem[1638] : 
                       (N432)? mem[1646] : 
                       (N434)? mem[1654] : 
                       (N436)? mem[1662] : 
                       (N438)? mem[1670] : 
                       (N440)? mem[1678] : 
                       (N442)? mem[1686] : 
                       (N444)? mem[1694] : 
                       (N446)? mem[1702] : 
                       (N448)? mem[1710] : 
                       (N450)? mem[1718] : 
                       (N452)? mem[1726] : 
                       (N454)? mem[1734] : 
                       (N456)? mem[1742] : 
                       (N458)? mem[1750] : 
                       (N460)? mem[1758] : 
                       (N462)? mem[1766] : 
                       (N464)? mem[1774] : 
                       (N466)? mem[1782] : 
                       (N468)? mem[1790] : 
                       (N470)? mem[1798] : 
                       (N472)? mem[1806] : 
                       (N474)? mem[1814] : 
                       (N476)? mem[1822] : 
                       (N478)? mem[1830] : 
                       (N480)? mem[1838] : 
                       (N482)? mem[1846] : 
                       (N484)? mem[1854] : 
                       (N486)? mem[1862] : 
                       (N488)? mem[1870] : 
                       (N490)? mem[1878] : 
                       (N492)? mem[1886] : 
                       (N494)? mem[1894] : 
                       (N496)? mem[1902] : 
                       (N498)? mem[1910] : 
                       (N500)? mem[1918] : 
                       (N502)? mem[1926] : 
                       (N504)? mem[1934] : 
                       (N506)? mem[1942] : 
                       (N508)? mem[1950] : 
                       (N510)? mem[1958] : 
                       (N512)? mem[1966] : 
                       (N514)? mem[1974] : 
                       (N516)? mem[1982] : 
                       (N518)? mem[1990] : 
                       (N520)? mem[1998] : 
                       (N522)? mem[2006] : 
                       (N524)? mem[2014] : 
                       (N526)? mem[2022] : 
                       (N528)? mem[2030] : 
                       (N530)? mem[2038] : 
                       (N532)? mem[2046] : 1'b0;
  assign data_out[5] = (N277)? mem[5] : 
                       (N279)? mem[13] : 
                       (N281)? mem[21] : 
                       (N283)? mem[29] : 
                       (N285)? mem[37] : 
                       (N287)? mem[45] : 
                       (N289)? mem[53] : 
                       (N291)? mem[61] : 
                       (N293)? mem[69] : 
                       (N295)? mem[77] : 
                       (N297)? mem[85] : 
                       (N299)? mem[93] : 
                       (N301)? mem[101] : 
                       (N303)? mem[109] : 
                       (N305)? mem[117] : 
                       (N307)? mem[125] : 
                       (N309)? mem[133] : 
                       (N311)? mem[141] : 
                       (N313)? mem[149] : 
                       (N315)? mem[157] : 
                       (N317)? mem[165] : 
                       (N319)? mem[173] : 
                       (N321)? mem[181] : 
                       (N323)? mem[189] : 
                       (N325)? mem[197] : 
                       (N327)? mem[205] : 
                       (N329)? mem[213] : 
                       (N331)? mem[221] : 
                       (N333)? mem[229] : 
                       (N335)? mem[237] : 
                       (N337)? mem[245] : 
                       (N339)? mem[253] : 
                       (N341)? mem[261] : 
                       (N343)? mem[269] : 
                       (N345)? mem[277] : 
                       (N347)? mem[285] : 
                       (N349)? mem[293] : 
                       (N351)? mem[301] : 
                       (N353)? mem[309] : 
                       (N355)? mem[317] : 
                       (N357)? mem[325] : 
                       (N359)? mem[333] : 
                       (N361)? mem[341] : 
                       (N363)? mem[349] : 
                       (N365)? mem[357] : 
                       (N367)? mem[365] : 
                       (N369)? mem[373] : 
                       (N371)? mem[381] : 
                       (N373)? mem[389] : 
                       (N375)? mem[397] : 
                       (N377)? mem[405] : 
                       (N379)? mem[413] : 
                       (N381)? mem[421] : 
                       (N383)? mem[429] : 
                       (N385)? mem[437] : 
                       (N387)? mem[445] : 
                       (N389)? mem[453] : 
                       (N391)? mem[461] : 
                       (N393)? mem[469] : 
                       (N395)? mem[477] : 
                       (N397)? mem[485] : 
                       (N399)? mem[493] : 
                       (N401)? mem[501] : 
                       (N403)? mem[509] : 
                       (N405)? mem[517] : 
                       (N407)? mem[525] : 
                       (N409)? mem[533] : 
                       (N411)? mem[541] : 
                       (N413)? mem[549] : 
                       (N415)? mem[557] : 
                       (N417)? mem[565] : 
                       (N419)? mem[573] : 
                       (N421)? mem[581] : 
                       (N423)? mem[589] : 
                       (N425)? mem[597] : 
                       (N427)? mem[605] : 
                       (N429)? mem[613] : 
                       (N431)? mem[621] : 
                       (N433)? mem[629] : 
                       (N435)? mem[637] : 
                       (N437)? mem[645] : 
                       (N439)? mem[653] : 
                       (N441)? mem[661] : 
                       (N443)? mem[669] : 
                       (N445)? mem[677] : 
                       (N447)? mem[685] : 
                       (N449)? mem[693] : 
                       (N451)? mem[701] : 
                       (N453)? mem[709] : 
                       (N455)? mem[717] : 
                       (N457)? mem[725] : 
                       (N459)? mem[733] : 
                       (N461)? mem[741] : 
                       (N463)? mem[749] : 
                       (N465)? mem[757] : 
                       (N467)? mem[765] : 
                       (N469)? mem[773] : 
                       (N471)? mem[781] : 
                       (N473)? mem[789] : 
                       (N475)? mem[797] : 
                       (N477)? mem[805] : 
                       (N479)? mem[813] : 
                       (N481)? mem[821] : 
                       (N483)? mem[829] : 
                       (N485)? mem[837] : 
                       (N487)? mem[845] : 
                       (N489)? mem[853] : 
                       (N491)? mem[861] : 
                       (N493)? mem[869] : 
                       (N495)? mem[877] : 
                       (N497)? mem[885] : 
                       (N499)? mem[893] : 
                       (N501)? mem[901] : 
                       (N503)? mem[909] : 
                       (N505)? mem[917] : 
                       (N507)? mem[925] : 
                       (N509)? mem[933] : 
                       (N511)? mem[941] : 
                       (N513)? mem[949] : 
                       (N515)? mem[957] : 
                       (N517)? mem[965] : 
                       (N519)? mem[973] : 
                       (N521)? mem[981] : 
                       (N523)? mem[989] : 
                       (N525)? mem[997] : 
                       (N527)? mem[1005] : 
                       (N529)? mem[1013] : 
                       (N531)? mem[1021] : 
                       (N278)? mem[1029] : 
                       (N280)? mem[1037] : 
                       (N282)? mem[1045] : 
                       (N284)? mem[1053] : 
                       (N286)? mem[1061] : 
                       (N288)? mem[1069] : 
                       (N290)? mem[1077] : 
                       (N292)? mem[1085] : 
                       (N294)? mem[1093] : 
                       (N296)? mem[1101] : 
                       (N298)? mem[1109] : 
                       (N300)? mem[1117] : 
                       (N302)? mem[1125] : 
                       (N304)? mem[1133] : 
                       (N306)? mem[1141] : 
                       (N308)? mem[1149] : 
                       (N310)? mem[1157] : 
                       (N312)? mem[1165] : 
                       (N314)? mem[1173] : 
                       (N316)? mem[1181] : 
                       (N318)? mem[1189] : 
                       (N320)? mem[1197] : 
                       (N322)? mem[1205] : 
                       (N324)? mem[1213] : 
                       (N326)? mem[1221] : 
                       (N328)? mem[1229] : 
                       (N330)? mem[1237] : 
                       (N332)? mem[1245] : 
                       (N334)? mem[1253] : 
                       (N336)? mem[1261] : 
                       (N338)? mem[1269] : 
                       (N340)? mem[1277] : 
                       (N342)? mem[1285] : 
                       (N344)? mem[1293] : 
                       (N346)? mem[1301] : 
                       (N348)? mem[1309] : 
                       (N350)? mem[1317] : 
                       (N352)? mem[1325] : 
                       (N354)? mem[1333] : 
                       (N356)? mem[1341] : 
                       (N358)? mem[1349] : 
                       (N360)? mem[1357] : 
                       (N362)? mem[1365] : 
                       (N364)? mem[1373] : 
                       (N366)? mem[1381] : 
                       (N368)? mem[1389] : 
                       (N370)? mem[1397] : 
                       (N372)? mem[1405] : 
                       (N374)? mem[1413] : 
                       (N376)? mem[1421] : 
                       (N378)? mem[1429] : 
                       (N380)? mem[1437] : 
                       (N382)? mem[1445] : 
                       (N384)? mem[1453] : 
                       (N386)? mem[1461] : 
                       (N388)? mem[1469] : 
                       (N390)? mem[1477] : 
                       (N392)? mem[1485] : 
                       (N394)? mem[1493] : 
                       (N396)? mem[1501] : 
                       (N398)? mem[1509] : 
                       (N400)? mem[1517] : 
                       (N402)? mem[1525] : 
                       (N404)? mem[1533] : 
                       (N406)? mem[1541] : 
                       (N408)? mem[1549] : 
                       (N410)? mem[1557] : 
                       (N412)? mem[1565] : 
                       (N414)? mem[1573] : 
                       (N416)? mem[1581] : 
                       (N418)? mem[1589] : 
                       (N420)? mem[1597] : 
                       (N422)? mem[1605] : 
                       (N424)? mem[1613] : 
                       (N426)? mem[1621] : 
                       (N428)? mem[1629] : 
                       (N430)? mem[1637] : 
                       (N432)? mem[1645] : 
                       (N434)? mem[1653] : 
                       (N436)? mem[1661] : 
                       (N438)? mem[1669] : 
                       (N440)? mem[1677] : 
                       (N442)? mem[1685] : 
                       (N444)? mem[1693] : 
                       (N446)? mem[1701] : 
                       (N448)? mem[1709] : 
                       (N450)? mem[1717] : 
                       (N452)? mem[1725] : 
                       (N454)? mem[1733] : 
                       (N456)? mem[1741] : 
                       (N458)? mem[1749] : 
                       (N460)? mem[1757] : 
                       (N462)? mem[1765] : 
                       (N464)? mem[1773] : 
                       (N466)? mem[1781] : 
                       (N468)? mem[1789] : 
                       (N470)? mem[1797] : 
                       (N472)? mem[1805] : 
                       (N474)? mem[1813] : 
                       (N476)? mem[1821] : 
                       (N478)? mem[1829] : 
                       (N480)? mem[1837] : 
                       (N482)? mem[1845] : 
                       (N484)? mem[1853] : 
                       (N486)? mem[1861] : 
                       (N488)? mem[1869] : 
                       (N490)? mem[1877] : 
                       (N492)? mem[1885] : 
                       (N494)? mem[1893] : 
                       (N496)? mem[1901] : 
                       (N498)? mem[1909] : 
                       (N500)? mem[1917] : 
                       (N502)? mem[1925] : 
                       (N504)? mem[1933] : 
                       (N506)? mem[1941] : 
                       (N508)? mem[1949] : 
                       (N510)? mem[1957] : 
                       (N512)? mem[1965] : 
                       (N514)? mem[1973] : 
                       (N516)? mem[1981] : 
                       (N518)? mem[1989] : 
                       (N520)? mem[1997] : 
                       (N522)? mem[2005] : 
                       (N524)? mem[2013] : 
                       (N526)? mem[2021] : 
                       (N528)? mem[2029] : 
                       (N530)? mem[2037] : 
                       (N532)? mem[2045] : 1'b0;
  assign data_out[4] = (N277)? mem[4] : 
                       (N279)? mem[12] : 
                       (N281)? mem[20] : 
                       (N283)? mem[28] : 
                       (N285)? mem[36] : 
                       (N287)? mem[44] : 
                       (N289)? mem[52] : 
                       (N291)? mem[60] : 
                       (N293)? mem[68] : 
                       (N295)? mem[76] : 
                       (N297)? mem[84] : 
                       (N299)? mem[92] : 
                       (N301)? mem[100] : 
                       (N303)? mem[108] : 
                       (N305)? mem[116] : 
                       (N307)? mem[124] : 
                       (N309)? mem[132] : 
                       (N311)? mem[140] : 
                       (N313)? mem[148] : 
                       (N315)? mem[156] : 
                       (N317)? mem[164] : 
                       (N319)? mem[172] : 
                       (N321)? mem[180] : 
                       (N323)? mem[188] : 
                       (N325)? mem[196] : 
                       (N327)? mem[204] : 
                       (N329)? mem[212] : 
                       (N331)? mem[220] : 
                       (N333)? mem[228] : 
                       (N335)? mem[236] : 
                       (N337)? mem[244] : 
                       (N339)? mem[252] : 
                       (N341)? mem[260] : 
                       (N343)? mem[268] : 
                       (N345)? mem[276] : 
                       (N347)? mem[284] : 
                       (N349)? mem[292] : 
                       (N351)? mem[300] : 
                       (N353)? mem[308] : 
                       (N355)? mem[316] : 
                       (N357)? mem[324] : 
                       (N359)? mem[332] : 
                       (N361)? mem[340] : 
                       (N363)? mem[348] : 
                       (N365)? mem[356] : 
                       (N367)? mem[364] : 
                       (N369)? mem[372] : 
                       (N371)? mem[380] : 
                       (N373)? mem[388] : 
                       (N375)? mem[396] : 
                       (N377)? mem[404] : 
                       (N379)? mem[412] : 
                       (N381)? mem[420] : 
                       (N383)? mem[428] : 
                       (N385)? mem[436] : 
                       (N387)? mem[444] : 
                       (N389)? mem[452] : 
                       (N391)? mem[460] : 
                       (N393)? mem[468] : 
                       (N395)? mem[476] : 
                       (N397)? mem[484] : 
                       (N399)? mem[492] : 
                       (N401)? mem[500] : 
                       (N403)? mem[508] : 
                       (N405)? mem[516] : 
                       (N407)? mem[524] : 
                       (N409)? mem[532] : 
                       (N411)? mem[540] : 
                       (N413)? mem[548] : 
                       (N415)? mem[556] : 
                       (N417)? mem[564] : 
                       (N419)? mem[572] : 
                       (N421)? mem[580] : 
                       (N423)? mem[588] : 
                       (N425)? mem[596] : 
                       (N427)? mem[604] : 
                       (N429)? mem[612] : 
                       (N431)? mem[620] : 
                       (N433)? mem[628] : 
                       (N435)? mem[636] : 
                       (N437)? mem[644] : 
                       (N439)? mem[652] : 
                       (N441)? mem[660] : 
                       (N443)? mem[668] : 
                       (N445)? mem[676] : 
                       (N447)? mem[684] : 
                       (N449)? mem[692] : 
                       (N451)? mem[700] : 
                       (N453)? mem[708] : 
                       (N455)? mem[716] : 
                       (N457)? mem[724] : 
                       (N459)? mem[732] : 
                       (N461)? mem[740] : 
                       (N463)? mem[748] : 
                       (N465)? mem[756] : 
                       (N467)? mem[764] : 
                       (N469)? mem[772] : 
                       (N471)? mem[780] : 
                       (N473)? mem[788] : 
                       (N475)? mem[796] : 
                       (N477)? mem[804] : 
                       (N479)? mem[812] : 
                       (N481)? mem[820] : 
                       (N483)? mem[828] : 
                       (N485)? mem[836] : 
                       (N487)? mem[844] : 
                       (N489)? mem[852] : 
                       (N491)? mem[860] : 
                       (N493)? mem[868] : 
                       (N495)? mem[876] : 
                       (N497)? mem[884] : 
                       (N499)? mem[892] : 
                       (N501)? mem[900] : 
                       (N503)? mem[908] : 
                       (N505)? mem[916] : 
                       (N507)? mem[924] : 
                       (N509)? mem[932] : 
                       (N511)? mem[940] : 
                       (N513)? mem[948] : 
                       (N515)? mem[956] : 
                       (N517)? mem[964] : 
                       (N519)? mem[972] : 
                       (N521)? mem[980] : 
                       (N523)? mem[988] : 
                       (N525)? mem[996] : 
                       (N527)? mem[1004] : 
                       (N529)? mem[1012] : 
                       (N531)? mem[1020] : 
                       (N278)? mem[1028] : 
                       (N280)? mem[1036] : 
                       (N282)? mem[1044] : 
                       (N284)? mem[1052] : 
                       (N286)? mem[1060] : 
                       (N288)? mem[1068] : 
                       (N290)? mem[1076] : 
                       (N292)? mem[1084] : 
                       (N294)? mem[1092] : 
                       (N296)? mem[1100] : 
                       (N298)? mem[1108] : 
                       (N300)? mem[1116] : 
                       (N302)? mem[1124] : 
                       (N304)? mem[1132] : 
                       (N306)? mem[1140] : 
                       (N308)? mem[1148] : 
                       (N310)? mem[1156] : 
                       (N312)? mem[1164] : 
                       (N314)? mem[1172] : 
                       (N316)? mem[1180] : 
                       (N318)? mem[1188] : 
                       (N320)? mem[1196] : 
                       (N322)? mem[1204] : 
                       (N324)? mem[1212] : 
                       (N326)? mem[1220] : 
                       (N328)? mem[1228] : 
                       (N330)? mem[1236] : 
                       (N332)? mem[1244] : 
                       (N334)? mem[1252] : 
                       (N336)? mem[1260] : 
                       (N338)? mem[1268] : 
                       (N340)? mem[1276] : 
                       (N342)? mem[1284] : 
                       (N344)? mem[1292] : 
                       (N346)? mem[1300] : 
                       (N348)? mem[1308] : 
                       (N350)? mem[1316] : 
                       (N352)? mem[1324] : 
                       (N354)? mem[1332] : 
                       (N356)? mem[1340] : 
                       (N358)? mem[1348] : 
                       (N360)? mem[1356] : 
                       (N362)? mem[1364] : 
                       (N364)? mem[1372] : 
                       (N366)? mem[1380] : 
                       (N368)? mem[1388] : 
                       (N370)? mem[1396] : 
                       (N372)? mem[1404] : 
                       (N374)? mem[1412] : 
                       (N376)? mem[1420] : 
                       (N378)? mem[1428] : 
                       (N380)? mem[1436] : 
                       (N382)? mem[1444] : 
                       (N384)? mem[1452] : 
                       (N386)? mem[1460] : 
                       (N388)? mem[1468] : 
                       (N390)? mem[1476] : 
                       (N392)? mem[1484] : 
                       (N394)? mem[1492] : 
                       (N396)? mem[1500] : 
                       (N398)? mem[1508] : 
                       (N400)? mem[1516] : 
                       (N402)? mem[1524] : 
                       (N404)? mem[1532] : 
                       (N406)? mem[1540] : 
                       (N408)? mem[1548] : 
                       (N410)? mem[1556] : 
                       (N412)? mem[1564] : 
                       (N414)? mem[1572] : 
                       (N416)? mem[1580] : 
                       (N418)? mem[1588] : 
                       (N420)? mem[1596] : 
                       (N422)? mem[1604] : 
                       (N424)? mem[1612] : 
                       (N426)? mem[1620] : 
                       (N428)? mem[1628] : 
                       (N430)? mem[1636] : 
                       (N432)? mem[1644] : 
                       (N434)? mem[1652] : 
                       (N436)? mem[1660] : 
                       (N438)? mem[1668] : 
                       (N440)? mem[1676] : 
                       (N442)? mem[1684] : 
                       (N444)? mem[1692] : 
                       (N446)? mem[1700] : 
                       (N448)? mem[1708] : 
                       (N450)? mem[1716] : 
                       (N452)? mem[1724] : 
                       (N454)? mem[1732] : 
                       (N456)? mem[1740] : 
                       (N458)? mem[1748] : 
                       (N460)? mem[1756] : 
                       (N462)? mem[1764] : 
                       (N464)? mem[1772] : 
                       (N466)? mem[1780] : 
                       (N468)? mem[1788] : 
                       (N470)? mem[1796] : 
                       (N472)? mem[1804] : 
                       (N474)? mem[1812] : 
                       (N476)? mem[1820] : 
                       (N478)? mem[1828] : 
                       (N480)? mem[1836] : 
                       (N482)? mem[1844] : 
                       (N484)? mem[1852] : 
                       (N486)? mem[1860] : 
                       (N488)? mem[1868] : 
                       (N490)? mem[1876] : 
                       (N492)? mem[1884] : 
                       (N494)? mem[1892] : 
                       (N496)? mem[1900] : 
                       (N498)? mem[1908] : 
                       (N500)? mem[1916] : 
                       (N502)? mem[1924] : 
                       (N504)? mem[1932] : 
                       (N506)? mem[1940] : 
                       (N508)? mem[1948] : 
                       (N510)? mem[1956] : 
                       (N512)? mem[1964] : 
                       (N514)? mem[1972] : 
                       (N516)? mem[1980] : 
                       (N518)? mem[1988] : 
                       (N520)? mem[1996] : 
                       (N522)? mem[2004] : 
                       (N524)? mem[2012] : 
                       (N526)? mem[2020] : 
                       (N528)? mem[2028] : 
                       (N530)? mem[2036] : 
                       (N532)? mem[2044] : 1'b0;
  assign data_out[3] = (N277)? mem[3] : 
                       (N279)? mem[11] : 
                       (N281)? mem[19] : 
                       (N283)? mem[27] : 
                       (N285)? mem[35] : 
                       (N287)? mem[43] : 
                       (N289)? mem[51] : 
                       (N291)? mem[59] : 
                       (N293)? mem[67] : 
                       (N295)? mem[75] : 
                       (N297)? mem[83] : 
                       (N299)? mem[91] : 
                       (N301)? mem[99] : 
                       (N303)? mem[107] : 
                       (N305)? mem[115] : 
                       (N307)? mem[123] : 
                       (N309)? mem[131] : 
                       (N311)? mem[139] : 
                       (N313)? mem[147] : 
                       (N315)? mem[155] : 
                       (N317)? mem[163] : 
                       (N319)? mem[171] : 
                       (N321)? mem[179] : 
                       (N323)? mem[187] : 
                       (N325)? mem[195] : 
                       (N327)? mem[203] : 
                       (N329)? mem[211] : 
                       (N331)? mem[219] : 
                       (N333)? mem[227] : 
                       (N335)? mem[235] : 
                       (N337)? mem[243] : 
                       (N339)? mem[251] : 
                       (N341)? mem[259] : 
                       (N343)? mem[267] : 
                       (N345)? mem[275] : 
                       (N347)? mem[283] : 
                       (N349)? mem[291] : 
                       (N351)? mem[299] : 
                       (N353)? mem[307] : 
                       (N355)? mem[315] : 
                       (N357)? mem[323] : 
                       (N359)? mem[331] : 
                       (N361)? mem[339] : 
                       (N363)? mem[347] : 
                       (N365)? mem[355] : 
                       (N367)? mem[363] : 
                       (N369)? mem[371] : 
                       (N371)? mem[379] : 
                       (N373)? mem[387] : 
                       (N375)? mem[395] : 
                       (N377)? mem[403] : 
                       (N379)? mem[411] : 
                       (N381)? mem[419] : 
                       (N383)? mem[427] : 
                       (N385)? mem[435] : 
                       (N387)? mem[443] : 
                       (N389)? mem[451] : 
                       (N391)? mem[459] : 
                       (N393)? mem[467] : 
                       (N395)? mem[475] : 
                       (N397)? mem[483] : 
                       (N399)? mem[491] : 
                       (N401)? mem[499] : 
                       (N403)? mem[507] : 
                       (N405)? mem[515] : 
                       (N407)? mem[523] : 
                       (N409)? mem[531] : 
                       (N411)? mem[539] : 
                       (N413)? mem[547] : 
                       (N415)? mem[555] : 
                       (N417)? mem[563] : 
                       (N419)? mem[571] : 
                       (N421)? mem[579] : 
                       (N423)? mem[587] : 
                       (N425)? mem[595] : 
                       (N427)? mem[603] : 
                       (N429)? mem[611] : 
                       (N431)? mem[619] : 
                       (N433)? mem[627] : 
                       (N435)? mem[635] : 
                       (N437)? mem[643] : 
                       (N439)? mem[651] : 
                       (N441)? mem[659] : 
                       (N443)? mem[667] : 
                       (N445)? mem[675] : 
                       (N447)? mem[683] : 
                       (N449)? mem[691] : 
                       (N451)? mem[699] : 
                       (N453)? mem[707] : 
                       (N455)? mem[715] : 
                       (N457)? mem[723] : 
                       (N459)? mem[731] : 
                       (N461)? mem[739] : 
                       (N463)? mem[747] : 
                       (N465)? mem[755] : 
                       (N467)? mem[763] : 
                       (N469)? mem[771] : 
                       (N471)? mem[779] : 
                       (N473)? mem[787] : 
                       (N475)? mem[795] : 
                       (N477)? mem[803] : 
                       (N479)? mem[811] : 
                       (N481)? mem[819] : 
                       (N483)? mem[827] : 
                       (N485)? mem[835] : 
                       (N487)? mem[843] : 
                       (N489)? mem[851] : 
                       (N491)? mem[859] : 
                       (N493)? mem[867] : 
                       (N495)? mem[875] : 
                       (N497)? mem[883] : 
                       (N499)? mem[891] : 
                       (N501)? mem[899] : 
                       (N503)? mem[907] : 
                       (N505)? mem[915] : 
                       (N507)? mem[923] : 
                       (N509)? mem[931] : 
                       (N511)? mem[939] : 
                       (N513)? mem[947] : 
                       (N515)? mem[955] : 
                       (N517)? mem[963] : 
                       (N519)? mem[971] : 
                       (N521)? mem[979] : 
                       (N523)? mem[987] : 
                       (N525)? mem[995] : 
                       (N527)? mem[1003] : 
                       (N529)? mem[1011] : 
                       (N531)? mem[1019] : 
                       (N278)? mem[1027] : 
                       (N280)? mem[1035] : 
                       (N282)? mem[1043] : 
                       (N284)? mem[1051] : 
                       (N286)? mem[1059] : 
                       (N288)? mem[1067] : 
                       (N290)? mem[1075] : 
                       (N292)? mem[1083] : 
                       (N294)? mem[1091] : 
                       (N296)? mem[1099] : 
                       (N298)? mem[1107] : 
                       (N300)? mem[1115] : 
                       (N302)? mem[1123] : 
                       (N304)? mem[1131] : 
                       (N306)? mem[1139] : 
                       (N308)? mem[1147] : 
                       (N310)? mem[1155] : 
                       (N312)? mem[1163] : 
                       (N314)? mem[1171] : 
                       (N316)? mem[1179] : 
                       (N318)? mem[1187] : 
                       (N320)? mem[1195] : 
                       (N322)? mem[1203] : 
                       (N324)? mem[1211] : 
                       (N326)? mem[1219] : 
                       (N328)? mem[1227] : 
                       (N330)? mem[1235] : 
                       (N332)? mem[1243] : 
                       (N334)? mem[1251] : 
                       (N336)? mem[1259] : 
                       (N338)? mem[1267] : 
                       (N340)? mem[1275] : 
                       (N342)? mem[1283] : 
                       (N344)? mem[1291] : 
                       (N346)? mem[1299] : 
                       (N348)? mem[1307] : 
                       (N350)? mem[1315] : 
                       (N352)? mem[1323] : 
                       (N354)? mem[1331] : 
                       (N356)? mem[1339] : 
                       (N358)? mem[1347] : 
                       (N360)? mem[1355] : 
                       (N362)? mem[1363] : 
                       (N364)? mem[1371] : 
                       (N366)? mem[1379] : 
                       (N368)? mem[1387] : 
                       (N370)? mem[1395] : 
                       (N372)? mem[1403] : 
                       (N374)? mem[1411] : 
                       (N376)? mem[1419] : 
                       (N378)? mem[1427] : 
                       (N380)? mem[1435] : 
                       (N382)? mem[1443] : 
                       (N384)? mem[1451] : 
                       (N386)? mem[1459] : 
                       (N388)? mem[1467] : 
                       (N390)? mem[1475] : 
                       (N392)? mem[1483] : 
                       (N394)? mem[1491] : 
                       (N396)? mem[1499] : 
                       (N398)? mem[1507] : 
                       (N400)? mem[1515] : 
                       (N402)? mem[1523] : 
                       (N404)? mem[1531] : 
                       (N406)? mem[1539] : 
                       (N408)? mem[1547] : 
                       (N410)? mem[1555] : 
                       (N412)? mem[1563] : 
                       (N414)? mem[1571] : 
                       (N416)? mem[1579] : 
                       (N418)? mem[1587] : 
                       (N420)? mem[1595] : 
                       (N422)? mem[1603] : 
                       (N424)? mem[1611] : 
                       (N426)? mem[1619] : 
                       (N428)? mem[1627] : 
                       (N430)? mem[1635] : 
                       (N432)? mem[1643] : 
                       (N434)? mem[1651] : 
                       (N436)? mem[1659] : 
                       (N438)? mem[1667] : 
                       (N440)? mem[1675] : 
                       (N442)? mem[1683] : 
                       (N444)? mem[1691] : 
                       (N446)? mem[1699] : 
                       (N448)? mem[1707] : 
                       (N450)? mem[1715] : 
                       (N452)? mem[1723] : 
                       (N454)? mem[1731] : 
                       (N456)? mem[1739] : 
                       (N458)? mem[1747] : 
                       (N460)? mem[1755] : 
                       (N462)? mem[1763] : 
                       (N464)? mem[1771] : 
                       (N466)? mem[1779] : 
                       (N468)? mem[1787] : 
                       (N470)? mem[1795] : 
                       (N472)? mem[1803] : 
                       (N474)? mem[1811] : 
                       (N476)? mem[1819] : 
                       (N478)? mem[1827] : 
                       (N480)? mem[1835] : 
                       (N482)? mem[1843] : 
                       (N484)? mem[1851] : 
                       (N486)? mem[1859] : 
                       (N488)? mem[1867] : 
                       (N490)? mem[1875] : 
                       (N492)? mem[1883] : 
                       (N494)? mem[1891] : 
                       (N496)? mem[1899] : 
                       (N498)? mem[1907] : 
                       (N500)? mem[1915] : 
                       (N502)? mem[1923] : 
                       (N504)? mem[1931] : 
                       (N506)? mem[1939] : 
                       (N508)? mem[1947] : 
                       (N510)? mem[1955] : 
                       (N512)? mem[1963] : 
                       (N514)? mem[1971] : 
                       (N516)? mem[1979] : 
                       (N518)? mem[1987] : 
                       (N520)? mem[1995] : 
                       (N522)? mem[2003] : 
                       (N524)? mem[2011] : 
                       (N526)? mem[2019] : 
                       (N528)? mem[2027] : 
                       (N530)? mem[2035] : 
                       (N532)? mem[2043] : 1'b0;
  assign data_out[2] = (N277)? mem[2] : 
                       (N279)? mem[10] : 
                       (N281)? mem[18] : 
                       (N283)? mem[26] : 
                       (N285)? mem[34] : 
                       (N287)? mem[42] : 
                       (N289)? mem[50] : 
                       (N291)? mem[58] : 
                       (N293)? mem[66] : 
                       (N295)? mem[74] : 
                       (N297)? mem[82] : 
                       (N299)? mem[90] : 
                       (N301)? mem[98] : 
                       (N303)? mem[106] : 
                       (N305)? mem[114] : 
                       (N307)? mem[122] : 
                       (N309)? mem[130] : 
                       (N311)? mem[138] : 
                       (N313)? mem[146] : 
                       (N315)? mem[154] : 
                       (N317)? mem[162] : 
                       (N319)? mem[170] : 
                       (N321)? mem[178] : 
                       (N323)? mem[186] : 
                       (N325)? mem[194] : 
                       (N327)? mem[202] : 
                       (N329)? mem[210] : 
                       (N331)? mem[218] : 
                       (N333)? mem[226] : 
                       (N335)? mem[234] : 
                       (N337)? mem[242] : 
                       (N339)? mem[250] : 
                       (N341)? mem[258] : 
                       (N343)? mem[266] : 
                       (N345)? mem[274] : 
                       (N347)? mem[282] : 
                       (N349)? mem[290] : 
                       (N351)? mem[298] : 
                       (N353)? mem[306] : 
                       (N355)? mem[314] : 
                       (N357)? mem[322] : 
                       (N359)? mem[330] : 
                       (N361)? mem[338] : 
                       (N363)? mem[346] : 
                       (N365)? mem[354] : 
                       (N367)? mem[362] : 
                       (N369)? mem[370] : 
                       (N371)? mem[378] : 
                       (N373)? mem[386] : 
                       (N375)? mem[394] : 
                       (N377)? mem[402] : 
                       (N379)? mem[410] : 
                       (N381)? mem[418] : 
                       (N383)? mem[426] : 
                       (N385)? mem[434] : 
                       (N387)? mem[442] : 
                       (N389)? mem[450] : 
                       (N391)? mem[458] : 
                       (N393)? mem[466] : 
                       (N395)? mem[474] : 
                       (N397)? mem[482] : 
                       (N399)? mem[490] : 
                       (N401)? mem[498] : 
                       (N403)? mem[506] : 
                       (N405)? mem[514] : 
                       (N407)? mem[522] : 
                       (N409)? mem[530] : 
                       (N411)? mem[538] : 
                       (N413)? mem[546] : 
                       (N415)? mem[554] : 
                       (N417)? mem[562] : 
                       (N419)? mem[570] : 
                       (N421)? mem[578] : 
                       (N423)? mem[586] : 
                       (N425)? mem[594] : 
                       (N427)? mem[602] : 
                       (N429)? mem[610] : 
                       (N431)? mem[618] : 
                       (N433)? mem[626] : 
                       (N435)? mem[634] : 
                       (N437)? mem[642] : 
                       (N439)? mem[650] : 
                       (N441)? mem[658] : 
                       (N443)? mem[666] : 
                       (N445)? mem[674] : 
                       (N447)? mem[682] : 
                       (N449)? mem[690] : 
                       (N451)? mem[698] : 
                       (N453)? mem[706] : 
                       (N455)? mem[714] : 
                       (N457)? mem[722] : 
                       (N459)? mem[730] : 
                       (N461)? mem[738] : 
                       (N463)? mem[746] : 
                       (N465)? mem[754] : 
                       (N467)? mem[762] : 
                       (N469)? mem[770] : 
                       (N471)? mem[778] : 
                       (N473)? mem[786] : 
                       (N475)? mem[794] : 
                       (N477)? mem[802] : 
                       (N479)? mem[810] : 
                       (N481)? mem[818] : 
                       (N483)? mem[826] : 
                       (N485)? mem[834] : 
                       (N487)? mem[842] : 
                       (N489)? mem[850] : 
                       (N491)? mem[858] : 
                       (N493)? mem[866] : 
                       (N495)? mem[874] : 
                       (N497)? mem[882] : 
                       (N499)? mem[890] : 
                       (N501)? mem[898] : 
                       (N503)? mem[906] : 
                       (N505)? mem[914] : 
                       (N507)? mem[922] : 
                       (N509)? mem[930] : 
                       (N511)? mem[938] : 
                       (N513)? mem[946] : 
                       (N515)? mem[954] : 
                       (N517)? mem[962] : 
                       (N519)? mem[970] : 
                       (N521)? mem[978] : 
                       (N523)? mem[986] : 
                       (N525)? mem[994] : 
                       (N527)? mem[1002] : 
                       (N529)? mem[1010] : 
                       (N531)? mem[1018] : 
                       (N278)? mem[1026] : 
                       (N280)? mem[1034] : 
                       (N282)? mem[1042] : 
                       (N284)? mem[1050] : 
                       (N286)? mem[1058] : 
                       (N288)? mem[1066] : 
                       (N290)? mem[1074] : 
                       (N292)? mem[1082] : 
                       (N294)? mem[1090] : 
                       (N296)? mem[1098] : 
                       (N298)? mem[1106] : 
                       (N300)? mem[1114] : 
                       (N302)? mem[1122] : 
                       (N304)? mem[1130] : 
                       (N306)? mem[1138] : 
                       (N308)? mem[1146] : 
                       (N310)? mem[1154] : 
                       (N312)? mem[1162] : 
                       (N314)? mem[1170] : 
                       (N316)? mem[1178] : 
                       (N318)? mem[1186] : 
                       (N320)? mem[1194] : 
                       (N322)? mem[1202] : 
                       (N324)? mem[1210] : 
                       (N326)? mem[1218] : 
                       (N328)? mem[1226] : 
                       (N330)? mem[1234] : 
                       (N332)? mem[1242] : 
                       (N334)? mem[1250] : 
                       (N336)? mem[1258] : 
                       (N338)? mem[1266] : 
                       (N340)? mem[1274] : 
                       (N342)? mem[1282] : 
                       (N344)? mem[1290] : 
                       (N346)? mem[1298] : 
                       (N348)? mem[1306] : 
                       (N350)? mem[1314] : 
                       (N352)? mem[1322] : 
                       (N354)? mem[1330] : 
                       (N356)? mem[1338] : 
                       (N358)? mem[1346] : 
                       (N360)? mem[1354] : 
                       (N362)? mem[1362] : 
                       (N364)? mem[1370] : 
                       (N366)? mem[1378] : 
                       (N368)? mem[1386] : 
                       (N370)? mem[1394] : 
                       (N372)? mem[1402] : 
                       (N374)? mem[1410] : 
                       (N376)? mem[1418] : 
                       (N378)? mem[1426] : 
                       (N380)? mem[1434] : 
                       (N382)? mem[1442] : 
                       (N384)? mem[1450] : 
                       (N386)? mem[1458] : 
                       (N388)? mem[1466] : 
                       (N390)? mem[1474] : 
                       (N392)? mem[1482] : 
                       (N394)? mem[1490] : 
                       (N396)? mem[1498] : 
                       (N398)? mem[1506] : 
                       (N400)? mem[1514] : 
                       (N402)? mem[1522] : 
                       (N404)? mem[1530] : 
                       (N406)? mem[1538] : 
                       (N408)? mem[1546] : 
                       (N410)? mem[1554] : 
                       (N412)? mem[1562] : 
                       (N414)? mem[1570] : 
                       (N416)? mem[1578] : 
                       (N418)? mem[1586] : 
                       (N420)? mem[1594] : 
                       (N422)? mem[1602] : 
                       (N424)? mem[1610] : 
                       (N426)? mem[1618] : 
                       (N428)? mem[1626] : 
                       (N430)? mem[1634] : 
                       (N432)? mem[1642] : 
                       (N434)? mem[1650] : 
                       (N436)? mem[1658] : 
                       (N438)? mem[1666] : 
                       (N440)? mem[1674] : 
                       (N442)? mem[1682] : 
                       (N444)? mem[1690] : 
                       (N446)? mem[1698] : 
                       (N448)? mem[1706] : 
                       (N450)? mem[1714] : 
                       (N452)? mem[1722] : 
                       (N454)? mem[1730] : 
                       (N456)? mem[1738] : 
                       (N458)? mem[1746] : 
                       (N460)? mem[1754] : 
                       (N462)? mem[1762] : 
                       (N464)? mem[1770] : 
                       (N466)? mem[1778] : 
                       (N468)? mem[1786] : 
                       (N470)? mem[1794] : 
                       (N472)? mem[1802] : 
                       (N474)? mem[1810] : 
                       (N476)? mem[1818] : 
                       (N478)? mem[1826] : 
                       (N480)? mem[1834] : 
                       (N482)? mem[1842] : 
                       (N484)? mem[1850] : 
                       (N486)? mem[1858] : 
                       (N488)? mem[1866] : 
                       (N490)? mem[1874] : 
                       (N492)? mem[1882] : 
                       (N494)? mem[1890] : 
                       (N496)? mem[1898] : 
                       (N498)? mem[1906] : 
                       (N500)? mem[1914] : 
                       (N502)? mem[1922] : 
                       (N504)? mem[1930] : 
                       (N506)? mem[1938] : 
                       (N508)? mem[1946] : 
                       (N510)? mem[1954] : 
                       (N512)? mem[1962] : 
                       (N514)? mem[1970] : 
                       (N516)? mem[1978] : 
                       (N518)? mem[1986] : 
                       (N520)? mem[1994] : 
                       (N522)? mem[2002] : 
                       (N524)? mem[2010] : 
                       (N526)? mem[2018] : 
                       (N528)? mem[2026] : 
                       (N530)? mem[2034] : 
                       (N532)? mem[2042] : 1'b0;
  assign data_out[1] = (N277)? mem[1] : 
                       (N279)? mem[9] : 
                       (N281)? mem[17] : 
                       (N283)? mem[25] : 
                       (N285)? mem[33] : 
                       (N287)? mem[41] : 
                       (N289)? mem[49] : 
                       (N291)? mem[57] : 
                       (N293)? mem[65] : 
                       (N295)? mem[73] : 
                       (N297)? mem[81] : 
                       (N299)? mem[89] : 
                       (N301)? mem[97] : 
                       (N303)? mem[105] : 
                       (N305)? mem[113] : 
                       (N307)? mem[121] : 
                       (N309)? mem[129] : 
                       (N311)? mem[137] : 
                       (N313)? mem[145] : 
                       (N315)? mem[153] : 
                       (N317)? mem[161] : 
                       (N319)? mem[169] : 
                       (N321)? mem[177] : 
                       (N323)? mem[185] : 
                       (N325)? mem[193] : 
                       (N327)? mem[201] : 
                       (N329)? mem[209] : 
                       (N331)? mem[217] : 
                       (N333)? mem[225] : 
                       (N335)? mem[233] : 
                       (N337)? mem[241] : 
                       (N339)? mem[249] : 
                       (N341)? mem[257] : 
                       (N343)? mem[265] : 
                       (N345)? mem[273] : 
                       (N347)? mem[281] : 
                       (N349)? mem[289] : 
                       (N351)? mem[297] : 
                       (N353)? mem[305] : 
                       (N355)? mem[313] : 
                       (N357)? mem[321] : 
                       (N359)? mem[329] : 
                       (N361)? mem[337] : 
                       (N363)? mem[345] : 
                       (N365)? mem[353] : 
                       (N367)? mem[361] : 
                       (N369)? mem[369] : 
                       (N371)? mem[377] : 
                       (N373)? mem[385] : 
                       (N375)? mem[393] : 
                       (N377)? mem[401] : 
                       (N379)? mem[409] : 
                       (N381)? mem[417] : 
                       (N383)? mem[425] : 
                       (N385)? mem[433] : 
                       (N387)? mem[441] : 
                       (N389)? mem[449] : 
                       (N391)? mem[457] : 
                       (N393)? mem[465] : 
                       (N395)? mem[473] : 
                       (N397)? mem[481] : 
                       (N399)? mem[489] : 
                       (N401)? mem[497] : 
                       (N403)? mem[505] : 
                       (N405)? mem[513] : 
                       (N407)? mem[521] : 
                       (N409)? mem[529] : 
                       (N411)? mem[537] : 
                       (N413)? mem[545] : 
                       (N415)? mem[553] : 
                       (N417)? mem[561] : 
                       (N419)? mem[569] : 
                       (N421)? mem[577] : 
                       (N423)? mem[585] : 
                       (N425)? mem[593] : 
                       (N427)? mem[601] : 
                       (N429)? mem[609] : 
                       (N431)? mem[617] : 
                       (N433)? mem[625] : 
                       (N435)? mem[633] : 
                       (N437)? mem[641] : 
                       (N439)? mem[649] : 
                       (N441)? mem[657] : 
                       (N443)? mem[665] : 
                       (N445)? mem[673] : 
                       (N447)? mem[681] : 
                       (N449)? mem[689] : 
                       (N451)? mem[697] : 
                       (N453)? mem[705] : 
                       (N455)? mem[713] : 
                       (N457)? mem[721] : 
                       (N459)? mem[729] : 
                       (N461)? mem[737] : 
                       (N463)? mem[745] : 
                       (N465)? mem[753] : 
                       (N467)? mem[761] : 
                       (N469)? mem[769] : 
                       (N471)? mem[777] : 
                       (N473)? mem[785] : 
                       (N475)? mem[793] : 
                       (N477)? mem[801] : 
                       (N479)? mem[809] : 
                       (N481)? mem[817] : 
                       (N483)? mem[825] : 
                       (N485)? mem[833] : 
                       (N487)? mem[841] : 
                       (N489)? mem[849] : 
                       (N491)? mem[857] : 
                       (N493)? mem[865] : 
                       (N495)? mem[873] : 
                       (N497)? mem[881] : 
                       (N499)? mem[889] : 
                       (N501)? mem[897] : 
                       (N503)? mem[905] : 
                       (N505)? mem[913] : 
                       (N507)? mem[921] : 
                       (N509)? mem[929] : 
                       (N511)? mem[937] : 
                       (N513)? mem[945] : 
                       (N515)? mem[953] : 
                       (N517)? mem[961] : 
                       (N519)? mem[969] : 
                       (N521)? mem[977] : 
                       (N523)? mem[985] : 
                       (N525)? mem[993] : 
                       (N527)? mem[1001] : 
                       (N529)? mem[1009] : 
                       (N531)? mem[1017] : 
                       (N278)? mem[1025] : 
                       (N280)? mem[1033] : 
                       (N282)? mem[1041] : 
                       (N284)? mem[1049] : 
                       (N286)? mem[1057] : 
                       (N288)? mem[1065] : 
                       (N290)? mem[1073] : 
                       (N292)? mem[1081] : 
                       (N294)? mem[1089] : 
                       (N296)? mem[1097] : 
                       (N298)? mem[1105] : 
                       (N300)? mem[1113] : 
                       (N302)? mem[1121] : 
                       (N304)? mem[1129] : 
                       (N306)? mem[1137] : 
                       (N308)? mem[1145] : 
                       (N310)? mem[1153] : 
                       (N312)? mem[1161] : 
                       (N314)? mem[1169] : 
                       (N316)? mem[1177] : 
                       (N318)? mem[1185] : 
                       (N320)? mem[1193] : 
                       (N322)? mem[1201] : 
                       (N324)? mem[1209] : 
                       (N326)? mem[1217] : 
                       (N328)? mem[1225] : 
                       (N330)? mem[1233] : 
                       (N332)? mem[1241] : 
                       (N334)? mem[1249] : 
                       (N336)? mem[1257] : 
                       (N338)? mem[1265] : 
                       (N340)? mem[1273] : 
                       (N342)? mem[1281] : 
                       (N344)? mem[1289] : 
                       (N346)? mem[1297] : 
                       (N348)? mem[1305] : 
                       (N350)? mem[1313] : 
                       (N352)? mem[1321] : 
                       (N354)? mem[1329] : 
                       (N356)? mem[1337] : 
                       (N358)? mem[1345] : 
                       (N360)? mem[1353] : 
                       (N362)? mem[1361] : 
                       (N364)? mem[1369] : 
                       (N366)? mem[1377] : 
                       (N368)? mem[1385] : 
                       (N370)? mem[1393] : 
                       (N372)? mem[1401] : 
                       (N374)? mem[1409] : 
                       (N376)? mem[1417] : 
                       (N378)? mem[1425] : 
                       (N380)? mem[1433] : 
                       (N382)? mem[1441] : 
                       (N384)? mem[1449] : 
                       (N386)? mem[1457] : 
                       (N388)? mem[1465] : 
                       (N390)? mem[1473] : 
                       (N392)? mem[1481] : 
                       (N394)? mem[1489] : 
                       (N396)? mem[1497] : 
                       (N398)? mem[1505] : 
                       (N400)? mem[1513] : 
                       (N402)? mem[1521] : 
                       (N404)? mem[1529] : 
                       (N406)? mem[1537] : 
                       (N408)? mem[1545] : 
                       (N410)? mem[1553] : 
                       (N412)? mem[1561] : 
                       (N414)? mem[1569] : 
                       (N416)? mem[1577] : 
                       (N418)? mem[1585] : 
                       (N420)? mem[1593] : 
                       (N422)? mem[1601] : 
                       (N424)? mem[1609] : 
                       (N426)? mem[1617] : 
                       (N428)? mem[1625] : 
                       (N430)? mem[1633] : 
                       (N432)? mem[1641] : 
                       (N434)? mem[1649] : 
                       (N436)? mem[1657] : 
                       (N438)? mem[1665] : 
                       (N440)? mem[1673] : 
                       (N442)? mem[1681] : 
                       (N444)? mem[1689] : 
                       (N446)? mem[1697] : 
                       (N448)? mem[1705] : 
                       (N450)? mem[1713] : 
                       (N452)? mem[1721] : 
                       (N454)? mem[1729] : 
                       (N456)? mem[1737] : 
                       (N458)? mem[1745] : 
                       (N460)? mem[1753] : 
                       (N462)? mem[1761] : 
                       (N464)? mem[1769] : 
                       (N466)? mem[1777] : 
                       (N468)? mem[1785] : 
                       (N470)? mem[1793] : 
                       (N472)? mem[1801] : 
                       (N474)? mem[1809] : 
                       (N476)? mem[1817] : 
                       (N478)? mem[1825] : 
                       (N480)? mem[1833] : 
                       (N482)? mem[1841] : 
                       (N484)? mem[1849] : 
                       (N486)? mem[1857] : 
                       (N488)? mem[1865] : 
                       (N490)? mem[1873] : 
                       (N492)? mem[1881] : 
                       (N494)? mem[1889] : 
                       (N496)? mem[1897] : 
                       (N498)? mem[1905] : 
                       (N500)? mem[1913] : 
                       (N502)? mem[1921] : 
                       (N504)? mem[1929] : 
                       (N506)? mem[1937] : 
                       (N508)? mem[1945] : 
                       (N510)? mem[1953] : 
                       (N512)? mem[1961] : 
                       (N514)? mem[1969] : 
                       (N516)? mem[1977] : 
                       (N518)? mem[1985] : 
                       (N520)? mem[1993] : 
                       (N522)? mem[2001] : 
                       (N524)? mem[2009] : 
                       (N526)? mem[2017] : 
                       (N528)? mem[2025] : 
                       (N530)? mem[2033] : 
                       (N532)? mem[2041] : 1'b0;
  assign data_out[0] = (N277)? mem[0] : 
                       (N279)? mem[8] : 
                       (N281)? mem[16] : 
                       (N283)? mem[24] : 
                       (N285)? mem[32] : 
                       (N287)? mem[40] : 
                       (N289)? mem[48] : 
                       (N291)? mem[56] : 
                       (N293)? mem[64] : 
                       (N295)? mem[72] : 
                       (N297)? mem[80] : 
                       (N299)? mem[88] : 
                       (N301)? mem[96] : 
                       (N303)? mem[104] : 
                       (N305)? mem[112] : 
                       (N307)? mem[120] : 
                       (N309)? mem[128] : 
                       (N311)? mem[136] : 
                       (N313)? mem[144] : 
                       (N315)? mem[152] : 
                       (N317)? mem[160] : 
                       (N319)? mem[168] : 
                       (N321)? mem[176] : 
                       (N323)? mem[184] : 
                       (N325)? mem[192] : 
                       (N327)? mem[200] : 
                       (N329)? mem[208] : 
                       (N331)? mem[216] : 
                       (N333)? mem[224] : 
                       (N335)? mem[232] : 
                       (N337)? mem[240] : 
                       (N339)? mem[248] : 
                       (N341)? mem[256] : 
                       (N343)? mem[264] : 
                       (N345)? mem[272] : 
                       (N347)? mem[280] : 
                       (N349)? mem[288] : 
                       (N351)? mem[296] : 
                       (N353)? mem[304] : 
                       (N355)? mem[312] : 
                       (N357)? mem[320] : 
                       (N359)? mem[328] : 
                       (N361)? mem[336] : 
                       (N363)? mem[344] : 
                       (N365)? mem[352] : 
                       (N367)? mem[360] : 
                       (N369)? mem[368] : 
                       (N371)? mem[376] : 
                       (N373)? mem[384] : 
                       (N375)? mem[392] : 
                       (N377)? mem[400] : 
                       (N379)? mem[408] : 
                       (N381)? mem[416] : 
                       (N383)? mem[424] : 
                       (N385)? mem[432] : 
                       (N387)? mem[440] : 
                       (N389)? mem[448] : 
                       (N391)? mem[456] : 
                       (N393)? mem[464] : 
                       (N395)? mem[472] : 
                       (N397)? mem[480] : 
                       (N399)? mem[488] : 
                       (N401)? mem[496] : 
                       (N403)? mem[504] : 
                       (N405)? mem[512] : 
                       (N407)? mem[520] : 
                       (N409)? mem[528] : 
                       (N411)? mem[536] : 
                       (N413)? mem[544] : 
                       (N415)? mem[552] : 
                       (N417)? mem[560] : 
                       (N419)? mem[568] : 
                       (N421)? mem[576] : 
                       (N423)? mem[584] : 
                       (N425)? mem[592] : 
                       (N427)? mem[600] : 
                       (N429)? mem[608] : 
                       (N431)? mem[616] : 
                       (N433)? mem[624] : 
                       (N435)? mem[632] : 
                       (N437)? mem[640] : 
                       (N439)? mem[648] : 
                       (N441)? mem[656] : 
                       (N443)? mem[664] : 
                       (N445)? mem[672] : 
                       (N447)? mem[680] : 
                       (N449)? mem[688] : 
                       (N451)? mem[696] : 
                       (N453)? mem[704] : 
                       (N455)? mem[712] : 
                       (N457)? mem[720] : 
                       (N459)? mem[728] : 
                       (N461)? mem[736] : 
                       (N463)? mem[744] : 
                       (N465)? mem[752] : 
                       (N467)? mem[760] : 
                       (N469)? mem[768] : 
                       (N471)? mem[776] : 
                       (N473)? mem[784] : 
                       (N475)? mem[792] : 
                       (N477)? mem[800] : 
                       (N479)? mem[808] : 
                       (N481)? mem[816] : 
                       (N483)? mem[824] : 
                       (N485)? mem[832] : 
                       (N487)? mem[840] : 
                       (N489)? mem[848] : 
                       (N491)? mem[856] : 
                       (N493)? mem[864] : 
                       (N495)? mem[872] : 
                       (N497)? mem[880] : 
                       (N499)? mem[888] : 
                       (N501)? mem[896] : 
                       (N503)? mem[904] : 
                       (N505)? mem[912] : 
                       (N507)? mem[920] : 
                       (N509)? mem[928] : 
                       (N511)? mem[936] : 
                       (N513)? mem[944] : 
                       (N515)? mem[952] : 
                       (N517)? mem[960] : 
                       (N519)? mem[968] : 
                       (N521)? mem[976] : 
                       (N523)? mem[984] : 
                       (N525)? mem[992] : 
                       (N527)? mem[1000] : 
                       (N529)? mem[1008] : 
                       (N531)? mem[1016] : 
                       (N278)? mem[1024] : 
                       (N280)? mem[1032] : 
                       (N282)? mem[1040] : 
                       (N284)? mem[1048] : 
                       (N286)? mem[1056] : 
                       (N288)? mem[1064] : 
                       (N290)? mem[1072] : 
                       (N292)? mem[1080] : 
                       (N294)? mem[1088] : 
                       (N296)? mem[1096] : 
                       (N298)? mem[1104] : 
                       (N300)? mem[1112] : 
                       (N302)? mem[1120] : 
                       (N304)? mem[1128] : 
                       (N306)? mem[1136] : 
                       (N308)? mem[1144] : 
                       (N310)? mem[1152] : 
                       (N312)? mem[1160] : 
                       (N314)? mem[1168] : 
                       (N316)? mem[1176] : 
                       (N318)? mem[1184] : 
                       (N320)? mem[1192] : 
                       (N322)? mem[1200] : 
                       (N324)? mem[1208] : 
                       (N326)? mem[1216] : 
                       (N328)? mem[1224] : 
                       (N330)? mem[1232] : 
                       (N332)? mem[1240] : 
                       (N334)? mem[1248] : 
                       (N336)? mem[1256] : 
                       (N338)? mem[1264] : 
                       (N340)? mem[1272] : 
                       (N342)? mem[1280] : 
                       (N344)? mem[1288] : 
                       (N346)? mem[1296] : 
                       (N348)? mem[1304] : 
                       (N350)? mem[1312] : 
                       (N352)? mem[1320] : 
                       (N354)? mem[1328] : 
                       (N356)? mem[1336] : 
                       (N358)? mem[1344] : 
                       (N360)? mem[1352] : 
                       (N362)? mem[1360] : 
                       (N364)? mem[1368] : 
                       (N366)? mem[1376] : 
                       (N368)? mem[1384] : 
                       (N370)? mem[1392] : 
                       (N372)? mem[1400] : 
                       (N374)? mem[1408] : 
                       (N376)? mem[1416] : 
                       (N378)? mem[1424] : 
                       (N380)? mem[1432] : 
                       (N382)? mem[1440] : 
                       (N384)? mem[1448] : 
                       (N386)? mem[1456] : 
                       (N388)? mem[1464] : 
                       (N390)? mem[1472] : 
                       (N392)? mem[1480] : 
                       (N394)? mem[1488] : 
                       (N396)? mem[1496] : 
                       (N398)? mem[1504] : 
                       (N400)? mem[1512] : 
                       (N402)? mem[1520] : 
                       (N404)? mem[1528] : 
                       (N406)? mem[1536] : 
                       (N408)? mem[1544] : 
                       (N410)? mem[1552] : 
                       (N412)? mem[1560] : 
                       (N414)? mem[1568] : 
                       (N416)? mem[1576] : 
                       (N418)? mem[1584] : 
                       (N420)? mem[1592] : 
                       (N422)? mem[1600] : 
                       (N424)? mem[1608] : 
                       (N426)? mem[1616] : 
                       (N428)? mem[1624] : 
                       (N430)? mem[1632] : 
                       (N432)? mem[1640] : 
                       (N434)? mem[1648] : 
                       (N436)? mem[1656] : 
                       (N438)? mem[1664] : 
                       (N440)? mem[1672] : 
                       (N442)? mem[1680] : 
                       (N444)? mem[1688] : 
                       (N446)? mem[1696] : 
                       (N448)? mem[1704] : 
                       (N450)? mem[1712] : 
                       (N452)? mem[1720] : 
                       (N454)? mem[1728] : 
                       (N456)? mem[1736] : 
                       (N458)? mem[1744] : 
                       (N460)? mem[1752] : 
                       (N462)? mem[1760] : 
                       (N464)? mem[1768] : 
                       (N466)? mem[1776] : 
                       (N468)? mem[1784] : 
                       (N470)? mem[1792] : 
                       (N472)? mem[1800] : 
                       (N474)? mem[1808] : 
                       (N476)? mem[1816] : 
                       (N478)? mem[1824] : 
                       (N480)? mem[1832] : 
                       (N482)? mem[1840] : 
                       (N484)? mem[1848] : 
                       (N486)? mem[1856] : 
                       (N488)? mem[1864] : 
                       (N490)? mem[1872] : 
                       (N492)? mem[1880] : 
                       (N494)? mem[1888] : 
                       (N496)? mem[1896] : 
                       (N498)? mem[1904] : 
                       (N500)? mem[1912] : 
                       (N502)? mem[1920] : 
                       (N504)? mem[1928] : 
                       (N506)? mem[1936] : 
                       (N508)? mem[1944] : 
                       (N510)? mem[1952] : 
                       (N512)? mem[1960] : 
                       (N514)? mem[1968] : 
                       (N516)? mem[1976] : 
                       (N518)? mem[1984] : 
                       (N520)? mem[1992] : 
                       (N522)? mem[2000] : 
                       (N524)? mem[2008] : 
                       (N526)? mem[2016] : 
                       (N528)? mem[2024] : 
                       (N530)? mem[2032] : 
                       (N532)? mem[2040] : 1'b0;

  bsg_dff_width_p1
  llr_read_en_dff
  (
    .clk_i(clk_i),
    .data_i(read_en),
    .data_o(llr_read_en_r)
  );


  bsg_dff_en_bypass_width_p8
  llr_dff_bypass
  (
    .clk_i(clk_i),
    .en_i(llr_read_en_r),
    .data_i(data_out),
    .data_o(data_o)
  );

  assign N1047 = addr_i[6] & addr_i[7];
  assign N1048 = N0 & addr_i[7];
  assign N0 = ~addr_i[6];
  assign N1049 = addr_i[6] & N1;
  assign N1 = ~addr_i[7];
  assign N1050 = N2 & N3;
  assign N2 = ~addr_i[6];
  assign N3 = ~addr_i[7];
  assign N1051 = addr_i[4] & addr_i[5];
  assign N1052 = N4 & addr_i[5];
  assign N4 = ~addr_i[4];
  assign N1053 = addr_i[4] & N5;
  assign N5 = ~addr_i[5];
  assign N1054 = N6 & N7;
  assign N6 = ~addr_i[4];
  assign N7 = ~addr_i[5];
  assign N1055 = N1047 & N1051;
  assign N1056 = N1047 & N1052;
  assign N1057 = N1047 & N1053;
  assign N1058 = N1047 & N1054;
  assign N1059 = N1048 & N1051;
  assign N1060 = N1048 & N1052;
  assign N1061 = N1048 & N1053;
  assign N1062 = N1048 & N1054;
  assign N1063 = N1049 & N1051;
  assign N1064 = N1049 & N1052;
  assign N1065 = N1049 & N1053;
  assign N1066 = N1049 & N1054;
  assign N1067 = N1050 & N1051;
  assign N1068 = N1050 & N1052;
  assign N1069 = N1050 & N1053;
  assign N1070 = N1050 & N1054;
  assign N1071 = addr_i[2] & addr_i[3];
  assign N1072 = N8 & addr_i[3];
  assign N8 = ~addr_i[2];
  assign N1073 = addr_i[2] & N9;
  assign N9 = ~addr_i[3];
  assign N1074 = N10 & N11;
  assign N10 = ~addr_i[2];
  assign N11 = ~addr_i[3];
  assign N1075 = addr_i[0] & addr_i[1];
  assign N1076 = N12 & addr_i[1];
  assign N12 = ~addr_i[0];
  assign N1077 = addr_i[0] & N13;
  assign N13 = ~addr_i[1];
  assign N1078 = N14 & N15;
  assign N14 = ~addr_i[0];
  assign N15 = ~addr_i[1];
  assign N1079 = N1071 & N1075;
  assign N1080 = N1071 & N1076;
  assign N1081 = N1071 & N1077;
  assign N1082 = N1071 & N1078;
  assign N1083 = N1072 & N1075;
  assign N1084 = N1072 & N1076;
  assign N1085 = N1072 & N1077;
  assign N1086 = N1072 & N1078;
  assign N1087 = N1073 & N1075;
  assign N1088 = N1073 & N1076;
  assign N1089 = N1073 & N1077;
  assign N1090 = N1073 & N1078;
  assign N1091 = N1074 & N1075;
  assign N1092 = N1074 & N1076;
  assign N1093 = N1074 & N1077;
  assign N1094 = N1074 & N1078;
  assign N790 = N1055 & N1079;
  assign N789 = N1055 & N1080;
  assign N788 = N1055 & N1081;
  assign N787 = N1055 & N1082;
  assign N786 = N1055 & N1083;
  assign N785 = N1055 & N1084;
  assign N784 = N1055 & N1085;
  assign N783 = N1055 & N1086;
  assign N782 = N1055 & N1087;
  assign N781 = N1055 & N1088;
  assign N780 = N1055 & N1089;
  assign N779 = N1055 & N1090;
  assign N778 = N1055 & N1091;
  assign N777 = N1055 & N1092;
  assign N776 = N1055 & N1093;
  assign N775 = N1055 & N1094;
  assign N774 = N1056 & N1079;
  assign N773 = N1056 & N1080;
  assign N772 = N1056 & N1081;
  assign N771 = N1056 & N1082;
  assign N770 = N1056 & N1083;
  assign N769 = N1056 & N1084;
  assign N768 = N1056 & N1085;
  assign N767 = N1056 & N1086;
  assign N766 = N1056 & N1087;
  assign N765 = N1056 & N1088;
  assign N764 = N1056 & N1089;
  assign N763 = N1056 & N1090;
  assign N762 = N1056 & N1091;
  assign N761 = N1056 & N1092;
  assign N760 = N1056 & N1093;
  assign N759 = N1056 & N1094;
  assign N758 = N1057 & N1079;
  assign N757 = N1057 & N1080;
  assign N756 = N1057 & N1081;
  assign N755 = N1057 & N1082;
  assign N754 = N1057 & N1083;
  assign N753 = N1057 & N1084;
  assign N752 = N1057 & N1085;
  assign N751 = N1057 & N1086;
  assign N750 = N1057 & N1087;
  assign N749 = N1057 & N1088;
  assign N748 = N1057 & N1089;
  assign N747 = N1057 & N1090;
  assign N746 = N1057 & N1091;
  assign N745 = N1057 & N1092;
  assign N744 = N1057 & N1093;
  assign N743 = N1057 & N1094;
  assign N742 = N1058 & N1079;
  assign N741 = N1058 & N1080;
  assign N740 = N1058 & N1081;
  assign N739 = N1058 & N1082;
  assign N738 = N1058 & N1083;
  assign N737 = N1058 & N1084;
  assign N736 = N1058 & N1085;
  assign N735 = N1058 & N1086;
  assign N734 = N1058 & N1087;
  assign N733 = N1058 & N1088;
  assign N732 = N1058 & N1089;
  assign N731 = N1058 & N1090;
  assign N730 = N1058 & N1091;
  assign N729 = N1058 & N1092;
  assign N728 = N1058 & N1093;
  assign N727 = N1058 & N1094;
  assign N726 = N1059 & N1079;
  assign N725 = N1059 & N1080;
  assign N724 = N1059 & N1081;
  assign N723 = N1059 & N1082;
  assign N722 = N1059 & N1083;
  assign N721 = N1059 & N1084;
  assign N720 = N1059 & N1085;
  assign N719 = N1059 & N1086;
  assign N718 = N1059 & N1087;
  assign N717 = N1059 & N1088;
  assign N716 = N1059 & N1089;
  assign N715 = N1059 & N1090;
  assign N714 = N1059 & N1091;
  assign N713 = N1059 & N1092;
  assign N712 = N1059 & N1093;
  assign N711 = N1059 & N1094;
  assign N710 = N1060 & N1079;
  assign N709 = N1060 & N1080;
  assign N708 = N1060 & N1081;
  assign N707 = N1060 & N1082;
  assign N706 = N1060 & N1083;
  assign N705 = N1060 & N1084;
  assign N704 = N1060 & N1085;
  assign N703 = N1060 & N1086;
  assign N702 = N1060 & N1087;
  assign N701 = N1060 & N1088;
  assign N700 = N1060 & N1089;
  assign N699 = N1060 & N1090;
  assign N698 = N1060 & N1091;
  assign N697 = N1060 & N1092;
  assign N696 = N1060 & N1093;
  assign N695 = N1060 & N1094;
  assign N694 = N1061 & N1079;
  assign N693 = N1061 & N1080;
  assign N692 = N1061 & N1081;
  assign N691 = N1061 & N1082;
  assign N690 = N1061 & N1083;
  assign N689 = N1061 & N1084;
  assign N688 = N1061 & N1085;
  assign N687 = N1061 & N1086;
  assign N686 = N1061 & N1087;
  assign N685 = N1061 & N1088;
  assign N684 = N1061 & N1089;
  assign N683 = N1061 & N1090;
  assign N682 = N1061 & N1091;
  assign N681 = N1061 & N1092;
  assign N680 = N1061 & N1093;
  assign N679 = N1061 & N1094;
  assign N678 = N1062 & N1079;
  assign N677 = N1062 & N1080;
  assign N676 = N1062 & N1081;
  assign N675 = N1062 & N1082;
  assign N674 = N1062 & N1083;
  assign N673 = N1062 & N1084;
  assign N672 = N1062 & N1085;
  assign N671 = N1062 & N1086;
  assign N670 = N1062 & N1087;
  assign N669 = N1062 & N1088;
  assign N668 = N1062 & N1089;
  assign N667 = N1062 & N1090;
  assign N666 = N1062 & N1091;
  assign N665 = N1062 & N1092;
  assign N664 = N1062 & N1093;
  assign N663 = N1062 & N1094;
  assign N662 = N1063 & N1079;
  assign N661 = N1063 & N1080;
  assign N660 = N1063 & N1081;
  assign N659 = N1063 & N1082;
  assign N658 = N1063 & N1083;
  assign N657 = N1063 & N1084;
  assign N656 = N1063 & N1085;
  assign N655 = N1063 & N1086;
  assign N654 = N1063 & N1087;
  assign N653 = N1063 & N1088;
  assign N652 = N1063 & N1089;
  assign N651 = N1063 & N1090;
  assign N650 = N1063 & N1091;
  assign N649 = N1063 & N1092;
  assign N648 = N1063 & N1093;
  assign N647 = N1063 & N1094;
  assign N646 = N1064 & N1079;
  assign N645 = N1064 & N1080;
  assign N644 = N1064 & N1081;
  assign N643 = N1064 & N1082;
  assign N642 = N1064 & N1083;
  assign N641 = N1064 & N1084;
  assign N640 = N1064 & N1085;
  assign N639 = N1064 & N1086;
  assign N638 = N1064 & N1087;
  assign N637 = N1064 & N1088;
  assign N636 = N1064 & N1089;
  assign N635 = N1064 & N1090;
  assign N634 = N1064 & N1091;
  assign N633 = N1064 & N1092;
  assign N632 = N1064 & N1093;
  assign N631 = N1064 & N1094;
  assign N630 = N1065 & N1079;
  assign N629 = N1065 & N1080;
  assign N628 = N1065 & N1081;
  assign N627 = N1065 & N1082;
  assign N626 = N1065 & N1083;
  assign N625 = N1065 & N1084;
  assign N624 = N1065 & N1085;
  assign N623 = N1065 & N1086;
  assign N622 = N1065 & N1087;
  assign N621 = N1065 & N1088;
  assign N620 = N1065 & N1089;
  assign N619 = N1065 & N1090;
  assign N618 = N1065 & N1091;
  assign N617 = N1065 & N1092;
  assign N616 = N1065 & N1093;
  assign N615 = N1065 & N1094;
  assign N614 = N1066 & N1079;
  assign N613 = N1066 & N1080;
  assign N612 = N1066 & N1081;
  assign N611 = N1066 & N1082;
  assign N610 = N1066 & N1083;
  assign N609 = N1066 & N1084;
  assign N608 = N1066 & N1085;
  assign N607 = N1066 & N1086;
  assign N606 = N1066 & N1087;
  assign N605 = N1066 & N1088;
  assign N604 = N1066 & N1089;
  assign N603 = N1066 & N1090;
  assign N602 = N1066 & N1091;
  assign N601 = N1066 & N1092;
  assign N600 = N1066 & N1093;
  assign N599 = N1066 & N1094;
  assign N598 = N1067 & N1079;
  assign N597 = N1067 & N1080;
  assign N596 = N1067 & N1081;
  assign N595 = N1067 & N1082;
  assign N594 = N1067 & N1083;
  assign N593 = N1067 & N1084;
  assign N592 = N1067 & N1085;
  assign N591 = N1067 & N1086;
  assign N590 = N1067 & N1087;
  assign N589 = N1067 & N1088;
  assign N588 = N1067 & N1089;
  assign N587 = N1067 & N1090;
  assign N586 = N1067 & N1091;
  assign N585 = N1067 & N1092;
  assign N584 = N1067 & N1093;
  assign N583 = N1067 & N1094;
  assign N582 = N1068 & N1079;
  assign N581 = N1068 & N1080;
  assign N580 = N1068 & N1081;
  assign N579 = N1068 & N1082;
  assign N578 = N1068 & N1083;
  assign N577 = N1068 & N1084;
  assign N576 = N1068 & N1085;
  assign N575 = N1068 & N1086;
  assign N574 = N1068 & N1087;
  assign N573 = N1068 & N1088;
  assign N572 = N1068 & N1089;
  assign N571 = N1068 & N1090;
  assign N570 = N1068 & N1091;
  assign N569 = N1068 & N1092;
  assign N568 = N1068 & N1093;
  assign N567 = N1068 & N1094;
  assign N566 = N1069 & N1079;
  assign N565 = N1069 & N1080;
  assign N564 = N1069 & N1081;
  assign N563 = N1069 & N1082;
  assign N562 = N1069 & N1083;
  assign N561 = N1069 & N1084;
  assign N560 = N1069 & N1085;
  assign N559 = N1069 & N1086;
  assign N558 = N1069 & N1087;
  assign N557 = N1069 & N1088;
  assign N556 = N1069 & N1089;
  assign N555 = N1069 & N1090;
  assign N554 = N1069 & N1091;
  assign N553 = N1069 & N1092;
  assign N552 = N1069 & N1093;
  assign N551 = N1069 & N1094;
  assign N550 = N1070 & N1079;
  assign N549 = N1070 & N1080;
  assign N548 = N1070 & N1081;
  assign N547 = N1070 & N1082;
  assign N546 = N1070 & N1083;
  assign N545 = N1070 & N1084;
  assign N544 = N1070 & N1085;
  assign N543 = N1070 & N1086;
  assign N542 = N1070 & N1087;
  assign N541 = N1070 & N1088;
  assign N540 = N1070 & N1089;
  assign N539 = N1070 & N1090;
  assign N538 = N1070 & N1091;
  assign N537 = N1070 & N1092;
  assign N536 = N1070 & N1093;
  assign N535 = N1070 & N1094;
  assign { N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791 } = (N16)? { N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             (N534)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = N533;
  assign read_en = v_i & N1095;
  assign N1095 = ~w_i;
  assign N17 = ~addr_r[0];
  assign N18 = ~addr_r[1];
  assign N19 = N17 & N18;
  assign N20 = N17 & addr_r[1];
  assign N21 = addr_r[0] & N18;
  assign N22 = addr_r[0] & addr_r[1];
  assign N23 = ~addr_r[2];
  assign N24 = N19 & N23;
  assign N25 = N19 & addr_r[2];
  assign N26 = N21 & N23;
  assign N27 = N21 & addr_r[2];
  assign N28 = N20 & N23;
  assign N29 = N20 & addr_r[2];
  assign N30 = N22 & N23;
  assign N31 = N22 & addr_r[2];
  assign N32 = ~addr_r[3];
  assign N33 = N24 & N32;
  assign N34 = N24 & addr_r[3];
  assign N35 = N26 & N32;
  assign N36 = N26 & addr_r[3];
  assign N37 = N28 & N32;
  assign N38 = N28 & addr_r[3];
  assign N39 = N30 & N32;
  assign N40 = N30 & addr_r[3];
  assign N41 = N25 & N32;
  assign N42 = N25 & addr_r[3];
  assign N43 = N27 & N32;
  assign N44 = N27 & addr_r[3];
  assign N45 = N29 & N32;
  assign N46 = N29 & addr_r[3];
  assign N47 = N31 & N32;
  assign N48 = N31 & addr_r[3];
  assign N49 = ~addr_r[4];
  assign N50 = N33 & N49;
  assign N51 = N33 & addr_r[4];
  assign N52 = N35 & N49;
  assign N53 = N35 & addr_r[4];
  assign N54 = N37 & N49;
  assign N55 = N37 & addr_r[4];
  assign N56 = N39 & N49;
  assign N57 = N39 & addr_r[4];
  assign N58 = N41 & N49;
  assign N59 = N41 & addr_r[4];
  assign N60 = N43 & N49;
  assign N61 = N43 & addr_r[4];
  assign N62 = N45 & N49;
  assign N63 = N45 & addr_r[4];
  assign N64 = N47 & N49;
  assign N65 = N47 & addr_r[4];
  assign N66 = N34 & N49;
  assign N67 = N34 & addr_r[4];
  assign N68 = N36 & N49;
  assign N69 = N36 & addr_r[4];
  assign N70 = N38 & N49;
  assign N71 = N38 & addr_r[4];
  assign N72 = N40 & N49;
  assign N73 = N40 & addr_r[4];
  assign N74 = N42 & N49;
  assign N75 = N42 & addr_r[4];
  assign N76 = N44 & N49;
  assign N77 = N44 & addr_r[4];
  assign N78 = N46 & N49;
  assign N79 = N46 & addr_r[4];
  assign N80 = N48 & N49;
  assign N81 = N48 & addr_r[4];
  assign N82 = ~addr_r[5];
  assign N83 = N50 & N82;
  assign N84 = N50 & addr_r[5];
  assign N85 = N52 & N82;
  assign N86 = N52 & addr_r[5];
  assign N87 = N54 & N82;
  assign N88 = N54 & addr_r[5];
  assign N89 = N56 & N82;
  assign N90 = N56 & addr_r[5];
  assign N91 = N58 & N82;
  assign N92 = N58 & addr_r[5];
  assign N93 = N60 & N82;
  assign N94 = N60 & addr_r[5];
  assign N95 = N62 & N82;
  assign N96 = N62 & addr_r[5];
  assign N97 = N64 & N82;
  assign N98 = N64 & addr_r[5];
  assign N99 = N66 & N82;
  assign N100 = N66 & addr_r[5];
  assign N101 = N68 & N82;
  assign N102 = N68 & addr_r[5];
  assign N103 = N70 & N82;
  assign N104 = N70 & addr_r[5];
  assign N105 = N72 & N82;
  assign N106 = N72 & addr_r[5];
  assign N107 = N74 & N82;
  assign N108 = N74 & addr_r[5];
  assign N109 = N76 & N82;
  assign N110 = N76 & addr_r[5];
  assign N111 = N78 & N82;
  assign N112 = N78 & addr_r[5];
  assign N113 = N80 & N82;
  assign N114 = N80 & addr_r[5];
  assign N115 = N51 & N82;
  assign N116 = N51 & addr_r[5];
  assign N117 = N53 & N82;
  assign N118 = N53 & addr_r[5];
  assign N119 = N55 & N82;
  assign N120 = N55 & addr_r[5];
  assign N121 = N57 & N82;
  assign N122 = N57 & addr_r[5];
  assign N123 = N59 & N82;
  assign N124 = N59 & addr_r[5];
  assign N125 = N61 & N82;
  assign N126 = N61 & addr_r[5];
  assign N127 = N63 & N82;
  assign N128 = N63 & addr_r[5];
  assign N129 = N65 & N82;
  assign N130 = N65 & addr_r[5];
  assign N131 = N67 & N82;
  assign N132 = N67 & addr_r[5];
  assign N133 = N69 & N82;
  assign N134 = N69 & addr_r[5];
  assign N135 = N71 & N82;
  assign N136 = N71 & addr_r[5];
  assign N137 = N73 & N82;
  assign N138 = N73 & addr_r[5];
  assign N139 = N75 & N82;
  assign N140 = N75 & addr_r[5];
  assign N141 = N77 & N82;
  assign N142 = N77 & addr_r[5];
  assign N143 = N79 & N82;
  assign N144 = N79 & addr_r[5];
  assign N145 = N81 & N82;
  assign N146 = N81 & addr_r[5];
  assign N147 = ~addr_r[6];
  assign N148 = N83 & N147;
  assign N149 = N83 & addr_r[6];
  assign N150 = N85 & N147;
  assign N151 = N85 & addr_r[6];
  assign N152 = N87 & N147;
  assign N153 = N87 & addr_r[6];
  assign N154 = N89 & N147;
  assign N155 = N89 & addr_r[6];
  assign N156 = N91 & N147;
  assign N157 = N91 & addr_r[6];
  assign N158 = N93 & N147;
  assign N159 = N93 & addr_r[6];
  assign N160 = N95 & N147;
  assign N161 = N95 & addr_r[6];
  assign N162 = N97 & N147;
  assign N163 = N97 & addr_r[6];
  assign N164 = N99 & N147;
  assign N165 = N99 & addr_r[6];
  assign N166 = N101 & N147;
  assign N167 = N101 & addr_r[6];
  assign N168 = N103 & N147;
  assign N169 = N103 & addr_r[6];
  assign N170 = N105 & N147;
  assign N171 = N105 & addr_r[6];
  assign N172 = N107 & N147;
  assign N173 = N107 & addr_r[6];
  assign N174 = N109 & N147;
  assign N175 = N109 & addr_r[6];
  assign N176 = N111 & N147;
  assign N177 = N111 & addr_r[6];
  assign N178 = N113 & N147;
  assign N179 = N113 & addr_r[6];
  assign N180 = N115 & N147;
  assign N181 = N115 & addr_r[6];
  assign N182 = N117 & N147;
  assign N183 = N117 & addr_r[6];
  assign N184 = N119 & N147;
  assign N185 = N119 & addr_r[6];
  assign N186 = N121 & N147;
  assign N187 = N121 & addr_r[6];
  assign N188 = N123 & N147;
  assign N189 = N123 & addr_r[6];
  assign N190 = N125 & N147;
  assign N191 = N125 & addr_r[6];
  assign N192 = N127 & N147;
  assign N193 = N127 & addr_r[6];
  assign N194 = N129 & N147;
  assign N195 = N129 & addr_r[6];
  assign N196 = N131 & N147;
  assign N197 = N131 & addr_r[6];
  assign N198 = N133 & N147;
  assign N199 = N133 & addr_r[6];
  assign N200 = N135 & N147;
  assign N201 = N135 & addr_r[6];
  assign N202 = N137 & N147;
  assign N203 = N137 & addr_r[6];
  assign N204 = N139 & N147;
  assign N205 = N139 & addr_r[6];
  assign N206 = N141 & N147;
  assign N207 = N141 & addr_r[6];
  assign N208 = N143 & N147;
  assign N209 = N143 & addr_r[6];
  assign N210 = N145 & N147;
  assign N211 = N145 & addr_r[6];
  assign N212 = N84 & N147;
  assign N213 = N84 & addr_r[6];
  assign N214 = N86 & N147;
  assign N215 = N86 & addr_r[6];
  assign N216 = N88 & N147;
  assign N217 = N88 & addr_r[6];
  assign N218 = N90 & N147;
  assign N219 = N90 & addr_r[6];
  assign N220 = N92 & N147;
  assign N221 = N92 & addr_r[6];
  assign N222 = N94 & N147;
  assign N223 = N94 & addr_r[6];
  assign N224 = N96 & N147;
  assign N225 = N96 & addr_r[6];
  assign N226 = N98 & N147;
  assign N227 = N98 & addr_r[6];
  assign N228 = N100 & N147;
  assign N229 = N100 & addr_r[6];
  assign N230 = N102 & N147;
  assign N231 = N102 & addr_r[6];
  assign N232 = N104 & N147;
  assign N233 = N104 & addr_r[6];
  assign N234 = N106 & N147;
  assign N235 = N106 & addr_r[6];
  assign N236 = N108 & N147;
  assign N237 = N108 & addr_r[6];
  assign N238 = N110 & N147;
  assign N239 = N110 & addr_r[6];
  assign N240 = N112 & N147;
  assign N241 = N112 & addr_r[6];
  assign N242 = N114 & N147;
  assign N243 = N114 & addr_r[6];
  assign N244 = N116 & N147;
  assign N245 = N116 & addr_r[6];
  assign N246 = N118 & N147;
  assign N247 = N118 & addr_r[6];
  assign N248 = N120 & N147;
  assign N249 = N120 & addr_r[6];
  assign N250 = N122 & N147;
  assign N251 = N122 & addr_r[6];
  assign N252 = N124 & N147;
  assign N253 = N124 & addr_r[6];
  assign N254 = N126 & N147;
  assign N255 = N126 & addr_r[6];
  assign N256 = N128 & N147;
  assign N257 = N128 & addr_r[6];
  assign N258 = N130 & N147;
  assign N259 = N130 & addr_r[6];
  assign N260 = N132 & N147;
  assign N261 = N132 & addr_r[6];
  assign N262 = N134 & N147;
  assign N263 = N134 & addr_r[6];
  assign N264 = N136 & N147;
  assign N265 = N136 & addr_r[6];
  assign N266 = N138 & N147;
  assign N267 = N138 & addr_r[6];
  assign N268 = N140 & N147;
  assign N269 = N140 & addr_r[6];
  assign N270 = N142 & N147;
  assign N271 = N142 & addr_r[6];
  assign N272 = N144 & N147;
  assign N273 = N144 & addr_r[6];
  assign N274 = N146 & N147;
  assign N275 = N146 & addr_r[6];
  assign N276 = ~addr_r[7];
  assign N277 = N148 & N276;
  assign N278 = N148 & addr_r[7];
  assign N279 = N150 & N276;
  assign N280 = N150 & addr_r[7];
  assign N281 = N152 & N276;
  assign N282 = N152 & addr_r[7];
  assign N283 = N154 & N276;
  assign N284 = N154 & addr_r[7];
  assign N285 = N156 & N276;
  assign N286 = N156 & addr_r[7];
  assign N287 = N158 & N276;
  assign N288 = N158 & addr_r[7];
  assign N289 = N160 & N276;
  assign N290 = N160 & addr_r[7];
  assign N291 = N162 & N276;
  assign N292 = N162 & addr_r[7];
  assign N293 = N164 & N276;
  assign N294 = N164 & addr_r[7];
  assign N295 = N166 & N276;
  assign N296 = N166 & addr_r[7];
  assign N297 = N168 & N276;
  assign N298 = N168 & addr_r[7];
  assign N299 = N170 & N276;
  assign N300 = N170 & addr_r[7];
  assign N301 = N172 & N276;
  assign N302 = N172 & addr_r[7];
  assign N303 = N174 & N276;
  assign N304 = N174 & addr_r[7];
  assign N305 = N176 & N276;
  assign N306 = N176 & addr_r[7];
  assign N307 = N178 & N276;
  assign N308 = N178 & addr_r[7];
  assign N309 = N180 & N276;
  assign N310 = N180 & addr_r[7];
  assign N311 = N182 & N276;
  assign N312 = N182 & addr_r[7];
  assign N313 = N184 & N276;
  assign N314 = N184 & addr_r[7];
  assign N315 = N186 & N276;
  assign N316 = N186 & addr_r[7];
  assign N317 = N188 & N276;
  assign N318 = N188 & addr_r[7];
  assign N319 = N190 & N276;
  assign N320 = N190 & addr_r[7];
  assign N321 = N192 & N276;
  assign N322 = N192 & addr_r[7];
  assign N323 = N194 & N276;
  assign N324 = N194 & addr_r[7];
  assign N325 = N196 & N276;
  assign N326 = N196 & addr_r[7];
  assign N327 = N198 & N276;
  assign N328 = N198 & addr_r[7];
  assign N329 = N200 & N276;
  assign N330 = N200 & addr_r[7];
  assign N331 = N202 & N276;
  assign N332 = N202 & addr_r[7];
  assign N333 = N204 & N276;
  assign N334 = N204 & addr_r[7];
  assign N335 = N206 & N276;
  assign N336 = N206 & addr_r[7];
  assign N337 = N208 & N276;
  assign N338 = N208 & addr_r[7];
  assign N339 = N210 & N276;
  assign N340 = N210 & addr_r[7];
  assign N341 = N212 & N276;
  assign N342 = N212 & addr_r[7];
  assign N343 = N214 & N276;
  assign N344 = N214 & addr_r[7];
  assign N345 = N216 & N276;
  assign N346 = N216 & addr_r[7];
  assign N347 = N218 & N276;
  assign N348 = N218 & addr_r[7];
  assign N349 = N220 & N276;
  assign N350 = N220 & addr_r[7];
  assign N351 = N222 & N276;
  assign N352 = N222 & addr_r[7];
  assign N353 = N224 & N276;
  assign N354 = N224 & addr_r[7];
  assign N355 = N226 & N276;
  assign N356 = N226 & addr_r[7];
  assign N357 = N228 & N276;
  assign N358 = N228 & addr_r[7];
  assign N359 = N230 & N276;
  assign N360 = N230 & addr_r[7];
  assign N361 = N232 & N276;
  assign N362 = N232 & addr_r[7];
  assign N363 = N234 & N276;
  assign N364 = N234 & addr_r[7];
  assign N365 = N236 & N276;
  assign N366 = N236 & addr_r[7];
  assign N367 = N238 & N276;
  assign N368 = N238 & addr_r[7];
  assign N369 = N240 & N276;
  assign N370 = N240 & addr_r[7];
  assign N371 = N242 & N276;
  assign N372 = N242 & addr_r[7];
  assign N373 = N244 & N276;
  assign N374 = N244 & addr_r[7];
  assign N375 = N246 & N276;
  assign N376 = N246 & addr_r[7];
  assign N377 = N248 & N276;
  assign N378 = N248 & addr_r[7];
  assign N379 = N250 & N276;
  assign N380 = N250 & addr_r[7];
  assign N381 = N252 & N276;
  assign N382 = N252 & addr_r[7];
  assign N383 = N254 & N276;
  assign N384 = N254 & addr_r[7];
  assign N385 = N256 & N276;
  assign N386 = N256 & addr_r[7];
  assign N387 = N258 & N276;
  assign N388 = N258 & addr_r[7];
  assign N389 = N260 & N276;
  assign N390 = N260 & addr_r[7];
  assign N391 = N262 & N276;
  assign N392 = N262 & addr_r[7];
  assign N393 = N264 & N276;
  assign N394 = N264 & addr_r[7];
  assign N395 = N266 & N276;
  assign N396 = N266 & addr_r[7];
  assign N397 = N268 & N276;
  assign N398 = N268 & addr_r[7];
  assign N399 = N270 & N276;
  assign N400 = N270 & addr_r[7];
  assign N401 = N272 & N276;
  assign N402 = N272 & addr_r[7];
  assign N403 = N274 & N276;
  assign N404 = N274 & addr_r[7];
  assign N405 = N149 & N276;
  assign N406 = N149 & addr_r[7];
  assign N407 = N151 & N276;
  assign N408 = N151 & addr_r[7];
  assign N409 = N153 & N276;
  assign N410 = N153 & addr_r[7];
  assign N411 = N155 & N276;
  assign N412 = N155 & addr_r[7];
  assign N413 = N157 & N276;
  assign N414 = N157 & addr_r[7];
  assign N415 = N159 & N276;
  assign N416 = N159 & addr_r[7];
  assign N417 = N161 & N276;
  assign N418 = N161 & addr_r[7];
  assign N419 = N163 & N276;
  assign N420 = N163 & addr_r[7];
  assign N421 = N165 & N276;
  assign N422 = N165 & addr_r[7];
  assign N423 = N167 & N276;
  assign N424 = N167 & addr_r[7];
  assign N425 = N169 & N276;
  assign N426 = N169 & addr_r[7];
  assign N427 = N171 & N276;
  assign N428 = N171 & addr_r[7];
  assign N429 = N173 & N276;
  assign N430 = N173 & addr_r[7];
  assign N431 = N175 & N276;
  assign N432 = N175 & addr_r[7];
  assign N433 = N177 & N276;
  assign N434 = N177 & addr_r[7];
  assign N435 = N179 & N276;
  assign N436 = N179 & addr_r[7];
  assign N437 = N181 & N276;
  assign N438 = N181 & addr_r[7];
  assign N439 = N183 & N276;
  assign N440 = N183 & addr_r[7];
  assign N441 = N185 & N276;
  assign N442 = N185 & addr_r[7];
  assign N443 = N187 & N276;
  assign N444 = N187 & addr_r[7];
  assign N445 = N189 & N276;
  assign N446 = N189 & addr_r[7];
  assign N447 = N191 & N276;
  assign N448 = N191 & addr_r[7];
  assign N449 = N193 & N276;
  assign N450 = N193 & addr_r[7];
  assign N451 = N195 & N276;
  assign N452 = N195 & addr_r[7];
  assign N453 = N197 & N276;
  assign N454 = N197 & addr_r[7];
  assign N455 = N199 & N276;
  assign N456 = N199 & addr_r[7];
  assign N457 = N201 & N276;
  assign N458 = N201 & addr_r[7];
  assign N459 = N203 & N276;
  assign N460 = N203 & addr_r[7];
  assign N461 = N205 & N276;
  assign N462 = N205 & addr_r[7];
  assign N463 = N207 & N276;
  assign N464 = N207 & addr_r[7];
  assign N465 = N209 & N276;
  assign N466 = N209 & addr_r[7];
  assign N467 = N211 & N276;
  assign N468 = N211 & addr_r[7];
  assign N469 = N213 & N276;
  assign N470 = N213 & addr_r[7];
  assign N471 = N215 & N276;
  assign N472 = N215 & addr_r[7];
  assign N473 = N217 & N276;
  assign N474 = N217 & addr_r[7];
  assign N475 = N219 & N276;
  assign N476 = N219 & addr_r[7];
  assign N477 = N221 & N276;
  assign N478 = N221 & addr_r[7];
  assign N479 = N223 & N276;
  assign N480 = N223 & addr_r[7];
  assign N481 = N225 & N276;
  assign N482 = N225 & addr_r[7];
  assign N483 = N227 & N276;
  assign N484 = N227 & addr_r[7];
  assign N485 = N229 & N276;
  assign N486 = N229 & addr_r[7];
  assign N487 = N231 & N276;
  assign N488 = N231 & addr_r[7];
  assign N489 = N233 & N276;
  assign N490 = N233 & addr_r[7];
  assign N491 = N235 & N276;
  assign N492 = N235 & addr_r[7];
  assign N493 = N237 & N276;
  assign N494 = N237 & addr_r[7];
  assign N495 = N239 & N276;
  assign N496 = N239 & addr_r[7];
  assign N497 = N241 & N276;
  assign N498 = N241 & addr_r[7];
  assign N499 = N243 & N276;
  assign N500 = N243 & addr_r[7];
  assign N501 = N245 & N276;
  assign N502 = N245 & addr_r[7];
  assign N503 = N247 & N276;
  assign N504 = N247 & addr_r[7];
  assign N505 = N249 & N276;
  assign N506 = N249 & addr_r[7];
  assign N507 = N251 & N276;
  assign N508 = N251 & addr_r[7];
  assign N509 = N253 & N276;
  assign N510 = N253 & addr_r[7];
  assign N511 = N255 & N276;
  assign N512 = N255 & addr_r[7];
  assign N513 = N257 & N276;
  assign N514 = N257 & addr_r[7];
  assign N515 = N259 & N276;
  assign N516 = N259 & addr_r[7];
  assign N517 = N261 & N276;
  assign N518 = N261 & addr_r[7];
  assign N519 = N263 & N276;
  assign N520 = N263 & addr_r[7];
  assign N521 = N265 & N276;
  assign N522 = N265 & addr_r[7];
  assign N523 = N267 & N276;
  assign N524 = N267 & addr_r[7];
  assign N525 = N269 & N276;
  assign N526 = N269 & addr_r[7];
  assign N527 = N271 & N276;
  assign N528 = N271 & addr_r[7];
  assign N529 = N273 & N276;
  assign N530 = N273 & addr_r[7];
  assign N531 = N275 & N276;
  assign N532 = N275 & addr_r[7];
  assign N533 = v_i & w_i;
  assign N534 = ~N533;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { addr_r[7:0] } <= { addr_i[7:0] };
    end 
    if(N1046) begin
      { mem[2047:2040] } <= { data_i[7:0] };
    end 
    if(N1045) begin
      { mem[2039:2032] } <= { data_i[7:0] };
    end 
    if(N1044) begin
      { mem[2031:2024] } <= { data_i[7:0] };
    end 
    if(N1043) begin
      { mem[2023:2016] } <= { data_i[7:0] };
    end 
    if(N1042) begin
      { mem[2015:2008] } <= { data_i[7:0] };
    end 
    if(N1041) begin
      { mem[2007:2000] } <= { data_i[7:0] };
    end 
    if(N1040) begin
      { mem[1999:1992] } <= { data_i[7:0] };
    end 
    if(N1039) begin
      { mem[1991:1984] } <= { data_i[7:0] };
    end 
    if(N1038) begin
      { mem[1983:1976] } <= { data_i[7:0] };
    end 
    if(N1037) begin
      { mem[1975:1968] } <= { data_i[7:0] };
    end 
    if(N1036) begin
      { mem[1967:1960] } <= { data_i[7:0] };
    end 
    if(N1035) begin
      { mem[1959:1952] } <= { data_i[7:0] };
    end 
    if(N1034) begin
      { mem[1951:1944] } <= { data_i[7:0] };
    end 
    if(N1033) begin
      { mem[1943:1936] } <= { data_i[7:0] };
    end 
    if(N1032) begin
      { mem[1935:1928] } <= { data_i[7:0] };
    end 
    if(N1031) begin
      { mem[1927:1920] } <= { data_i[7:0] };
    end 
    if(N1030) begin
      { mem[1919:1912] } <= { data_i[7:0] };
    end 
    if(N1029) begin
      { mem[1911:1904] } <= { data_i[7:0] };
    end 
    if(N1028) begin
      { mem[1903:1896] } <= { data_i[7:0] };
    end 
    if(N1027) begin
      { mem[1895:1888] } <= { data_i[7:0] };
    end 
    if(N1026) begin
      { mem[1887:1880] } <= { data_i[7:0] };
    end 
    if(N1025) begin
      { mem[1879:1872] } <= { data_i[7:0] };
    end 
    if(N1024) begin
      { mem[1871:1864] } <= { data_i[7:0] };
    end 
    if(N1023) begin
      { mem[1863:1856] } <= { data_i[7:0] };
    end 
    if(N1022) begin
      { mem[1855:1848] } <= { data_i[7:0] };
    end 
    if(N1021) begin
      { mem[1847:1840] } <= { data_i[7:0] };
    end 
    if(N1020) begin
      { mem[1839:1832] } <= { data_i[7:0] };
    end 
    if(N1019) begin
      { mem[1831:1824] } <= { data_i[7:0] };
    end 
    if(N1018) begin
      { mem[1823:1816] } <= { data_i[7:0] };
    end 
    if(N1017) begin
      { mem[1815:1808] } <= { data_i[7:0] };
    end 
    if(N1016) begin
      { mem[1807:1800] } <= { data_i[7:0] };
    end 
    if(N1015) begin
      { mem[1799:1792] } <= { data_i[7:0] };
    end 
    if(N1014) begin
      { mem[1791:1784] } <= { data_i[7:0] };
    end 
    if(N1013) begin
      { mem[1783:1776] } <= { data_i[7:0] };
    end 
    if(N1012) begin
      { mem[1775:1768] } <= { data_i[7:0] };
    end 
    if(N1011) begin
      { mem[1767:1760] } <= { data_i[7:0] };
    end 
    if(N1010) begin
      { mem[1759:1752] } <= { data_i[7:0] };
    end 
    if(N1009) begin
      { mem[1751:1744] } <= { data_i[7:0] };
    end 
    if(N1008) begin
      { mem[1743:1736] } <= { data_i[7:0] };
    end 
    if(N1007) begin
      { mem[1735:1728] } <= { data_i[7:0] };
    end 
    if(N1006) begin
      { mem[1727:1720] } <= { data_i[7:0] };
    end 
    if(N1005) begin
      { mem[1719:1712] } <= { data_i[7:0] };
    end 
    if(N1004) begin
      { mem[1711:1704] } <= { data_i[7:0] };
    end 
    if(N1003) begin
      { mem[1703:1696] } <= { data_i[7:0] };
    end 
    if(N1002) begin
      { mem[1695:1688] } <= { data_i[7:0] };
    end 
    if(N1001) begin
      { mem[1687:1680] } <= { data_i[7:0] };
    end 
    if(N1000) begin
      { mem[1679:1672] } <= { data_i[7:0] };
    end 
    if(N999) begin
      { mem[1671:1664] } <= { data_i[7:0] };
    end 
    if(N998) begin
      { mem[1663:1656] } <= { data_i[7:0] };
    end 
    if(N997) begin
      { mem[1655:1648] } <= { data_i[7:0] };
    end 
    if(N996) begin
      { mem[1647:1640] } <= { data_i[7:0] };
    end 
    if(N995) begin
      { mem[1639:1632] } <= { data_i[7:0] };
    end 
    if(N994) begin
      { mem[1631:1624] } <= { data_i[7:0] };
    end 
    if(N993) begin
      { mem[1623:1616] } <= { data_i[7:0] };
    end 
    if(N992) begin
      { mem[1615:1608] } <= { data_i[7:0] };
    end 
    if(N991) begin
      { mem[1607:1600] } <= { data_i[7:0] };
    end 
    if(N990) begin
      { mem[1599:1592] } <= { data_i[7:0] };
    end 
    if(N989) begin
      { mem[1591:1584] } <= { data_i[7:0] };
    end 
    if(N988) begin
      { mem[1583:1576] } <= { data_i[7:0] };
    end 
    if(N987) begin
      { mem[1575:1568] } <= { data_i[7:0] };
    end 
    if(N986) begin
      { mem[1567:1560] } <= { data_i[7:0] };
    end 
    if(N985) begin
      { mem[1559:1552] } <= { data_i[7:0] };
    end 
    if(N984) begin
      { mem[1551:1544] } <= { data_i[7:0] };
    end 
    if(N983) begin
      { mem[1543:1536] } <= { data_i[7:0] };
    end 
    if(N982) begin
      { mem[1535:1528] } <= { data_i[7:0] };
    end 
    if(N981) begin
      { mem[1527:1520] } <= { data_i[7:0] };
    end 
    if(N980) begin
      { mem[1519:1512] } <= { data_i[7:0] };
    end 
    if(N979) begin
      { mem[1511:1504] } <= { data_i[7:0] };
    end 
    if(N978) begin
      { mem[1503:1496] } <= { data_i[7:0] };
    end 
    if(N977) begin
      { mem[1495:1488] } <= { data_i[7:0] };
    end 
    if(N976) begin
      { mem[1487:1480] } <= { data_i[7:0] };
    end 
    if(N975) begin
      { mem[1479:1472] } <= { data_i[7:0] };
    end 
    if(N974) begin
      { mem[1471:1464] } <= { data_i[7:0] };
    end 
    if(N973) begin
      { mem[1463:1456] } <= { data_i[7:0] };
    end 
    if(N972) begin
      { mem[1455:1448] } <= { data_i[7:0] };
    end 
    if(N971) begin
      { mem[1447:1440] } <= { data_i[7:0] };
    end 
    if(N970) begin
      { mem[1439:1432] } <= { data_i[7:0] };
    end 
    if(N969) begin
      { mem[1431:1424] } <= { data_i[7:0] };
    end 
    if(N968) begin
      { mem[1423:1416] } <= { data_i[7:0] };
    end 
    if(N967) begin
      { mem[1415:1408] } <= { data_i[7:0] };
    end 
    if(N966) begin
      { mem[1407:1400] } <= { data_i[7:0] };
    end 
    if(N965) begin
      { mem[1399:1392] } <= { data_i[7:0] };
    end 
    if(N964) begin
      { mem[1391:1384] } <= { data_i[7:0] };
    end 
    if(N963) begin
      { mem[1383:1376] } <= { data_i[7:0] };
    end 
    if(N962) begin
      { mem[1375:1368] } <= { data_i[7:0] };
    end 
    if(N961) begin
      { mem[1367:1360] } <= { data_i[7:0] };
    end 
    if(N960) begin
      { mem[1359:1352] } <= { data_i[7:0] };
    end 
    if(N959) begin
      { mem[1351:1344] } <= { data_i[7:0] };
    end 
    if(N958) begin
      { mem[1343:1336] } <= { data_i[7:0] };
    end 
    if(N957) begin
      { mem[1335:1328] } <= { data_i[7:0] };
    end 
    if(N956) begin
      { mem[1327:1320] } <= { data_i[7:0] };
    end 
    if(N955) begin
      { mem[1319:1312] } <= { data_i[7:0] };
    end 
    if(N954) begin
      { mem[1311:1304] } <= { data_i[7:0] };
    end 
    if(N953) begin
      { mem[1303:1296] } <= { data_i[7:0] };
    end 
    if(N952) begin
      { mem[1295:1288] } <= { data_i[7:0] };
    end 
    if(N951) begin
      { mem[1287:1280] } <= { data_i[7:0] };
    end 
    if(N950) begin
      { mem[1279:1272] } <= { data_i[7:0] };
    end 
    if(N949) begin
      { mem[1271:1264] } <= { data_i[7:0] };
    end 
    if(N948) begin
      { mem[1263:1256] } <= { data_i[7:0] };
    end 
    if(N947) begin
      { mem[1255:1248] } <= { data_i[7:0] };
    end 
    if(N946) begin
      { mem[1247:1240] } <= { data_i[7:0] };
    end 
    if(N945) begin
      { mem[1239:1232] } <= { data_i[7:0] };
    end 
    if(N944) begin
      { mem[1231:1224] } <= { data_i[7:0] };
    end 
    if(N943) begin
      { mem[1223:1216] } <= { data_i[7:0] };
    end 
    if(N942) begin
      { mem[1215:1208] } <= { data_i[7:0] };
    end 
    if(N941) begin
      { mem[1207:1200] } <= { data_i[7:0] };
    end 
    if(N940) begin
      { mem[1199:1192] } <= { data_i[7:0] };
    end 
    if(N939) begin
      { mem[1191:1184] } <= { data_i[7:0] };
    end 
    if(N938) begin
      { mem[1183:1176] } <= { data_i[7:0] };
    end 
    if(N937) begin
      { mem[1175:1168] } <= { data_i[7:0] };
    end 
    if(N936) begin
      { mem[1167:1160] } <= { data_i[7:0] };
    end 
    if(N935) begin
      { mem[1159:1152] } <= { data_i[7:0] };
    end 
    if(N934) begin
      { mem[1151:1144] } <= { data_i[7:0] };
    end 
    if(N933) begin
      { mem[1143:1136] } <= { data_i[7:0] };
    end 
    if(N932) begin
      { mem[1135:1128] } <= { data_i[7:0] };
    end 
    if(N931) begin
      { mem[1127:1120] } <= { data_i[7:0] };
    end 
    if(N930) begin
      { mem[1119:1112] } <= { data_i[7:0] };
    end 
    if(N929) begin
      { mem[1111:1104] } <= { data_i[7:0] };
    end 
    if(N928) begin
      { mem[1103:1096] } <= { data_i[7:0] };
    end 
    if(N927) begin
      { mem[1095:1088] } <= { data_i[7:0] };
    end 
    if(N926) begin
      { mem[1087:1080] } <= { data_i[7:0] };
    end 
    if(N925) begin
      { mem[1079:1072] } <= { data_i[7:0] };
    end 
    if(N924) begin
      { mem[1071:1064] } <= { data_i[7:0] };
    end 
    if(N923) begin
      { mem[1063:1056] } <= { data_i[7:0] };
    end 
    if(N922) begin
      { mem[1055:1048] } <= { data_i[7:0] };
    end 
    if(N921) begin
      { mem[1047:1040] } <= { data_i[7:0] };
    end 
    if(N920) begin
      { mem[1039:1032] } <= { data_i[7:0] };
    end 
    if(N919) begin
      { mem[1031:1024] } <= { data_i[7:0] };
    end 
    if(N918) begin
      { mem[1023:1016] } <= { data_i[7:0] };
    end 
    if(N917) begin
      { mem[1015:1008] } <= { data_i[7:0] };
    end 
    if(N916) begin
      { mem[1007:1000] } <= { data_i[7:0] };
    end 
    if(N915) begin
      { mem[999:992] } <= { data_i[7:0] };
    end 
    if(N914) begin
      { mem[991:984] } <= { data_i[7:0] };
    end 
    if(N913) begin
      { mem[983:976] } <= { data_i[7:0] };
    end 
    if(N912) begin
      { mem[975:968] } <= { data_i[7:0] };
    end 
    if(N911) begin
      { mem[967:960] } <= { data_i[7:0] };
    end 
    if(N910) begin
      { mem[959:952] } <= { data_i[7:0] };
    end 
    if(N909) begin
      { mem[951:944] } <= { data_i[7:0] };
    end 
    if(N908) begin
      { mem[943:936] } <= { data_i[7:0] };
    end 
    if(N907) begin
      { mem[935:928] } <= { data_i[7:0] };
    end 
    if(N906) begin
      { mem[927:920] } <= { data_i[7:0] };
    end 
    if(N905) begin
      { mem[919:912] } <= { data_i[7:0] };
    end 
    if(N904) begin
      { mem[911:904] } <= { data_i[7:0] };
    end 
    if(N903) begin
      { mem[903:896] } <= { data_i[7:0] };
    end 
    if(N902) begin
      { mem[895:888] } <= { data_i[7:0] };
    end 
    if(N901) begin
      { mem[887:880] } <= { data_i[7:0] };
    end 
    if(N900) begin
      { mem[879:872] } <= { data_i[7:0] };
    end 
    if(N899) begin
      { mem[871:864] } <= { data_i[7:0] };
    end 
    if(N898) begin
      { mem[863:856] } <= { data_i[7:0] };
    end 
    if(N897) begin
      { mem[855:848] } <= { data_i[7:0] };
    end 
    if(N896) begin
      { mem[847:840] } <= { data_i[7:0] };
    end 
    if(N895) begin
      { mem[839:832] } <= { data_i[7:0] };
    end 
    if(N894) begin
      { mem[831:824] } <= { data_i[7:0] };
    end 
    if(N893) begin
      { mem[823:816] } <= { data_i[7:0] };
    end 
    if(N892) begin
      { mem[815:808] } <= { data_i[7:0] };
    end 
    if(N891) begin
      { mem[807:800] } <= { data_i[7:0] };
    end 
    if(N890) begin
      { mem[799:792] } <= { data_i[7:0] };
    end 
    if(N889) begin
      { mem[791:784] } <= { data_i[7:0] };
    end 
    if(N888) begin
      { mem[783:776] } <= { data_i[7:0] };
    end 
    if(N887) begin
      { mem[775:768] } <= { data_i[7:0] };
    end 
    if(N886) begin
      { mem[767:760] } <= { data_i[7:0] };
    end 
    if(N885) begin
      { mem[759:752] } <= { data_i[7:0] };
    end 
    if(N884) begin
      { mem[751:744] } <= { data_i[7:0] };
    end 
    if(N883) begin
      { mem[743:736] } <= { data_i[7:0] };
    end 
    if(N882) begin
      { mem[735:728] } <= { data_i[7:0] };
    end 
    if(N881) begin
      { mem[727:720] } <= { data_i[7:0] };
    end 
    if(N880) begin
      { mem[719:712] } <= { data_i[7:0] };
    end 
    if(N879) begin
      { mem[711:704] } <= { data_i[7:0] };
    end 
    if(N878) begin
      { mem[703:696] } <= { data_i[7:0] };
    end 
    if(N877) begin
      { mem[695:688] } <= { data_i[7:0] };
    end 
    if(N876) begin
      { mem[687:680] } <= { data_i[7:0] };
    end 
    if(N875) begin
      { mem[679:672] } <= { data_i[7:0] };
    end 
    if(N874) begin
      { mem[671:664] } <= { data_i[7:0] };
    end 
    if(N873) begin
      { mem[663:656] } <= { data_i[7:0] };
    end 
    if(N872) begin
      { mem[655:648] } <= { data_i[7:0] };
    end 
    if(N871) begin
      { mem[647:640] } <= { data_i[7:0] };
    end 
    if(N870) begin
      { mem[639:632] } <= { data_i[7:0] };
    end 
    if(N869) begin
      { mem[631:624] } <= { data_i[7:0] };
    end 
    if(N868) begin
      { mem[623:616] } <= { data_i[7:0] };
    end 
    if(N867) begin
      { mem[615:608] } <= { data_i[7:0] };
    end 
    if(N866) begin
      { mem[607:600] } <= { data_i[7:0] };
    end 
    if(N865) begin
      { mem[599:592] } <= { data_i[7:0] };
    end 
    if(N864) begin
      { mem[591:584] } <= { data_i[7:0] };
    end 
    if(N863) begin
      { mem[583:576] } <= { data_i[7:0] };
    end 
    if(N862) begin
      { mem[575:568] } <= { data_i[7:0] };
    end 
    if(N861) begin
      { mem[567:560] } <= { data_i[7:0] };
    end 
    if(N860) begin
      { mem[559:552] } <= { data_i[7:0] };
    end 
    if(N859) begin
      { mem[551:544] } <= { data_i[7:0] };
    end 
    if(N858) begin
      { mem[543:536] } <= { data_i[7:0] };
    end 
    if(N857) begin
      { mem[535:528] } <= { data_i[7:0] };
    end 
    if(N856) begin
      { mem[527:520] } <= { data_i[7:0] };
    end 
    if(N855) begin
      { mem[519:512] } <= { data_i[7:0] };
    end 
    if(N854) begin
      { mem[511:504] } <= { data_i[7:0] };
    end 
    if(N853) begin
      { mem[503:496] } <= { data_i[7:0] };
    end 
    if(N852) begin
      { mem[495:488] } <= { data_i[7:0] };
    end 
    if(N851) begin
      { mem[487:480] } <= { data_i[7:0] };
    end 
    if(N850) begin
      { mem[479:472] } <= { data_i[7:0] };
    end 
    if(N849) begin
      { mem[471:464] } <= { data_i[7:0] };
    end 
    if(N848) begin
      { mem[463:456] } <= { data_i[7:0] };
    end 
    if(N847) begin
      { mem[455:448] } <= { data_i[7:0] };
    end 
    if(N846) begin
      { mem[447:440] } <= { data_i[7:0] };
    end 
    if(N845) begin
      { mem[439:432] } <= { data_i[7:0] };
    end 
    if(N844) begin
      { mem[431:424] } <= { data_i[7:0] };
    end 
    if(N843) begin
      { mem[423:416] } <= { data_i[7:0] };
    end 
    if(N842) begin
      { mem[415:408] } <= { data_i[7:0] };
    end 
    if(N841) begin
      { mem[407:400] } <= { data_i[7:0] };
    end 
    if(N840) begin
      { mem[399:392] } <= { data_i[7:0] };
    end 
    if(N839) begin
      { mem[391:384] } <= { data_i[7:0] };
    end 
    if(N838) begin
      { mem[383:376] } <= { data_i[7:0] };
    end 
    if(N837) begin
      { mem[375:368] } <= { data_i[7:0] };
    end 
    if(N836) begin
      { mem[367:360] } <= { data_i[7:0] };
    end 
    if(N835) begin
      { mem[359:352] } <= { data_i[7:0] };
    end 
    if(N834) begin
      { mem[351:344] } <= { data_i[7:0] };
    end 
    if(N833) begin
      { mem[343:336] } <= { data_i[7:0] };
    end 
    if(N832) begin
      { mem[335:328] } <= { data_i[7:0] };
    end 
    if(N831) begin
      { mem[327:320] } <= { data_i[7:0] };
    end 
    if(N830) begin
      { mem[319:312] } <= { data_i[7:0] };
    end 
    if(N829) begin
      { mem[311:304] } <= { data_i[7:0] };
    end 
    if(N828) begin
      { mem[303:296] } <= { data_i[7:0] };
    end 
    if(N827) begin
      { mem[295:288] } <= { data_i[7:0] };
    end 
    if(N826) begin
      { mem[287:280] } <= { data_i[7:0] };
    end 
    if(N825) begin
      { mem[279:272] } <= { data_i[7:0] };
    end 
    if(N824) begin
      { mem[271:264] } <= { data_i[7:0] };
    end 
    if(N823) begin
      { mem[263:256] } <= { data_i[7:0] };
    end 
    if(N822) begin
      { mem[255:248] } <= { data_i[7:0] };
    end 
    if(N821) begin
      { mem[247:240] } <= { data_i[7:0] };
    end 
    if(N820) begin
      { mem[239:232] } <= { data_i[7:0] };
    end 
    if(N819) begin
      { mem[231:224] } <= { data_i[7:0] };
    end 
    if(N818) begin
      { mem[223:216] } <= { data_i[7:0] };
    end 
    if(N817) begin
      { mem[215:208] } <= { data_i[7:0] };
    end 
    if(N816) begin
      { mem[207:200] } <= { data_i[7:0] };
    end 
    if(N815) begin
      { mem[199:192] } <= { data_i[7:0] };
    end 
    if(N814) begin
      { mem[191:184] } <= { data_i[7:0] };
    end 
    if(N813) begin
      { mem[183:176] } <= { data_i[7:0] };
    end 
    if(N812) begin
      { mem[175:168] } <= { data_i[7:0] };
    end 
    if(N811) begin
      { mem[167:160] } <= { data_i[7:0] };
    end 
    if(N810) begin
      { mem[159:152] } <= { data_i[7:0] };
    end 
    if(N809) begin
      { mem[151:144] } <= { data_i[7:0] };
    end 
    if(N808) begin
      { mem[143:136] } <= { data_i[7:0] };
    end 
    if(N807) begin
      { mem[135:128] } <= { data_i[7:0] };
    end 
    if(N806) begin
      { mem[127:120] } <= { data_i[7:0] };
    end 
    if(N805) begin
      { mem[119:112] } <= { data_i[7:0] };
    end 
    if(N804) begin
      { mem[111:104] } <= { data_i[7:0] };
    end 
    if(N803) begin
      { mem[103:96] } <= { data_i[7:0] };
    end 
    if(N802) begin
      { mem[95:88] } <= { data_i[7:0] };
    end 
    if(N801) begin
      { mem[87:80] } <= { data_i[7:0] };
    end 
    if(N800) begin
      { mem[79:72] } <= { data_i[7:0] };
    end 
    if(N799) begin
      { mem[71:64] } <= { data_i[7:0] };
    end 
    if(N798) begin
      { mem[63:56] } <= { data_i[7:0] };
    end 
    if(N797) begin
      { mem[55:48] } <= { data_i[7:0] };
    end 
    if(N796) begin
      { mem[47:40] } <= { data_i[7:0] };
    end 
    if(N795) begin
      { mem[39:32] } <= { data_i[7:0] };
    end 
    if(N794) begin
      { mem[31:24] } <= { data_i[7:0] };
    end 
    if(N793) begin
      { mem[23:16] } <= { data_i[7:0] };
    end 
    if(N792) begin
      { mem[15:8] } <= { data_i[7:0] };
    end 
    if(N791) begin
      { mem[7:0] } <= { data_i[7:0] };
    end 
  end


endmodule



module bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_i,
  data_o
);

  input [7:0] data_i;
  input [7:0] addr_i;
  output [7:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [7:0] data_o;

  bsg_mem_1rw_sync_synth_width_p8_els_p256_latch_last_read_p1
  synth
  (
    .clk_i(clk_i),
    .v_i(v_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_mem_1rw_sync_mask_write_byte_synth_els_p256_latch_last_read_p1_data_width_p128
(
  clk_i,
  reset_i,
  v_i,
  w_i,
  addr_i,
  data_i,
  write_mask_i,
  data_o
);

  input [7:0] addr_i;
  input [127:0] data_i;
  input [15:0] write_mask_i;
  output [127:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [127:0] data_o;
  wire n_0_net_,n_1_net_,n_2_net_,n_3_net_,n_4_net_,n_5_net_,n_6_net_,n_7_net_,
  n_8_net_,n_9_net_,n_10_net_,n_11_net_,n_12_net_,n_13_net_,n_14_net_,n_15_net_;

  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_0__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[7:0]),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(n_0_net_),
    .data_o(data_o[7:0])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_1__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[15:8]),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(n_1_net_),
    .data_o(data_o[15:8])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_2__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[23:16]),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(n_2_net_),
    .data_o(data_o[23:16])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_3__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[31:24]),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(n_3_net_),
    .data_o(data_o[31:24])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_4__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[39:32]),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(n_4_net_),
    .data_o(data_o[39:32])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_5__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[47:40]),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(n_5_net_),
    .data_o(data_o[47:40])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_6__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[55:48]),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(n_6_net_),
    .data_o(data_o[55:48])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_7__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[63:56]),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(n_7_net_),
    .data_o(data_o[63:56])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_8__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[71:64]),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(n_8_net_),
    .data_o(data_o[71:64])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_9__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[79:72]),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(n_9_net_),
    .data_o(data_o[79:72])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_10__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[87:80]),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(n_10_net_),
    .data_o(data_o[87:80])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_11__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[95:88]),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(n_11_net_),
    .data_o(data_o[95:88])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_12__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[103:96]),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(n_12_net_),
    .data_o(data_o[103:96])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_13__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[111:104]),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(n_13_net_),
    .data_o(data_o[111:104])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_14__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[119:112]),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(n_14_net_),
    .data_o(data_o[119:112])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_15__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[127:120]),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(n_15_net_),
    .data_o(data_o[127:120])
  );

  assign n_0_net_ = w_i & write_mask_i[0];
  assign n_1_net_ = w_i & write_mask_i[1];
  assign n_2_net_ = w_i & write_mask_i[2];
  assign n_3_net_ = w_i & write_mask_i[3];
  assign n_4_net_ = w_i & write_mask_i[4];
  assign n_5_net_ = w_i & write_mask_i[5];
  assign n_6_net_ = w_i & write_mask_i[6];
  assign n_7_net_ = w_i & write_mask_i[7];
  assign n_8_net_ = w_i & write_mask_i[8];
  assign n_9_net_ = w_i & write_mask_i[9];
  assign n_10_net_ = w_i & write_mask_i[10];
  assign n_11_net_ = w_i & write_mask_i[11];
  assign n_12_net_ = w_i & write_mask_i[12];
  assign n_13_net_ = w_i & write_mask_i[13];
  assign n_14_net_ = w_i & write_mask_i[14];
  assign n_15_net_ = w_i & write_mask_i[15];

endmodule



module bsg_mem_1rw_sync_mask_write_byte_els_p256_data_width_p128_latch_last_read_p1
(
  clk_i,
  reset_i,
  v_i,
  w_i,
  addr_i,
  data_i,
  write_mask_i,
  data_o
);

  input [7:0] addr_i;
  input [127:0] data_i;
  input [15:0] write_mask_i;
  output [127:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [127:0] data_o;

  bsg_mem_1rw_sync_mask_write_byte_synth_els_p256_latch_last_read_p1_data_width_p128
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .w_i(w_i),
    .addr_i(addr_i),
    .data_i(data_i),
    .write_mask_i(write_mask_i),
    .data_o(data_o)
  );


endmodule



module bsg_scan_width_p4_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [3:0] i;
  output [3:0] o;
  wire [3:0] o;
  wire t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__3_ = i[0] | 1'b0;
  assign t_1__2_ = i[1] | i[0];
  assign t_1__1_ = i[2] | i[1];
  assign t_1__0_ = i[3] | i[2];
  assign o[0] = t_1__3_ | 1'b0;
  assign o[1] = t_1__2_ | 1'b0;
  assign o[2] = t_1__1_ | t_1__3_;
  assign o[3] = t_1__0_ | t_1__2_;

endmodule



module bsg_priority_encode_one_hot_out_width_p4_lo_to_hi_p1
(
  i,
  o
);

  input [3:0] i;
  output [3:0] o;
  wire [3:0] o;
  wire N0,N1,N2;
  wire [3:1] scan_lo;

  bsg_scan_width_p4_or_p1_lo_to_hi_p1
  genblk1_scan
  (
    .i(i),
    .o({ scan_lo, o[0:0] })
  );

  assign o[3] = scan_lo[3] & N0;
  assign N0 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N1;
  assign N1 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N2;
  assign N2 = ~o[0];

endmodule



module bsg_encode_one_hot_width_p1
(
  i,
  addr_o,
  v_o
);

  input [0:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  assign v_o = i[0];
  assign addr_o[0] = 1'b0;

endmodule



module bsg_encode_one_hot_width_p2
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o,aligned_vs;
  wire v_o;
  wire [1:0] aligned_addrs;

  bsg_encode_one_hot_width_p1
  aligned_left
  (
    .i(i[0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p1
  aligned_right
  (
    .i(i[1]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[0])
  );

  assign v_o = addr_o[0] | aligned_vs[0];

endmodule



module bsg_encode_one_hot_width_p4_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [3:0] i;
  output [1:0] addr_o;
  output v_o;
  wire [1:0] addr_o,aligned_addrs;
  wire v_o;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p2
  aligned_left
  (
    .i(i[1:0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p2
  aligned_right
  (
    .i(i[3:2]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[1])
  );

  assign v_o = addr_o[1] | aligned_vs[0];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[1];

endmodule



module bsg_priority_encode_width_p4_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [3:0] i;
  output [1:0] addr_o;
  output v_o;
  wire [1:0] addr_o;
  wire v_o;
  wire [3:0] enc_lo;

  bsg_priority_encode_one_hot_out_width_p4_lo_to_hi_p1
  a
  (
    .i(i),
    .o(enc_lo)
  );


  bsg_encode_one_hot_width_p4_lo_to_hi_p1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o),
    .v_o(v_o)
  );


endmodule



module bsg_dff_en_width_p7_harden_p0_strength_p0
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [6:0] data_i;
  output [6:0] data_o;
  input clk_i;
  input en_i;
  reg [6:0] data_o;

  always @(posedge clk_i) begin
    if(en_i) begin
      { data_o[6:0] } <= { data_i[6:0] };
    end 
  end


endmodule



module bsg_dff_en_bypass_width_p7
(
  clk_i,
  en_i,
  data_i,
  data_o
);

  input [6:0] data_i;
  output [6:0] data_o;
  input clk_i;
  input en_i;
  wire [6:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_en_width_p7_harden_p0_strength_p0
  dff
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .en_i(en_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_mem_1rw_sync_mask_write_bit_synth_width_p7_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [6:0] data_i;
  input [5:0] addr_i;
  input [6:0] w_mask_i;
  output [6:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [6:0] data_o,data_out;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,read_en,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,
  llr_read_en_r,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,
  N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
  N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,
  N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
  N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,
  N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,
  N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,
  N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,
  N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,
  N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,
  N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,
  N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,
  N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,
  N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,
  N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,
  N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,
  N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,
  N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,
  N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,
  N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,
  N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,
  N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,
  N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,
  N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,
  N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,
  N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,
  N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,
  N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,
  N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,
  N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,
  N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,
  N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,
  N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,
  N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,
  N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,
  N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,
  N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,
  N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
  N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,
  N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,
  N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,
  N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,
  N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,
  N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,
  N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,
  N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,
  N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,
  N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,
  N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,
  N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,
  N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,
  N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,
  N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,
  N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,
  N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,
  N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,
  N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,
  N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,
  N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,
  N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,
  N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,
  N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,
  N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,
  N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,
  N1141;
  reg [5:0] addr_r;
  reg [447:0] mem;
  assign data_out[6] = (N82)? mem[6] : 
                       (N84)? mem[13] : 
                       (N86)? mem[20] : 
                       (N88)? mem[27] : 
                       (N90)? mem[34] : 
                       (N92)? mem[41] : 
                       (N94)? mem[48] : 
                       (N96)? mem[55] : 
                       (N98)? mem[62] : 
                       (N100)? mem[69] : 
                       (N102)? mem[76] : 
                       (N104)? mem[83] : 
                       (N106)? mem[90] : 
                       (N108)? mem[97] : 
                       (N110)? mem[104] : 
                       (N112)? mem[111] : 
                       (N114)? mem[118] : 
                       (N116)? mem[125] : 
                       (N118)? mem[132] : 
                       (N120)? mem[139] : 
                       (N122)? mem[146] : 
                       (N124)? mem[153] : 
                       (N126)? mem[160] : 
                       (N128)? mem[167] : 
                       (N130)? mem[174] : 
                       (N132)? mem[181] : 
                       (N134)? mem[188] : 
                       (N136)? mem[195] : 
                       (N138)? mem[202] : 
                       (N140)? mem[209] : 
                       (N142)? mem[216] : 
                       (N144)? mem[223] : 
                       (N83)? mem[230] : 
                       (N85)? mem[237] : 
                       (N87)? mem[244] : 
                       (N89)? mem[251] : 
                       (N91)? mem[258] : 
                       (N93)? mem[265] : 
                       (N95)? mem[272] : 
                       (N97)? mem[279] : 
                       (N99)? mem[286] : 
                       (N101)? mem[293] : 
                       (N103)? mem[300] : 
                       (N105)? mem[307] : 
                       (N107)? mem[314] : 
                       (N109)? mem[321] : 
                       (N111)? mem[328] : 
                       (N113)? mem[335] : 
                       (N115)? mem[342] : 
                       (N117)? mem[349] : 
                       (N119)? mem[356] : 
                       (N121)? mem[363] : 
                       (N123)? mem[370] : 
                       (N125)? mem[377] : 
                       (N127)? mem[384] : 
                       (N129)? mem[391] : 
                       (N131)? mem[398] : 
                       (N133)? mem[405] : 
                       (N135)? mem[412] : 
                       (N137)? mem[419] : 
                       (N139)? mem[426] : 
                       (N141)? mem[433] : 
                       (N143)? mem[440] : 
                       (N145)? mem[447] : 1'b0;
  assign data_out[5] = (N82)? mem[5] : 
                       (N84)? mem[12] : 
                       (N86)? mem[19] : 
                       (N88)? mem[26] : 
                       (N90)? mem[33] : 
                       (N92)? mem[40] : 
                       (N94)? mem[47] : 
                       (N96)? mem[54] : 
                       (N98)? mem[61] : 
                       (N100)? mem[68] : 
                       (N102)? mem[75] : 
                       (N104)? mem[82] : 
                       (N106)? mem[89] : 
                       (N108)? mem[96] : 
                       (N110)? mem[103] : 
                       (N112)? mem[110] : 
                       (N114)? mem[117] : 
                       (N116)? mem[124] : 
                       (N118)? mem[131] : 
                       (N120)? mem[138] : 
                       (N122)? mem[145] : 
                       (N124)? mem[152] : 
                       (N126)? mem[159] : 
                       (N128)? mem[166] : 
                       (N130)? mem[173] : 
                       (N132)? mem[180] : 
                       (N134)? mem[187] : 
                       (N136)? mem[194] : 
                       (N138)? mem[201] : 
                       (N140)? mem[208] : 
                       (N142)? mem[215] : 
                       (N144)? mem[222] : 
                       (N83)? mem[229] : 
                       (N85)? mem[236] : 
                       (N87)? mem[243] : 
                       (N89)? mem[250] : 
                       (N91)? mem[257] : 
                       (N93)? mem[264] : 
                       (N95)? mem[271] : 
                       (N97)? mem[278] : 
                       (N99)? mem[285] : 
                       (N101)? mem[292] : 
                       (N103)? mem[299] : 
                       (N105)? mem[306] : 
                       (N107)? mem[313] : 
                       (N109)? mem[320] : 
                       (N111)? mem[327] : 
                       (N113)? mem[334] : 
                       (N115)? mem[341] : 
                       (N117)? mem[348] : 
                       (N119)? mem[355] : 
                       (N121)? mem[362] : 
                       (N123)? mem[369] : 
                       (N125)? mem[376] : 
                       (N127)? mem[383] : 
                       (N129)? mem[390] : 
                       (N131)? mem[397] : 
                       (N133)? mem[404] : 
                       (N135)? mem[411] : 
                       (N137)? mem[418] : 
                       (N139)? mem[425] : 
                       (N141)? mem[432] : 
                       (N143)? mem[439] : 
                       (N145)? mem[446] : 1'b0;
  assign data_out[4] = (N82)? mem[4] : 
                       (N84)? mem[11] : 
                       (N86)? mem[18] : 
                       (N88)? mem[25] : 
                       (N90)? mem[32] : 
                       (N92)? mem[39] : 
                       (N94)? mem[46] : 
                       (N96)? mem[53] : 
                       (N98)? mem[60] : 
                       (N100)? mem[67] : 
                       (N102)? mem[74] : 
                       (N104)? mem[81] : 
                       (N106)? mem[88] : 
                       (N108)? mem[95] : 
                       (N110)? mem[102] : 
                       (N112)? mem[109] : 
                       (N114)? mem[116] : 
                       (N116)? mem[123] : 
                       (N118)? mem[130] : 
                       (N120)? mem[137] : 
                       (N122)? mem[144] : 
                       (N124)? mem[151] : 
                       (N126)? mem[158] : 
                       (N128)? mem[165] : 
                       (N130)? mem[172] : 
                       (N132)? mem[179] : 
                       (N134)? mem[186] : 
                       (N136)? mem[193] : 
                       (N138)? mem[200] : 
                       (N140)? mem[207] : 
                       (N142)? mem[214] : 
                       (N144)? mem[221] : 
                       (N83)? mem[228] : 
                       (N85)? mem[235] : 
                       (N87)? mem[242] : 
                       (N89)? mem[249] : 
                       (N91)? mem[256] : 
                       (N93)? mem[263] : 
                       (N95)? mem[270] : 
                       (N97)? mem[277] : 
                       (N99)? mem[284] : 
                       (N101)? mem[291] : 
                       (N103)? mem[298] : 
                       (N105)? mem[305] : 
                       (N107)? mem[312] : 
                       (N109)? mem[319] : 
                       (N111)? mem[326] : 
                       (N113)? mem[333] : 
                       (N115)? mem[340] : 
                       (N117)? mem[347] : 
                       (N119)? mem[354] : 
                       (N121)? mem[361] : 
                       (N123)? mem[368] : 
                       (N125)? mem[375] : 
                       (N127)? mem[382] : 
                       (N129)? mem[389] : 
                       (N131)? mem[396] : 
                       (N133)? mem[403] : 
                       (N135)? mem[410] : 
                       (N137)? mem[417] : 
                       (N139)? mem[424] : 
                       (N141)? mem[431] : 
                       (N143)? mem[438] : 
                       (N145)? mem[445] : 1'b0;
  assign data_out[3] = (N82)? mem[3] : 
                       (N84)? mem[10] : 
                       (N86)? mem[17] : 
                       (N88)? mem[24] : 
                       (N90)? mem[31] : 
                       (N92)? mem[38] : 
                       (N94)? mem[45] : 
                       (N96)? mem[52] : 
                       (N98)? mem[59] : 
                       (N100)? mem[66] : 
                       (N102)? mem[73] : 
                       (N104)? mem[80] : 
                       (N106)? mem[87] : 
                       (N108)? mem[94] : 
                       (N110)? mem[101] : 
                       (N112)? mem[108] : 
                       (N114)? mem[115] : 
                       (N116)? mem[122] : 
                       (N118)? mem[129] : 
                       (N120)? mem[136] : 
                       (N122)? mem[143] : 
                       (N124)? mem[150] : 
                       (N126)? mem[157] : 
                       (N128)? mem[164] : 
                       (N130)? mem[171] : 
                       (N132)? mem[178] : 
                       (N134)? mem[185] : 
                       (N136)? mem[192] : 
                       (N138)? mem[199] : 
                       (N140)? mem[206] : 
                       (N142)? mem[213] : 
                       (N144)? mem[220] : 
                       (N83)? mem[227] : 
                       (N85)? mem[234] : 
                       (N87)? mem[241] : 
                       (N89)? mem[248] : 
                       (N91)? mem[255] : 
                       (N93)? mem[262] : 
                       (N95)? mem[269] : 
                       (N97)? mem[276] : 
                       (N99)? mem[283] : 
                       (N101)? mem[290] : 
                       (N103)? mem[297] : 
                       (N105)? mem[304] : 
                       (N107)? mem[311] : 
                       (N109)? mem[318] : 
                       (N111)? mem[325] : 
                       (N113)? mem[332] : 
                       (N115)? mem[339] : 
                       (N117)? mem[346] : 
                       (N119)? mem[353] : 
                       (N121)? mem[360] : 
                       (N123)? mem[367] : 
                       (N125)? mem[374] : 
                       (N127)? mem[381] : 
                       (N129)? mem[388] : 
                       (N131)? mem[395] : 
                       (N133)? mem[402] : 
                       (N135)? mem[409] : 
                       (N137)? mem[416] : 
                       (N139)? mem[423] : 
                       (N141)? mem[430] : 
                       (N143)? mem[437] : 
                       (N145)? mem[444] : 1'b0;
  assign data_out[2] = (N82)? mem[2] : 
                       (N84)? mem[9] : 
                       (N86)? mem[16] : 
                       (N88)? mem[23] : 
                       (N90)? mem[30] : 
                       (N92)? mem[37] : 
                       (N94)? mem[44] : 
                       (N96)? mem[51] : 
                       (N98)? mem[58] : 
                       (N100)? mem[65] : 
                       (N102)? mem[72] : 
                       (N104)? mem[79] : 
                       (N106)? mem[86] : 
                       (N108)? mem[93] : 
                       (N110)? mem[100] : 
                       (N112)? mem[107] : 
                       (N114)? mem[114] : 
                       (N116)? mem[121] : 
                       (N118)? mem[128] : 
                       (N120)? mem[135] : 
                       (N122)? mem[142] : 
                       (N124)? mem[149] : 
                       (N126)? mem[156] : 
                       (N128)? mem[163] : 
                       (N130)? mem[170] : 
                       (N132)? mem[177] : 
                       (N134)? mem[184] : 
                       (N136)? mem[191] : 
                       (N138)? mem[198] : 
                       (N140)? mem[205] : 
                       (N142)? mem[212] : 
                       (N144)? mem[219] : 
                       (N83)? mem[226] : 
                       (N85)? mem[233] : 
                       (N87)? mem[240] : 
                       (N89)? mem[247] : 
                       (N91)? mem[254] : 
                       (N93)? mem[261] : 
                       (N95)? mem[268] : 
                       (N97)? mem[275] : 
                       (N99)? mem[282] : 
                       (N101)? mem[289] : 
                       (N103)? mem[296] : 
                       (N105)? mem[303] : 
                       (N107)? mem[310] : 
                       (N109)? mem[317] : 
                       (N111)? mem[324] : 
                       (N113)? mem[331] : 
                       (N115)? mem[338] : 
                       (N117)? mem[345] : 
                       (N119)? mem[352] : 
                       (N121)? mem[359] : 
                       (N123)? mem[366] : 
                       (N125)? mem[373] : 
                       (N127)? mem[380] : 
                       (N129)? mem[387] : 
                       (N131)? mem[394] : 
                       (N133)? mem[401] : 
                       (N135)? mem[408] : 
                       (N137)? mem[415] : 
                       (N139)? mem[422] : 
                       (N141)? mem[429] : 
                       (N143)? mem[436] : 
                       (N145)? mem[443] : 1'b0;
  assign data_out[1] = (N82)? mem[1] : 
                       (N84)? mem[8] : 
                       (N86)? mem[15] : 
                       (N88)? mem[22] : 
                       (N90)? mem[29] : 
                       (N92)? mem[36] : 
                       (N94)? mem[43] : 
                       (N96)? mem[50] : 
                       (N98)? mem[57] : 
                       (N100)? mem[64] : 
                       (N102)? mem[71] : 
                       (N104)? mem[78] : 
                       (N106)? mem[85] : 
                       (N108)? mem[92] : 
                       (N110)? mem[99] : 
                       (N112)? mem[106] : 
                       (N114)? mem[113] : 
                       (N116)? mem[120] : 
                       (N118)? mem[127] : 
                       (N120)? mem[134] : 
                       (N122)? mem[141] : 
                       (N124)? mem[148] : 
                       (N126)? mem[155] : 
                       (N128)? mem[162] : 
                       (N130)? mem[169] : 
                       (N132)? mem[176] : 
                       (N134)? mem[183] : 
                       (N136)? mem[190] : 
                       (N138)? mem[197] : 
                       (N140)? mem[204] : 
                       (N142)? mem[211] : 
                       (N144)? mem[218] : 
                       (N83)? mem[225] : 
                       (N85)? mem[232] : 
                       (N87)? mem[239] : 
                       (N89)? mem[246] : 
                       (N91)? mem[253] : 
                       (N93)? mem[260] : 
                       (N95)? mem[267] : 
                       (N97)? mem[274] : 
                       (N99)? mem[281] : 
                       (N101)? mem[288] : 
                       (N103)? mem[295] : 
                       (N105)? mem[302] : 
                       (N107)? mem[309] : 
                       (N109)? mem[316] : 
                       (N111)? mem[323] : 
                       (N113)? mem[330] : 
                       (N115)? mem[337] : 
                       (N117)? mem[344] : 
                       (N119)? mem[351] : 
                       (N121)? mem[358] : 
                       (N123)? mem[365] : 
                       (N125)? mem[372] : 
                       (N127)? mem[379] : 
                       (N129)? mem[386] : 
                       (N131)? mem[393] : 
                       (N133)? mem[400] : 
                       (N135)? mem[407] : 
                       (N137)? mem[414] : 
                       (N139)? mem[421] : 
                       (N141)? mem[428] : 
                       (N143)? mem[435] : 
                       (N145)? mem[442] : 1'b0;
  assign data_out[0] = (N82)? mem[0] : 
                       (N84)? mem[7] : 
                       (N86)? mem[14] : 
                       (N88)? mem[21] : 
                       (N90)? mem[28] : 
                       (N92)? mem[35] : 
                       (N94)? mem[42] : 
                       (N96)? mem[49] : 
                       (N98)? mem[56] : 
                       (N100)? mem[63] : 
                       (N102)? mem[70] : 
                       (N104)? mem[77] : 
                       (N106)? mem[84] : 
                       (N108)? mem[91] : 
                       (N110)? mem[98] : 
                       (N112)? mem[105] : 
                       (N114)? mem[112] : 
                       (N116)? mem[119] : 
                       (N118)? mem[126] : 
                       (N120)? mem[133] : 
                       (N122)? mem[140] : 
                       (N124)? mem[147] : 
                       (N126)? mem[154] : 
                       (N128)? mem[161] : 
                       (N130)? mem[168] : 
                       (N132)? mem[175] : 
                       (N134)? mem[182] : 
                       (N136)? mem[189] : 
                       (N138)? mem[196] : 
                       (N140)? mem[203] : 
                       (N142)? mem[210] : 
                       (N144)? mem[217] : 
                       (N83)? mem[224] : 
                       (N85)? mem[231] : 
                       (N87)? mem[238] : 
                       (N89)? mem[245] : 
                       (N91)? mem[252] : 
                       (N93)? mem[259] : 
                       (N95)? mem[266] : 
                       (N97)? mem[273] : 
                       (N99)? mem[280] : 
                       (N101)? mem[287] : 
                       (N103)? mem[294] : 
                       (N105)? mem[301] : 
                       (N107)? mem[308] : 
                       (N109)? mem[315] : 
                       (N111)? mem[322] : 
                       (N113)? mem[329] : 
                       (N115)? mem[336] : 
                       (N117)? mem[343] : 
                       (N119)? mem[350] : 
                       (N121)? mem[357] : 
                       (N123)? mem[364] : 
                       (N125)? mem[371] : 
                       (N127)? mem[378] : 
                       (N129)? mem[385] : 
                       (N131)? mem[392] : 
                       (N133)? mem[399] : 
                       (N135)? mem[406] : 
                       (N137)? mem[413] : 
                       (N139)? mem[420] : 
                       (N141)? mem[427] : 
                       (N143)? mem[434] : 
                       (N145)? mem[441] : 1'b0;

  bsg_dff_width_p1
  llr_read_en_dff
  (
    .clk_i(clk_i),
    .data_i(read_en),
    .data_o(llr_read_en_r)
  );


  bsg_dff_en_bypass_width_p7
  llr_dff_bypass
  (
    .clk_i(clk_i),
    .en_i(llr_read_en_r),
    .data_i(data_out),
    .data_o(data_o)
  );

  assign N1115 = ~addr_i[5];
  assign N1116 = addr_i[3] & addr_i[4];
  assign N1117 = N0 & addr_i[4];
  assign N0 = ~addr_i[3];
  assign N1118 = addr_i[3] & N1;
  assign N1 = ~addr_i[4];
  assign N1119 = N2 & N3;
  assign N2 = ~addr_i[3];
  assign N3 = ~addr_i[4];
  assign N1120 = addr_i[5] & N1116;
  assign N1121 = addr_i[5] & N1117;
  assign N1122 = addr_i[5] & N1118;
  assign N1123 = addr_i[5] & N1119;
  assign N1124 = N1115 & N1116;
  assign N1125 = N1115 & N1117;
  assign N1126 = N1115 & N1118;
  assign N1127 = N1115 & N1119;
  assign N1128 = ~addr_i[2];
  assign N1129 = addr_i[0] & addr_i[1];
  assign N1130 = N4 & addr_i[1];
  assign N4 = ~addr_i[0];
  assign N1131 = addr_i[0] & N5;
  assign N5 = ~addr_i[1];
  assign N1132 = N6 & N7;
  assign N6 = ~addr_i[0];
  assign N7 = ~addr_i[1];
  assign N1133 = addr_i[2] & N1129;
  assign N1134 = addr_i[2] & N1130;
  assign N1135 = addr_i[2] & N1131;
  assign N1136 = addr_i[2] & N1132;
  assign N1137 = N1128 & N1129;
  assign N1138 = N1128 & N1130;
  assign N1139 = N1128 & N1131;
  assign N1140 = N1128 & N1132;
  assign N602 = N1120 & N1133;
  assign N601 = N1120 & N1134;
  assign N600 = N1120 & N1135;
  assign N599 = N1120 & N1136;
  assign N598 = N1120 & N1137;
  assign N597 = N1120 & N1138;
  assign N596 = N1120 & N1139;
  assign N595 = N1120 & N1140;
  assign N594 = N1121 & N1133;
  assign N593 = N1121 & N1134;
  assign N592 = N1121 & N1135;
  assign N591 = N1121 & N1136;
  assign N590 = N1121 & N1137;
  assign N589 = N1121 & N1138;
  assign N588 = N1121 & N1139;
  assign N587 = N1121 & N1140;
  assign N586 = N1122 & N1133;
  assign N585 = N1122 & N1134;
  assign N584 = N1122 & N1135;
  assign N583 = N1122 & N1136;
  assign N582 = N1122 & N1137;
  assign N581 = N1122 & N1138;
  assign N580 = N1122 & N1139;
  assign N579 = N1122 & N1140;
  assign N578 = N1123 & N1133;
  assign N577 = N1123 & N1134;
  assign N576 = N1123 & N1135;
  assign N575 = N1123 & N1136;
  assign N574 = N1123 & N1137;
  assign N573 = N1123 & N1138;
  assign N572 = N1123 & N1139;
  assign N571 = N1123 & N1140;
  assign N570 = N1124 & N1133;
  assign N569 = N1124 & N1134;
  assign N568 = N1124 & N1135;
  assign N567 = N1124 & N1136;
  assign N566 = N1124 & N1137;
  assign N565 = N1124 & N1138;
  assign N564 = N1124 & N1139;
  assign N563 = N1124 & N1140;
  assign N562 = N1125 & N1133;
  assign N561 = N1125 & N1134;
  assign N560 = N1125 & N1135;
  assign N559 = N1125 & N1136;
  assign N558 = N1125 & N1137;
  assign N557 = N1125 & N1138;
  assign N556 = N1125 & N1139;
  assign N555 = N1125 & N1140;
  assign N554 = N1126 & N1133;
  assign N553 = N1126 & N1134;
  assign N552 = N1126 & N1135;
  assign N551 = N1126 & N1136;
  assign N550 = N1126 & N1137;
  assign N549 = N1126 & N1138;
  assign N548 = N1126 & N1139;
  assign N547 = N1126 & N1140;
  assign N546 = N1127 & N1133;
  assign N545 = N1127 & N1134;
  assign N544 = N1127 & N1135;
  assign N543 = N1127 & N1136;
  assign N542 = N1127 & N1137;
  assign N541 = N1127 & N1138;
  assign N540 = N1127 & N1139;
  assign N539 = N1127 & N1140;
  assign { N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149 } = (N8)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N148)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_mask_i[0];
  assign { N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214 } = (N9)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N213)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N9 = w_mask_i[1];
  assign { N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279 } = (N10)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N278)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = w_mask_i[2];
  assign { N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344 } = (N11)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N343)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = w_mask_i[3];
  assign { N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409 } = (N12)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N408)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = w_mask_i[4];
  assign { N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474 } = (N13)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N473)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = w_mask_i[5];
  assign { N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603 } = (N14)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N538)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N14 = w_mask_i[6];
  assign { N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667 } = (N15)? { N666, N537, N472, N407, N342, N277, N212, N665, N536, N471, N406, N341, N276, N211, N664, N535, N470, N405, N340, N275, N210, N663, N534, N469, N404, N339, N274, N209, N662, N533, N468, N403, N338, N273, N208, N661, N532, N467, N402, N337, N272, N207, N660, N531, N466, N401, N336, N271, N206, N659, N530, N465, N400, N335, N270, N205, N658, N529, N464, N399, N334, N269, N204, N657, N528, N463, N398, N333, N268, N203, N656, N527, N462, N397, N332, N267, N202, N655, N526, N461, N396, N331, N266, N201, N654, N525, N460, N395, N330, N265, N200, N653, N524, N459, N394, N329, N264, N199, N652, N523, N458, N393, N328, N263, N198, N651, N522, N457, N392, N327, N262, N197, N650, N521, N456, N391, N326, N261, N196, N649, N520, N455, N390, N325, N260, N195, N648, N519, N454, N389, N324, N259, N194, N647, N518, N453, N388, N323, N258, N193, N646, N517, N452, N387, N322, N257, N192, N645, N516, N451, N386, N321, N256, N191, N644, N515, N450, N385, N320, N255, N190, N643, N514, N449, N384, N319, N254, N189, N642, N513, N448, N383, N318, N253, N188, N641, N512, N447, N382, N317, N252, N187, N640, N511, N446, N381, N316, N251, N186, N639, N510, N445, N380, N315, N250, N185, N638, N509, N444, N379, N314, N249, N184, N637, N508, N443, N378, N313, N248, N183, N636, N507, N442, N377, N312, N247, N182, N635, N506, N441, N376, N311, N246, N181, N634, N505, N440, N375, N310, N245, N180, N633, N504, N439, N374, N309, N244, N179, N632, N503, N438, N373, N308, N243, N178, N631, N502, N437, N372, N307, N242, N177, N630, N501, N436, N371, N306, N241, N176, N629, N500, N435, N370, N305, N240, N175, N628, N499, N434, N369, N304, N239, N174, N627, N498, N433, N368, N303, N238, N173, N626, N497, N432, N367, N302, N237, N172, N625, N496, N431, N366, N301, N236, N171, N624, N495, N430, N365, N300, N235, N170, N623, N494, N429, N364, N299, N234, N169, N622, N493, N428, N363, N298, N233, N168, N621, N492, N427, N362, N297, N232, N167, N620, N491, N426, N361, N296, N231, N166, N619, N490, N425, N360, N295, N230, N165, N618, N489, N424, N359, N294, N229, N164, N617, N488, N423, N358, N293, N228, N163, N616, N487, N422, N357, N292, N227, N162, N615, N486, N421, N356, N291, N226, N161, N614, N485, N420, N355, N290, N225, N160, N613, N484, N419, N354, N289, N224, N159, N612, N483, N418, N353, N288, N223, N158, N611, N482, N417, N352, N287, N222, N157, N610, N481, N416, N351, N286, N221, N156, N609, N480, N415, N350, N285, N220, N155, N608, N479, N414, N349, N284, N219, N154, N607, N478, N413, N348, N283, N218, N153, N606, N477, N412, N347, N282, N217, N152, N605, N476, N411, N346, N281, N216, N151, N604, N475, N410, N345, N280, N215, N150, N603, N474, N409, N344, N279, N214, N149 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 (N147)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = N146;
  assign read_en = v_i & N1141;
  assign N1141 = ~w_i;
  assign N16 = ~addr_r[0];
  assign N17 = ~addr_r[1];
  assign N18 = N16 & N17;
  assign N19 = N16 & addr_r[1];
  assign N20 = addr_r[0] & N17;
  assign N21 = addr_r[0] & addr_r[1];
  assign N22 = ~addr_r[2];
  assign N23 = N18 & N22;
  assign N24 = N18 & addr_r[2];
  assign N25 = N20 & N22;
  assign N26 = N20 & addr_r[2];
  assign N27 = N19 & N22;
  assign N28 = N19 & addr_r[2];
  assign N29 = N21 & N22;
  assign N30 = N21 & addr_r[2];
  assign N31 = ~addr_r[3];
  assign N32 = N23 & N31;
  assign N33 = N23 & addr_r[3];
  assign N34 = N25 & N31;
  assign N35 = N25 & addr_r[3];
  assign N36 = N27 & N31;
  assign N37 = N27 & addr_r[3];
  assign N38 = N29 & N31;
  assign N39 = N29 & addr_r[3];
  assign N40 = N24 & N31;
  assign N41 = N24 & addr_r[3];
  assign N42 = N26 & N31;
  assign N43 = N26 & addr_r[3];
  assign N44 = N28 & N31;
  assign N45 = N28 & addr_r[3];
  assign N46 = N30 & N31;
  assign N47 = N30 & addr_r[3];
  assign N48 = ~addr_r[4];
  assign N49 = N32 & N48;
  assign N50 = N32 & addr_r[4];
  assign N51 = N34 & N48;
  assign N52 = N34 & addr_r[4];
  assign N53 = N36 & N48;
  assign N54 = N36 & addr_r[4];
  assign N55 = N38 & N48;
  assign N56 = N38 & addr_r[4];
  assign N57 = N40 & N48;
  assign N58 = N40 & addr_r[4];
  assign N59 = N42 & N48;
  assign N60 = N42 & addr_r[4];
  assign N61 = N44 & N48;
  assign N62 = N44 & addr_r[4];
  assign N63 = N46 & N48;
  assign N64 = N46 & addr_r[4];
  assign N65 = N33 & N48;
  assign N66 = N33 & addr_r[4];
  assign N67 = N35 & N48;
  assign N68 = N35 & addr_r[4];
  assign N69 = N37 & N48;
  assign N70 = N37 & addr_r[4];
  assign N71 = N39 & N48;
  assign N72 = N39 & addr_r[4];
  assign N73 = N41 & N48;
  assign N74 = N41 & addr_r[4];
  assign N75 = N43 & N48;
  assign N76 = N43 & addr_r[4];
  assign N77 = N45 & N48;
  assign N78 = N45 & addr_r[4];
  assign N79 = N47 & N48;
  assign N80 = N47 & addr_r[4];
  assign N81 = ~addr_r[5];
  assign N82 = N49 & N81;
  assign N83 = N49 & addr_r[5];
  assign N84 = N51 & N81;
  assign N85 = N51 & addr_r[5];
  assign N86 = N53 & N81;
  assign N87 = N53 & addr_r[5];
  assign N88 = N55 & N81;
  assign N89 = N55 & addr_r[5];
  assign N90 = N57 & N81;
  assign N91 = N57 & addr_r[5];
  assign N92 = N59 & N81;
  assign N93 = N59 & addr_r[5];
  assign N94 = N61 & N81;
  assign N95 = N61 & addr_r[5];
  assign N96 = N63 & N81;
  assign N97 = N63 & addr_r[5];
  assign N98 = N65 & N81;
  assign N99 = N65 & addr_r[5];
  assign N100 = N67 & N81;
  assign N101 = N67 & addr_r[5];
  assign N102 = N69 & N81;
  assign N103 = N69 & addr_r[5];
  assign N104 = N71 & N81;
  assign N105 = N71 & addr_r[5];
  assign N106 = N73 & N81;
  assign N107 = N73 & addr_r[5];
  assign N108 = N75 & N81;
  assign N109 = N75 & addr_r[5];
  assign N110 = N77 & N81;
  assign N111 = N77 & addr_r[5];
  assign N112 = N79 & N81;
  assign N113 = N79 & addr_r[5];
  assign N114 = N50 & N81;
  assign N115 = N50 & addr_r[5];
  assign N116 = N52 & N81;
  assign N117 = N52 & addr_r[5];
  assign N118 = N54 & N81;
  assign N119 = N54 & addr_r[5];
  assign N120 = N56 & N81;
  assign N121 = N56 & addr_r[5];
  assign N122 = N58 & N81;
  assign N123 = N58 & addr_r[5];
  assign N124 = N60 & N81;
  assign N125 = N60 & addr_r[5];
  assign N126 = N62 & N81;
  assign N127 = N62 & addr_r[5];
  assign N128 = N64 & N81;
  assign N129 = N64 & addr_r[5];
  assign N130 = N66 & N81;
  assign N131 = N66 & addr_r[5];
  assign N132 = N68 & N81;
  assign N133 = N68 & addr_r[5];
  assign N134 = N70 & N81;
  assign N135 = N70 & addr_r[5];
  assign N136 = N72 & N81;
  assign N137 = N72 & addr_r[5];
  assign N138 = N74 & N81;
  assign N139 = N74 & addr_r[5];
  assign N140 = N76 & N81;
  assign N141 = N76 & addr_r[5];
  assign N142 = N78 & N81;
  assign N143 = N78 & addr_r[5];
  assign N144 = N80 & N81;
  assign N145 = N80 & addr_r[5];
  assign N146 = v_i & w_i;
  assign N147 = ~N146;
  assign N148 = ~w_mask_i[0];
  assign N213 = ~w_mask_i[1];
  assign N278 = ~w_mask_i[2];
  assign N343 = ~w_mask_i[3];
  assign N408 = ~w_mask_i[4];
  assign N473 = ~w_mask_i[5];
  assign N538 = ~w_mask_i[6];

  always @(posedge clk_i) begin
    if(1'b1) begin
      { addr_r[5:0] } <= { addr_i[5:0] };
    end 
    if(N1114) begin
      { mem[447:447] } <= { data_i[6:6] };
    end 
    if(N1113) begin
      { mem[446:446] } <= { data_i[5:5] };
    end 
    if(N1112) begin
      { mem[445:445] } <= { data_i[4:4] };
    end 
    if(N1111) begin
      { mem[444:444] } <= { data_i[3:3] };
    end 
    if(N1110) begin
      { mem[443:443] } <= { data_i[2:2] };
    end 
    if(N1109) begin
      { mem[442:442] } <= { data_i[1:1] };
    end 
    if(N1108) begin
      { mem[441:441] } <= { data_i[0:0] };
    end 
    if(N1107) begin
      { mem[440:440] } <= { data_i[6:6] };
    end 
    if(N1106) begin
      { mem[439:439] } <= { data_i[5:5] };
    end 
    if(N1105) begin
      { mem[438:438] } <= { data_i[4:4] };
    end 
    if(N1104) begin
      { mem[437:437] } <= { data_i[3:3] };
    end 
    if(N1103) begin
      { mem[436:436] } <= { data_i[2:2] };
    end 
    if(N1102) begin
      { mem[435:435] } <= { data_i[1:1] };
    end 
    if(N1101) begin
      { mem[434:434] } <= { data_i[0:0] };
    end 
    if(N1100) begin
      { mem[433:433] } <= { data_i[6:6] };
    end 
    if(N1099) begin
      { mem[432:432] } <= { data_i[5:5] };
    end 
    if(N1098) begin
      { mem[431:431] } <= { data_i[4:4] };
    end 
    if(N1097) begin
      { mem[430:430] } <= { data_i[3:3] };
    end 
    if(N1096) begin
      { mem[429:429] } <= { data_i[2:2] };
    end 
    if(N1095) begin
      { mem[428:428] } <= { data_i[1:1] };
    end 
    if(N1094) begin
      { mem[427:427] } <= { data_i[0:0] };
    end 
    if(N1093) begin
      { mem[426:426] } <= { data_i[6:6] };
    end 
    if(N1092) begin
      { mem[425:425] } <= { data_i[5:5] };
    end 
    if(N1091) begin
      { mem[424:424] } <= { data_i[4:4] };
    end 
    if(N1090) begin
      { mem[423:423] } <= { data_i[3:3] };
    end 
    if(N1089) begin
      { mem[422:422] } <= { data_i[2:2] };
    end 
    if(N1088) begin
      { mem[421:421] } <= { data_i[1:1] };
    end 
    if(N1087) begin
      { mem[420:420] } <= { data_i[0:0] };
    end 
    if(N1086) begin
      { mem[419:419] } <= { data_i[6:6] };
    end 
    if(N1085) begin
      { mem[418:418] } <= { data_i[5:5] };
    end 
    if(N1084) begin
      { mem[417:417] } <= { data_i[4:4] };
    end 
    if(N1083) begin
      { mem[416:416] } <= { data_i[3:3] };
    end 
    if(N1082) begin
      { mem[415:415] } <= { data_i[2:2] };
    end 
    if(N1081) begin
      { mem[414:414] } <= { data_i[1:1] };
    end 
    if(N1080) begin
      { mem[413:413] } <= { data_i[0:0] };
    end 
    if(N1079) begin
      { mem[412:412] } <= { data_i[6:6] };
    end 
    if(N1078) begin
      { mem[411:411] } <= { data_i[5:5] };
    end 
    if(N1077) begin
      { mem[410:410] } <= { data_i[4:4] };
    end 
    if(N1076) begin
      { mem[409:409] } <= { data_i[3:3] };
    end 
    if(N1075) begin
      { mem[408:408] } <= { data_i[2:2] };
    end 
    if(N1074) begin
      { mem[407:407] } <= { data_i[1:1] };
    end 
    if(N1073) begin
      { mem[406:406] } <= { data_i[0:0] };
    end 
    if(N1072) begin
      { mem[405:405] } <= { data_i[6:6] };
    end 
    if(N1071) begin
      { mem[404:404] } <= { data_i[5:5] };
    end 
    if(N1070) begin
      { mem[403:403] } <= { data_i[4:4] };
    end 
    if(N1069) begin
      { mem[402:402] } <= { data_i[3:3] };
    end 
    if(N1068) begin
      { mem[401:401] } <= { data_i[2:2] };
    end 
    if(N1067) begin
      { mem[400:400] } <= { data_i[1:1] };
    end 
    if(N1066) begin
      { mem[399:399] } <= { data_i[0:0] };
    end 
    if(N1065) begin
      { mem[398:398] } <= { data_i[6:6] };
    end 
    if(N1064) begin
      { mem[397:397] } <= { data_i[5:5] };
    end 
    if(N1063) begin
      { mem[396:396] } <= { data_i[4:4] };
    end 
    if(N1062) begin
      { mem[395:395] } <= { data_i[3:3] };
    end 
    if(N1061) begin
      { mem[394:394] } <= { data_i[2:2] };
    end 
    if(N1060) begin
      { mem[393:393] } <= { data_i[1:1] };
    end 
    if(N1059) begin
      { mem[392:392] } <= { data_i[0:0] };
    end 
    if(N1058) begin
      { mem[391:391] } <= { data_i[6:6] };
    end 
    if(N1057) begin
      { mem[390:390] } <= { data_i[5:5] };
    end 
    if(N1056) begin
      { mem[389:389] } <= { data_i[4:4] };
    end 
    if(N1055) begin
      { mem[388:388] } <= { data_i[3:3] };
    end 
    if(N1054) begin
      { mem[387:387] } <= { data_i[2:2] };
    end 
    if(N1053) begin
      { mem[386:386] } <= { data_i[1:1] };
    end 
    if(N1052) begin
      { mem[385:385] } <= { data_i[0:0] };
    end 
    if(N1051) begin
      { mem[384:384] } <= { data_i[6:6] };
    end 
    if(N1050) begin
      { mem[383:383] } <= { data_i[5:5] };
    end 
    if(N1049) begin
      { mem[382:382] } <= { data_i[4:4] };
    end 
    if(N1048) begin
      { mem[381:381] } <= { data_i[3:3] };
    end 
    if(N1047) begin
      { mem[380:380] } <= { data_i[2:2] };
    end 
    if(N1046) begin
      { mem[379:379] } <= { data_i[1:1] };
    end 
    if(N1045) begin
      { mem[378:378] } <= { data_i[0:0] };
    end 
    if(N1044) begin
      { mem[377:377] } <= { data_i[6:6] };
    end 
    if(N1043) begin
      { mem[376:376] } <= { data_i[5:5] };
    end 
    if(N1042) begin
      { mem[375:375] } <= { data_i[4:4] };
    end 
    if(N1041) begin
      { mem[374:374] } <= { data_i[3:3] };
    end 
    if(N1040) begin
      { mem[373:373] } <= { data_i[2:2] };
    end 
    if(N1039) begin
      { mem[372:372] } <= { data_i[1:1] };
    end 
    if(N1038) begin
      { mem[371:371] } <= { data_i[0:0] };
    end 
    if(N1037) begin
      { mem[370:370] } <= { data_i[6:6] };
    end 
    if(N1036) begin
      { mem[369:369] } <= { data_i[5:5] };
    end 
    if(N1035) begin
      { mem[368:368] } <= { data_i[4:4] };
    end 
    if(N1034) begin
      { mem[367:367] } <= { data_i[3:3] };
    end 
    if(N1033) begin
      { mem[366:366] } <= { data_i[2:2] };
    end 
    if(N1032) begin
      { mem[365:365] } <= { data_i[1:1] };
    end 
    if(N1031) begin
      { mem[364:364] } <= { data_i[0:0] };
    end 
    if(N1030) begin
      { mem[363:363] } <= { data_i[6:6] };
    end 
    if(N1029) begin
      { mem[362:362] } <= { data_i[5:5] };
    end 
    if(N1028) begin
      { mem[361:361] } <= { data_i[4:4] };
    end 
    if(N1027) begin
      { mem[360:360] } <= { data_i[3:3] };
    end 
    if(N1026) begin
      { mem[359:359] } <= { data_i[2:2] };
    end 
    if(N1025) begin
      { mem[358:358] } <= { data_i[1:1] };
    end 
    if(N1024) begin
      { mem[357:357] } <= { data_i[0:0] };
    end 
    if(N1023) begin
      { mem[356:356] } <= { data_i[6:6] };
    end 
    if(N1022) begin
      { mem[355:355] } <= { data_i[5:5] };
    end 
    if(N1021) begin
      { mem[354:354] } <= { data_i[4:4] };
    end 
    if(N1020) begin
      { mem[353:353] } <= { data_i[3:3] };
    end 
    if(N1019) begin
      { mem[352:352] } <= { data_i[2:2] };
    end 
    if(N1018) begin
      { mem[351:351] } <= { data_i[1:1] };
    end 
    if(N1017) begin
      { mem[350:350] } <= { data_i[0:0] };
    end 
    if(N1016) begin
      { mem[349:349] } <= { data_i[6:6] };
    end 
    if(N1015) begin
      { mem[348:348] } <= { data_i[5:5] };
    end 
    if(N1014) begin
      { mem[347:347] } <= { data_i[4:4] };
    end 
    if(N1013) begin
      { mem[346:346] } <= { data_i[3:3] };
    end 
    if(N1012) begin
      { mem[345:345] } <= { data_i[2:2] };
    end 
    if(N1011) begin
      { mem[344:344] } <= { data_i[1:1] };
    end 
    if(N1010) begin
      { mem[343:343] } <= { data_i[0:0] };
    end 
    if(N1009) begin
      { mem[342:342] } <= { data_i[6:6] };
    end 
    if(N1008) begin
      { mem[341:341] } <= { data_i[5:5] };
    end 
    if(N1007) begin
      { mem[340:340] } <= { data_i[4:4] };
    end 
    if(N1006) begin
      { mem[339:339] } <= { data_i[3:3] };
    end 
    if(N1005) begin
      { mem[338:338] } <= { data_i[2:2] };
    end 
    if(N1004) begin
      { mem[337:337] } <= { data_i[1:1] };
    end 
    if(N1003) begin
      { mem[336:336] } <= { data_i[0:0] };
    end 
    if(N1002) begin
      { mem[335:335] } <= { data_i[6:6] };
    end 
    if(N1001) begin
      { mem[334:334] } <= { data_i[5:5] };
    end 
    if(N1000) begin
      { mem[333:333] } <= { data_i[4:4] };
    end 
    if(N999) begin
      { mem[332:332] } <= { data_i[3:3] };
    end 
    if(N998) begin
      { mem[331:331] } <= { data_i[2:2] };
    end 
    if(N997) begin
      { mem[330:330] } <= { data_i[1:1] };
    end 
    if(N996) begin
      { mem[329:329] } <= { data_i[0:0] };
    end 
    if(N995) begin
      { mem[328:328] } <= { data_i[6:6] };
    end 
    if(N994) begin
      { mem[327:327] } <= { data_i[5:5] };
    end 
    if(N993) begin
      { mem[326:326] } <= { data_i[4:4] };
    end 
    if(N992) begin
      { mem[325:325] } <= { data_i[3:3] };
    end 
    if(N991) begin
      { mem[324:324] } <= { data_i[2:2] };
    end 
    if(N990) begin
      { mem[323:323] } <= { data_i[1:1] };
    end 
    if(N989) begin
      { mem[322:322] } <= { data_i[0:0] };
    end 
    if(N988) begin
      { mem[321:321] } <= { data_i[6:6] };
    end 
    if(N987) begin
      { mem[320:320] } <= { data_i[5:5] };
    end 
    if(N986) begin
      { mem[319:319] } <= { data_i[4:4] };
    end 
    if(N985) begin
      { mem[318:318] } <= { data_i[3:3] };
    end 
    if(N984) begin
      { mem[317:317] } <= { data_i[2:2] };
    end 
    if(N983) begin
      { mem[316:316] } <= { data_i[1:1] };
    end 
    if(N982) begin
      { mem[315:315] } <= { data_i[0:0] };
    end 
    if(N981) begin
      { mem[314:314] } <= { data_i[6:6] };
    end 
    if(N980) begin
      { mem[313:313] } <= { data_i[5:5] };
    end 
    if(N979) begin
      { mem[312:312] } <= { data_i[4:4] };
    end 
    if(N978) begin
      { mem[311:311] } <= { data_i[3:3] };
    end 
    if(N977) begin
      { mem[310:310] } <= { data_i[2:2] };
    end 
    if(N976) begin
      { mem[309:309] } <= { data_i[1:1] };
    end 
    if(N975) begin
      { mem[308:308] } <= { data_i[0:0] };
    end 
    if(N974) begin
      { mem[307:307] } <= { data_i[6:6] };
    end 
    if(N973) begin
      { mem[306:306] } <= { data_i[5:5] };
    end 
    if(N972) begin
      { mem[305:305] } <= { data_i[4:4] };
    end 
    if(N971) begin
      { mem[304:304] } <= { data_i[3:3] };
    end 
    if(N970) begin
      { mem[303:303] } <= { data_i[2:2] };
    end 
    if(N969) begin
      { mem[302:302] } <= { data_i[1:1] };
    end 
    if(N968) begin
      { mem[301:301] } <= { data_i[0:0] };
    end 
    if(N967) begin
      { mem[300:300] } <= { data_i[6:6] };
    end 
    if(N966) begin
      { mem[299:299] } <= { data_i[5:5] };
    end 
    if(N965) begin
      { mem[298:298] } <= { data_i[4:4] };
    end 
    if(N964) begin
      { mem[297:297] } <= { data_i[3:3] };
    end 
    if(N963) begin
      { mem[296:296] } <= { data_i[2:2] };
    end 
    if(N962) begin
      { mem[295:295] } <= { data_i[1:1] };
    end 
    if(N961) begin
      { mem[294:294] } <= { data_i[0:0] };
    end 
    if(N960) begin
      { mem[293:293] } <= { data_i[6:6] };
    end 
    if(N959) begin
      { mem[292:292] } <= { data_i[5:5] };
    end 
    if(N958) begin
      { mem[291:291] } <= { data_i[4:4] };
    end 
    if(N957) begin
      { mem[290:290] } <= { data_i[3:3] };
    end 
    if(N956) begin
      { mem[289:289] } <= { data_i[2:2] };
    end 
    if(N955) begin
      { mem[288:288] } <= { data_i[1:1] };
    end 
    if(N954) begin
      { mem[287:287] } <= { data_i[0:0] };
    end 
    if(N953) begin
      { mem[286:286] } <= { data_i[6:6] };
    end 
    if(N952) begin
      { mem[285:285] } <= { data_i[5:5] };
    end 
    if(N951) begin
      { mem[284:284] } <= { data_i[4:4] };
    end 
    if(N950) begin
      { mem[283:283] } <= { data_i[3:3] };
    end 
    if(N949) begin
      { mem[282:282] } <= { data_i[2:2] };
    end 
    if(N948) begin
      { mem[281:281] } <= { data_i[1:1] };
    end 
    if(N947) begin
      { mem[280:280] } <= { data_i[0:0] };
    end 
    if(N946) begin
      { mem[279:279] } <= { data_i[6:6] };
    end 
    if(N945) begin
      { mem[278:278] } <= { data_i[5:5] };
    end 
    if(N944) begin
      { mem[277:277] } <= { data_i[4:4] };
    end 
    if(N943) begin
      { mem[276:276] } <= { data_i[3:3] };
    end 
    if(N942) begin
      { mem[275:275] } <= { data_i[2:2] };
    end 
    if(N941) begin
      { mem[274:274] } <= { data_i[1:1] };
    end 
    if(N940) begin
      { mem[273:273] } <= { data_i[0:0] };
    end 
    if(N939) begin
      { mem[272:272] } <= { data_i[6:6] };
    end 
    if(N938) begin
      { mem[271:271] } <= { data_i[5:5] };
    end 
    if(N937) begin
      { mem[270:270] } <= { data_i[4:4] };
    end 
    if(N936) begin
      { mem[269:269] } <= { data_i[3:3] };
    end 
    if(N935) begin
      { mem[268:268] } <= { data_i[2:2] };
    end 
    if(N934) begin
      { mem[267:267] } <= { data_i[1:1] };
    end 
    if(N933) begin
      { mem[266:266] } <= { data_i[0:0] };
    end 
    if(N932) begin
      { mem[265:265] } <= { data_i[6:6] };
    end 
    if(N931) begin
      { mem[264:264] } <= { data_i[5:5] };
    end 
    if(N930) begin
      { mem[263:263] } <= { data_i[4:4] };
    end 
    if(N929) begin
      { mem[262:262] } <= { data_i[3:3] };
    end 
    if(N928) begin
      { mem[261:261] } <= { data_i[2:2] };
    end 
    if(N927) begin
      { mem[260:260] } <= { data_i[1:1] };
    end 
    if(N926) begin
      { mem[259:259] } <= { data_i[0:0] };
    end 
    if(N925) begin
      { mem[258:258] } <= { data_i[6:6] };
    end 
    if(N924) begin
      { mem[257:257] } <= { data_i[5:5] };
    end 
    if(N923) begin
      { mem[256:256] } <= { data_i[4:4] };
    end 
    if(N922) begin
      { mem[255:255] } <= { data_i[3:3] };
    end 
    if(N921) begin
      { mem[254:254] } <= { data_i[2:2] };
    end 
    if(N920) begin
      { mem[253:253] } <= { data_i[1:1] };
    end 
    if(N919) begin
      { mem[252:252] } <= { data_i[0:0] };
    end 
    if(N918) begin
      { mem[251:251] } <= { data_i[6:6] };
    end 
    if(N917) begin
      { mem[250:250] } <= { data_i[5:5] };
    end 
    if(N916) begin
      { mem[249:249] } <= { data_i[4:4] };
    end 
    if(N915) begin
      { mem[248:248] } <= { data_i[3:3] };
    end 
    if(N914) begin
      { mem[247:247] } <= { data_i[2:2] };
    end 
    if(N913) begin
      { mem[246:246] } <= { data_i[1:1] };
    end 
    if(N912) begin
      { mem[245:245] } <= { data_i[0:0] };
    end 
    if(N911) begin
      { mem[244:244] } <= { data_i[6:6] };
    end 
    if(N910) begin
      { mem[243:243] } <= { data_i[5:5] };
    end 
    if(N909) begin
      { mem[242:242] } <= { data_i[4:4] };
    end 
    if(N908) begin
      { mem[241:241] } <= { data_i[3:3] };
    end 
    if(N907) begin
      { mem[240:240] } <= { data_i[2:2] };
    end 
    if(N906) begin
      { mem[239:239] } <= { data_i[1:1] };
    end 
    if(N905) begin
      { mem[238:238] } <= { data_i[0:0] };
    end 
    if(N904) begin
      { mem[237:237] } <= { data_i[6:6] };
    end 
    if(N903) begin
      { mem[236:236] } <= { data_i[5:5] };
    end 
    if(N902) begin
      { mem[235:235] } <= { data_i[4:4] };
    end 
    if(N901) begin
      { mem[234:234] } <= { data_i[3:3] };
    end 
    if(N900) begin
      { mem[233:233] } <= { data_i[2:2] };
    end 
    if(N899) begin
      { mem[232:232] } <= { data_i[1:1] };
    end 
    if(N898) begin
      { mem[231:231] } <= { data_i[0:0] };
    end 
    if(N897) begin
      { mem[230:230] } <= { data_i[6:6] };
    end 
    if(N896) begin
      { mem[229:229] } <= { data_i[5:5] };
    end 
    if(N895) begin
      { mem[228:228] } <= { data_i[4:4] };
    end 
    if(N894) begin
      { mem[227:227] } <= { data_i[3:3] };
    end 
    if(N893) begin
      { mem[226:226] } <= { data_i[2:2] };
    end 
    if(N892) begin
      { mem[225:225] } <= { data_i[1:1] };
    end 
    if(N891) begin
      { mem[224:224] } <= { data_i[0:0] };
    end 
    if(N890) begin
      { mem[223:223] } <= { data_i[6:6] };
    end 
    if(N889) begin
      { mem[222:222] } <= { data_i[5:5] };
    end 
    if(N888) begin
      { mem[221:221] } <= { data_i[4:4] };
    end 
    if(N887) begin
      { mem[220:220] } <= { data_i[3:3] };
    end 
    if(N886) begin
      { mem[219:219] } <= { data_i[2:2] };
    end 
    if(N885) begin
      { mem[218:218] } <= { data_i[1:1] };
    end 
    if(N884) begin
      { mem[217:217] } <= { data_i[0:0] };
    end 
    if(N883) begin
      { mem[216:216] } <= { data_i[6:6] };
    end 
    if(N882) begin
      { mem[215:215] } <= { data_i[5:5] };
    end 
    if(N881) begin
      { mem[214:214] } <= { data_i[4:4] };
    end 
    if(N880) begin
      { mem[213:213] } <= { data_i[3:3] };
    end 
    if(N879) begin
      { mem[212:212] } <= { data_i[2:2] };
    end 
    if(N878) begin
      { mem[211:211] } <= { data_i[1:1] };
    end 
    if(N877) begin
      { mem[210:210] } <= { data_i[0:0] };
    end 
    if(N876) begin
      { mem[209:209] } <= { data_i[6:6] };
    end 
    if(N875) begin
      { mem[208:208] } <= { data_i[5:5] };
    end 
    if(N874) begin
      { mem[207:207] } <= { data_i[4:4] };
    end 
    if(N873) begin
      { mem[206:206] } <= { data_i[3:3] };
    end 
    if(N872) begin
      { mem[205:205] } <= { data_i[2:2] };
    end 
    if(N871) begin
      { mem[204:204] } <= { data_i[1:1] };
    end 
    if(N870) begin
      { mem[203:203] } <= { data_i[0:0] };
    end 
    if(N869) begin
      { mem[202:202] } <= { data_i[6:6] };
    end 
    if(N868) begin
      { mem[201:201] } <= { data_i[5:5] };
    end 
    if(N867) begin
      { mem[200:200] } <= { data_i[4:4] };
    end 
    if(N866) begin
      { mem[199:199] } <= { data_i[3:3] };
    end 
    if(N865) begin
      { mem[198:198] } <= { data_i[2:2] };
    end 
    if(N864) begin
      { mem[197:197] } <= { data_i[1:1] };
    end 
    if(N863) begin
      { mem[196:196] } <= { data_i[0:0] };
    end 
    if(N862) begin
      { mem[195:195] } <= { data_i[6:6] };
    end 
    if(N861) begin
      { mem[194:194] } <= { data_i[5:5] };
    end 
    if(N860) begin
      { mem[193:193] } <= { data_i[4:4] };
    end 
    if(N859) begin
      { mem[192:192] } <= { data_i[3:3] };
    end 
    if(N858) begin
      { mem[191:191] } <= { data_i[2:2] };
    end 
    if(N857) begin
      { mem[190:190] } <= { data_i[1:1] };
    end 
    if(N856) begin
      { mem[189:189] } <= { data_i[0:0] };
    end 
    if(N855) begin
      { mem[188:188] } <= { data_i[6:6] };
    end 
    if(N854) begin
      { mem[187:187] } <= { data_i[5:5] };
    end 
    if(N853) begin
      { mem[186:186] } <= { data_i[4:4] };
    end 
    if(N852) begin
      { mem[185:185] } <= { data_i[3:3] };
    end 
    if(N851) begin
      { mem[184:184] } <= { data_i[2:2] };
    end 
    if(N850) begin
      { mem[183:183] } <= { data_i[1:1] };
    end 
    if(N849) begin
      { mem[182:182] } <= { data_i[0:0] };
    end 
    if(N848) begin
      { mem[181:181] } <= { data_i[6:6] };
    end 
    if(N847) begin
      { mem[180:180] } <= { data_i[5:5] };
    end 
    if(N846) begin
      { mem[179:179] } <= { data_i[4:4] };
    end 
    if(N845) begin
      { mem[178:178] } <= { data_i[3:3] };
    end 
    if(N844) begin
      { mem[177:177] } <= { data_i[2:2] };
    end 
    if(N843) begin
      { mem[176:176] } <= { data_i[1:1] };
    end 
    if(N842) begin
      { mem[175:175] } <= { data_i[0:0] };
    end 
    if(N841) begin
      { mem[174:174] } <= { data_i[6:6] };
    end 
    if(N840) begin
      { mem[173:173] } <= { data_i[5:5] };
    end 
    if(N839) begin
      { mem[172:172] } <= { data_i[4:4] };
    end 
    if(N838) begin
      { mem[171:171] } <= { data_i[3:3] };
    end 
    if(N837) begin
      { mem[170:170] } <= { data_i[2:2] };
    end 
    if(N836) begin
      { mem[169:169] } <= { data_i[1:1] };
    end 
    if(N835) begin
      { mem[168:168] } <= { data_i[0:0] };
    end 
    if(N834) begin
      { mem[167:167] } <= { data_i[6:6] };
    end 
    if(N833) begin
      { mem[166:166] } <= { data_i[5:5] };
    end 
    if(N832) begin
      { mem[165:165] } <= { data_i[4:4] };
    end 
    if(N831) begin
      { mem[164:164] } <= { data_i[3:3] };
    end 
    if(N830) begin
      { mem[163:163] } <= { data_i[2:2] };
    end 
    if(N829) begin
      { mem[162:162] } <= { data_i[1:1] };
    end 
    if(N828) begin
      { mem[161:161] } <= { data_i[0:0] };
    end 
    if(N827) begin
      { mem[160:160] } <= { data_i[6:6] };
    end 
    if(N826) begin
      { mem[159:159] } <= { data_i[5:5] };
    end 
    if(N825) begin
      { mem[158:158] } <= { data_i[4:4] };
    end 
    if(N824) begin
      { mem[157:157] } <= { data_i[3:3] };
    end 
    if(N823) begin
      { mem[156:156] } <= { data_i[2:2] };
    end 
    if(N822) begin
      { mem[155:155] } <= { data_i[1:1] };
    end 
    if(N821) begin
      { mem[154:154] } <= { data_i[0:0] };
    end 
    if(N820) begin
      { mem[153:153] } <= { data_i[6:6] };
    end 
    if(N819) begin
      { mem[152:152] } <= { data_i[5:5] };
    end 
    if(N818) begin
      { mem[151:151] } <= { data_i[4:4] };
    end 
    if(N817) begin
      { mem[150:150] } <= { data_i[3:3] };
    end 
    if(N816) begin
      { mem[149:149] } <= { data_i[2:2] };
    end 
    if(N815) begin
      { mem[148:148] } <= { data_i[1:1] };
    end 
    if(N814) begin
      { mem[147:147] } <= { data_i[0:0] };
    end 
    if(N813) begin
      { mem[146:146] } <= { data_i[6:6] };
    end 
    if(N812) begin
      { mem[145:145] } <= { data_i[5:5] };
    end 
    if(N811) begin
      { mem[144:144] } <= { data_i[4:4] };
    end 
    if(N810) begin
      { mem[143:143] } <= { data_i[3:3] };
    end 
    if(N809) begin
      { mem[142:142] } <= { data_i[2:2] };
    end 
    if(N808) begin
      { mem[141:141] } <= { data_i[1:1] };
    end 
    if(N807) begin
      { mem[140:140] } <= { data_i[0:0] };
    end 
    if(N806) begin
      { mem[139:139] } <= { data_i[6:6] };
    end 
    if(N805) begin
      { mem[138:138] } <= { data_i[5:5] };
    end 
    if(N804) begin
      { mem[137:137] } <= { data_i[4:4] };
    end 
    if(N803) begin
      { mem[136:136] } <= { data_i[3:3] };
    end 
    if(N802) begin
      { mem[135:135] } <= { data_i[2:2] };
    end 
    if(N801) begin
      { mem[134:134] } <= { data_i[1:1] };
    end 
    if(N800) begin
      { mem[133:133] } <= { data_i[0:0] };
    end 
    if(N799) begin
      { mem[132:132] } <= { data_i[6:6] };
    end 
    if(N798) begin
      { mem[131:131] } <= { data_i[5:5] };
    end 
    if(N797) begin
      { mem[130:130] } <= { data_i[4:4] };
    end 
    if(N796) begin
      { mem[129:129] } <= { data_i[3:3] };
    end 
    if(N795) begin
      { mem[128:128] } <= { data_i[2:2] };
    end 
    if(N794) begin
      { mem[127:127] } <= { data_i[1:1] };
    end 
    if(N793) begin
      { mem[126:126] } <= { data_i[0:0] };
    end 
    if(N792) begin
      { mem[125:125] } <= { data_i[6:6] };
    end 
    if(N791) begin
      { mem[124:124] } <= { data_i[5:5] };
    end 
    if(N790) begin
      { mem[123:123] } <= { data_i[4:4] };
    end 
    if(N789) begin
      { mem[122:122] } <= { data_i[3:3] };
    end 
    if(N788) begin
      { mem[121:121] } <= { data_i[2:2] };
    end 
    if(N787) begin
      { mem[120:120] } <= { data_i[1:1] };
    end 
    if(N786) begin
      { mem[119:119] } <= { data_i[0:0] };
    end 
    if(N785) begin
      { mem[118:118] } <= { data_i[6:6] };
    end 
    if(N784) begin
      { mem[117:117] } <= { data_i[5:5] };
    end 
    if(N783) begin
      { mem[116:116] } <= { data_i[4:4] };
    end 
    if(N782) begin
      { mem[115:115] } <= { data_i[3:3] };
    end 
    if(N781) begin
      { mem[114:114] } <= { data_i[2:2] };
    end 
    if(N780) begin
      { mem[113:113] } <= { data_i[1:1] };
    end 
    if(N779) begin
      { mem[112:112] } <= { data_i[0:0] };
    end 
    if(N778) begin
      { mem[111:111] } <= { data_i[6:6] };
    end 
    if(N777) begin
      { mem[110:110] } <= { data_i[5:5] };
    end 
    if(N776) begin
      { mem[109:109] } <= { data_i[4:4] };
    end 
    if(N775) begin
      { mem[108:108] } <= { data_i[3:3] };
    end 
    if(N774) begin
      { mem[107:107] } <= { data_i[2:2] };
    end 
    if(N773) begin
      { mem[106:106] } <= { data_i[1:1] };
    end 
    if(N772) begin
      { mem[105:105] } <= { data_i[0:0] };
    end 
    if(N771) begin
      { mem[104:104] } <= { data_i[6:6] };
    end 
    if(N770) begin
      { mem[103:103] } <= { data_i[5:5] };
    end 
    if(N769) begin
      { mem[102:102] } <= { data_i[4:4] };
    end 
    if(N768) begin
      { mem[101:101] } <= { data_i[3:3] };
    end 
    if(N767) begin
      { mem[100:100] } <= { data_i[2:2] };
    end 
    if(N766) begin
      { mem[99:99] } <= { data_i[1:1] };
    end 
    if(N765) begin
      { mem[98:98] } <= { data_i[0:0] };
    end 
    if(N764) begin
      { mem[97:97] } <= { data_i[6:6] };
    end 
    if(N763) begin
      { mem[96:96] } <= { data_i[5:5] };
    end 
    if(N762) begin
      { mem[95:95] } <= { data_i[4:4] };
    end 
    if(N761) begin
      { mem[94:94] } <= { data_i[3:3] };
    end 
    if(N760) begin
      { mem[93:93] } <= { data_i[2:2] };
    end 
    if(N759) begin
      { mem[92:92] } <= { data_i[1:1] };
    end 
    if(N758) begin
      { mem[91:91] } <= { data_i[0:0] };
    end 
    if(N757) begin
      { mem[90:90] } <= { data_i[6:6] };
    end 
    if(N756) begin
      { mem[89:89] } <= { data_i[5:5] };
    end 
    if(N755) begin
      { mem[88:88] } <= { data_i[4:4] };
    end 
    if(N754) begin
      { mem[87:87] } <= { data_i[3:3] };
    end 
    if(N753) begin
      { mem[86:86] } <= { data_i[2:2] };
    end 
    if(N752) begin
      { mem[85:85] } <= { data_i[1:1] };
    end 
    if(N751) begin
      { mem[84:84] } <= { data_i[0:0] };
    end 
    if(N750) begin
      { mem[83:83] } <= { data_i[6:6] };
    end 
    if(N749) begin
      { mem[82:82] } <= { data_i[5:5] };
    end 
    if(N748) begin
      { mem[81:81] } <= { data_i[4:4] };
    end 
    if(N747) begin
      { mem[80:80] } <= { data_i[3:3] };
    end 
    if(N746) begin
      { mem[79:79] } <= { data_i[2:2] };
    end 
    if(N745) begin
      { mem[78:78] } <= { data_i[1:1] };
    end 
    if(N744) begin
      { mem[77:77] } <= { data_i[0:0] };
    end 
    if(N743) begin
      { mem[76:76] } <= { data_i[6:6] };
    end 
    if(N742) begin
      { mem[75:75] } <= { data_i[5:5] };
    end 
    if(N741) begin
      { mem[74:74] } <= { data_i[4:4] };
    end 
    if(N740) begin
      { mem[73:73] } <= { data_i[3:3] };
    end 
    if(N739) begin
      { mem[72:72] } <= { data_i[2:2] };
    end 
    if(N738) begin
      { mem[71:71] } <= { data_i[1:1] };
    end 
    if(N737) begin
      { mem[70:70] } <= { data_i[0:0] };
    end 
    if(N736) begin
      { mem[69:69] } <= { data_i[6:6] };
    end 
    if(N735) begin
      { mem[68:68] } <= { data_i[5:5] };
    end 
    if(N734) begin
      { mem[67:67] } <= { data_i[4:4] };
    end 
    if(N733) begin
      { mem[66:66] } <= { data_i[3:3] };
    end 
    if(N732) begin
      { mem[65:65] } <= { data_i[2:2] };
    end 
    if(N731) begin
      { mem[64:64] } <= { data_i[1:1] };
    end 
    if(N730) begin
      { mem[63:63] } <= { data_i[0:0] };
    end 
    if(N729) begin
      { mem[62:62] } <= { data_i[6:6] };
    end 
    if(N728) begin
      { mem[61:61] } <= { data_i[5:5] };
    end 
    if(N727) begin
      { mem[60:60] } <= { data_i[4:4] };
    end 
    if(N726) begin
      { mem[59:59] } <= { data_i[3:3] };
    end 
    if(N725) begin
      { mem[58:58] } <= { data_i[2:2] };
    end 
    if(N724) begin
      { mem[57:57] } <= { data_i[1:1] };
    end 
    if(N723) begin
      { mem[56:56] } <= { data_i[0:0] };
    end 
    if(N722) begin
      { mem[55:55] } <= { data_i[6:6] };
    end 
    if(N721) begin
      { mem[54:54] } <= { data_i[5:5] };
    end 
    if(N720) begin
      { mem[53:53] } <= { data_i[4:4] };
    end 
    if(N719) begin
      { mem[52:52] } <= { data_i[3:3] };
    end 
    if(N718) begin
      { mem[51:51] } <= { data_i[2:2] };
    end 
    if(N717) begin
      { mem[50:50] } <= { data_i[1:1] };
    end 
    if(N716) begin
      { mem[49:49] } <= { data_i[0:0] };
    end 
    if(N715) begin
      { mem[48:48] } <= { data_i[6:6] };
    end 
    if(N714) begin
      { mem[47:47] } <= { data_i[5:5] };
    end 
    if(N713) begin
      { mem[46:46] } <= { data_i[4:4] };
    end 
    if(N712) begin
      { mem[45:45] } <= { data_i[3:3] };
    end 
    if(N711) begin
      { mem[44:44] } <= { data_i[2:2] };
    end 
    if(N710) begin
      { mem[43:43] } <= { data_i[1:1] };
    end 
    if(N709) begin
      { mem[42:42] } <= { data_i[0:0] };
    end 
    if(N708) begin
      { mem[41:41] } <= { data_i[6:6] };
    end 
    if(N707) begin
      { mem[40:40] } <= { data_i[5:5] };
    end 
    if(N706) begin
      { mem[39:39] } <= { data_i[4:4] };
    end 
    if(N705) begin
      { mem[38:38] } <= { data_i[3:3] };
    end 
    if(N704) begin
      { mem[37:37] } <= { data_i[2:2] };
    end 
    if(N703) begin
      { mem[36:36] } <= { data_i[1:1] };
    end 
    if(N702) begin
      { mem[35:35] } <= { data_i[0:0] };
    end 
    if(N701) begin
      { mem[34:34] } <= { data_i[6:6] };
    end 
    if(N700) begin
      { mem[33:33] } <= { data_i[5:5] };
    end 
    if(N699) begin
      { mem[32:32] } <= { data_i[4:4] };
    end 
    if(N698) begin
      { mem[31:31] } <= { data_i[3:3] };
    end 
    if(N697) begin
      { mem[30:30] } <= { data_i[2:2] };
    end 
    if(N696) begin
      { mem[29:29] } <= { data_i[1:1] };
    end 
    if(N695) begin
      { mem[28:28] } <= { data_i[0:0] };
    end 
    if(N694) begin
      { mem[27:27] } <= { data_i[6:6] };
    end 
    if(N693) begin
      { mem[26:26] } <= { data_i[5:5] };
    end 
    if(N692) begin
      { mem[25:25] } <= { data_i[4:4] };
    end 
    if(N691) begin
      { mem[24:24] } <= { data_i[3:3] };
    end 
    if(N690) begin
      { mem[23:23] } <= { data_i[2:2] };
    end 
    if(N689) begin
      { mem[22:22] } <= { data_i[1:1] };
    end 
    if(N688) begin
      { mem[21:21] } <= { data_i[0:0] };
    end 
    if(N687) begin
      { mem[20:20] } <= { data_i[6:6] };
    end 
    if(N686) begin
      { mem[19:19] } <= { data_i[5:5] };
    end 
    if(N685) begin
      { mem[18:18] } <= { data_i[4:4] };
    end 
    if(N684) begin
      { mem[17:17] } <= { data_i[3:3] };
    end 
    if(N683) begin
      { mem[16:16] } <= { data_i[2:2] };
    end 
    if(N682) begin
      { mem[15:15] } <= { data_i[1:1] };
    end 
    if(N681) begin
      { mem[14:14] } <= { data_i[0:0] };
    end 
    if(N680) begin
      { mem[13:13] } <= { data_i[6:6] };
    end 
    if(N679) begin
      { mem[12:12] } <= { data_i[5:5] };
    end 
    if(N678) begin
      { mem[11:11] } <= { data_i[4:4] };
    end 
    if(N677) begin
      { mem[10:10] } <= { data_i[3:3] };
    end 
    if(N676) begin
      { mem[9:9] } <= { data_i[2:2] };
    end 
    if(N675) begin
      { mem[8:8] } <= { data_i[1:1] };
    end 
    if(N674) begin
      { mem[7:7] } <= { data_i[0:0] };
    end 
    if(N673) begin
      { mem[6:6] } <= { data_i[6:6] };
    end 
    if(N672) begin
      { mem[5:5] } <= { data_i[5:5] };
    end 
    if(N671) begin
      { mem[4:4] } <= { data_i[4:4] };
    end 
    if(N670) begin
      { mem[3:3] } <= { data_i[3:3] };
    end 
    if(N669) begin
      { mem[2:2] } <= { data_i[2:2] };
    end 
    if(N668) begin
      { mem[1:1] } <= { data_i[1:1] };
    end 
    if(N667) begin
      { mem[0:0] } <= { data_i[0:0] };
    end 
  end


endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p7_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [6:0] data_i;
  input [5:0] addr_i;
  input [6:0] w_mask_i;
  output [6:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [6:0] data_o;

  bsg_mem_1rw_sync_mask_write_bit_synth_width_p7_els_p64_latch_last_read_p1
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_mux_width_p1_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [1:0] data_i;
  input [0:0] sel_i;
  output [0:0] data_o;
  wire [0:0] data_o;
  wire N0,N1;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[1] : 1'b0;
  assign N0 = sel_i[0];
  assign N1 = ~sel_i[0];

endmodule



module bsg_lru_pseudo_tree_encode_ways_p4
(
  lru_i,
  way_id_o
);

  input [2:0] lru_i;
  output [1:0] way_id_o;
  wire [1:0] way_id_o;
  assign way_id_o[1] = lru_i[0];

  bsg_mux_width_p1_els_p2
  rank_1__nz_mux
  (
    .data_i(lru_i[2:1]),
    .sel_i(lru_i[0]),
    .data_o(way_id_o[0])
  );


endmodule



module bsg_lru_pseudo_tree_decode_ways_p4
(
  way_id_i,
  data_o,
  mask_o
);

  input [1:0] way_id_i;
  output [2:0] data_o;
  output [2:0] mask_o;
  wire [2:0] data_o,mask_o;
  wire N0,N1;
  assign mask_o[0] = 1'b1;
  assign data_o[0] = 1'b1 & N0;
  assign N0 = ~way_id_i[1];
  assign mask_o[1] = 1'b1 & N0;
  assign data_o[1] = mask_o[1] & N1;
  assign N1 = ~way_id_i[0];
  assign mask_o[2] = 1'b1 & way_id_i[1];
  assign data_o[2] = mask_o[2] & N1;

endmodule



module bsg_decode_num_out_p4
(
  i,
  o
);

  input [1:0] i;
  output [3:0] o;
  wire [3:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_cache_miss_addr_width_p28_data_width_p32_block_size_in_words_p4_sets_p64_ways_p4
(
  clk_i,
  reset_i,
  miss_v_i,
  decode_v_i,
  addr_v_i,
  tag_v_i,
  valid_v_i,
  lock_v_i,
  tag_hit_way_id_i,
  tag_hit_found_i,
  sbuf_empty_i,
  dma_cmd_o,
  dma_way_o,
  dma_addr_o,
  dma_done_i,
  stat_info_i,
  stat_mem_v_o,
  stat_mem_w_o,
  stat_mem_addr_o,
  stat_mem_data_o,
  stat_mem_w_mask_o,
  tag_mem_v_o,
  tag_mem_w_o,
  tag_mem_addr_o,
  tag_mem_data_o,
  tag_mem_w_mask_o,
  done_o,
  recover_o,
  chosen_way_o,
  ack_i
);

  input [15:0] decode_v_i;
  input [27:0] addr_v_i;
  input [71:0] tag_v_i;
  input [3:0] valid_v_i;
  input [3:0] lock_v_i;
  input [1:0] tag_hit_way_id_i;
  output [3:0] dma_cmd_o;
  output [1:0] dma_way_o;
  output [27:0] dma_addr_o;
  input [6:0] stat_info_i;
  output [5:0] stat_mem_addr_o;
  output [6:0] stat_mem_data_o;
  output [6:0] stat_mem_w_mask_o;
  output [5:0] tag_mem_addr_o;
  output [79:0] tag_mem_data_o;
  output [79:0] tag_mem_w_mask_o;
  output [1:0] chosen_way_o;
  input clk_i;
  input reset_i;
  input miss_v_i;
  input tag_hit_found_i;
  input sbuf_empty_i;
  input dma_done_i;
  input ack_i;
  output stat_mem_v_o;
  output stat_mem_w_o;
  output tag_mem_v_o;
  output tag_mem_w_o;
  output done_o;
  output recover_o;
  wire [3:0] dma_cmd_o,chosen_way_decode,miss_state_n;
  wire [27:0] dma_addr_o;
  wire [5:0] stat_mem_addr_o,tag_mem_addr_o;
  wire [6:0] stat_mem_data_o,stat_mem_w_mask_o;
  wire [79:0] tag_mem_data_o,tag_mem_w_mask_o;
  wire [1:0] chosen_way_o,invalid_way_id,lru_way_id,backup_lru_way_id;
  wire stat_mem_v_o,stat_mem_w_o,tag_mem_v_o,tag_mem_w_o,done_o,recover_o,N0,N1,N2,N3,
  N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,n_0_net__3_,n_0_net__2_,
  n_0_net__1_,n_0_net__0_,invalid_exist,goto_flush_op,goto_lock_op,n_2_net__3_,n_2_net__2_,
  n_2_net__1_,n_2_net__0_,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,
  N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,
  N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,
  N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,
  N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,
  N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,
  N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,
  N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,
  N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,
  N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,
  N189,N190,N191,N192,N193,N194;
  wire [2:0] chosen_way_lru_data,chosen_way_lru_mask;
  reg [1:0] dma_way_o;
  reg [3:0] miss_state_r;
  assign dma_addr_o[0] = 1'b0;
  assign dma_addr_o[1] = 1'b0;
  assign tag_mem_addr_o[5] = addr_v_i[9];
  assign stat_mem_addr_o[5] = addr_v_i[9];
  assign tag_mem_addr_o[4] = addr_v_i[8];
  assign stat_mem_addr_o[4] = addr_v_i[8];
  assign tag_mem_addr_o[3] = addr_v_i[7];
  assign stat_mem_addr_o[3] = addr_v_i[7];
  assign tag_mem_addr_o[2] = addr_v_i[6];
  assign stat_mem_addr_o[2] = addr_v_i[6];
  assign tag_mem_addr_o[1] = addr_v_i[5];
  assign stat_mem_addr_o[1] = addr_v_i[5];
  assign tag_mem_addr_o[0] = addr_v_i[4];
  assign stat_mem_addr_o[0] = addr_v_i[4];
  assign dma_cmd_o[0] = tag_mem_data_o[79];
  assign tag_mem_data_o[19] = tag_mem_data_o[79];
  assign tag_mem_data_o[39] = tag_mem_data_o[79];
  assign tag_mem_data_o[59] = tag_mem_data_o[79];

  bsg_priority_encode_width_p4_lo_to_hi_p1
  invalid_way_pe
  (
    .i({ n_0_net__3_, n_0_net__2_, n_0_net__1_, n_0_net__0_ }),
    .addr_o(invalid_way_id),
    .v_o(invalid_exist)
  );


  bsg_lru_pseudo_tree_encode_ways_p4
  lru_encode
  (
    .lru_i(stat_info_i[2:0]),
    .way_id_o(lru_way_id)
  );


  bsg_lru_pseudo_tree_decode_ways_p4
  chosen_way_lru_decode
  (
    .way_id_i(chosen_way_o),
    .data_o(chosen_way_lru_data),
    .mask_o(chosen_way_lru_mask)
  );


  bsg_priority_encode_width_p4_lo_to_hi_p1
  backup_lru_pe
  (
    .i({ n_2_net__3_, n_2_net__2_, n_2_net__1_, n_2_net__0_ }),
    .addr_o(backup_lru_way_id)
  );


  bsg_decode_num_out_p4
  chosen_way_demux
  (
    .i(chosen_way_o),
    .o(chosen_way_decode)
  );

  assign N21 = N17 & N18;
  assign N22 = N19 & N20;
  assign N23 = N21 & N22;
  assign N24 = miss_state_r[3] | N18;
  assign N25 = miss_state_r[1] | miss_state_r[0];
  assign N26 = N24 | N25;
  assign N28 = miss_state_r[3] | miss_state_r[2];
  assign N29 = miss_state_r[1] | N20;
  assign N30 = N28 | N29;
  assign N32 = miss_state_r[3] | miss_state_r[2];
  assign N33 = N19 | miss_state_r[0];
  assign N34 = N32 | N33;
  assign N36 = miss_state_r[3] | miss_state_r[2];
  assign N37 = N19 | N20;
  assign N38 = N36 | N37;
  assign N40 = miss_state_r[3] | N18;
  assign N41 = miss_state_r[1] | N20;
  assign N42 = N40 | N41;
  assign N44 = miss_state_r[3] | N18;
  assign N45 = N19 | miss_state_r[0];
  assign N46 = N44 | N45;
  assign N48 = miss_state_r[3] | N18;
  assign N49 = N19 | N20;
  assign N50 = N48 | N49;
  assign N52 = N17 | miss_state_r[2];
  assign N53 = miss_state_r[1] | miss_state_r[0];
  assign N54 = N52 | N53;
  assign N56 = miss_state_r[3] & miss_state_r[0];
  assign N57 = miss_state_r[3] & miss_state_r[1];
  assign N58 = miss_state_r[3] & miss_state_r[2];
  assign N75 = (N71)? lock_v_i[0] : 
               (N73)? lock_v_i[1] : 
               (N72)? lock_v_i[2] : 
               (N74)? lock_v_i[3] : 1'b0;
  assign N86 = (N82)? stat_info_i[3] : 
               (N84)? stat_info_i[4] : 
               (N83)? stat_info_i[5] : 
               (N85)? stat_info_i[6] : 1'b0;
  assign N87 = (N82)? valid_v_i[0] : 
               (N84)? valid_v_i[1] : 
               (N83)? valid_v_i[2] : 
               (N85)? valid_v_i[3] : 1'b0;
  assign N109 = (N105)? stat_info_i[3] : 
                (N107)? stat_info_i[4] : 
                (N106)? stat_info_i[5] : 
                (N108)? stat_info_i[6] : 1'b0;
  assign N110 = (N105)? valid_v_i[0] : 
                (N107)? valid_v_i[1] : 
                (N106)? valid_v_i[2] : 
                (N108)? valid_v_i[3] : 1'b0;
  assign N119 = (N115)? tag_v_i[17] : 
                (N117)? tag_v_i[35] : 
                (N116)? tag_v_i[53] : 
                (N118)? tag_v_i[71] : 1'b0;
  assign N120 = (N115)? tag_v_i[16] : 
                (N117)? tag_v_i[34] : 
                (N116)? tag_v_i[52] : 
                (N118)? tag_v_i[70] : 1'b0;
  assign N121 = (N115)? tag_v_i[15] : 
                (N117)? tag_v_i[33] : 
                (N116)? tag_v_i[51] : 
                (N118)? tag_v_i[69] : 1'b0;
  assign N122 = (N115)? tag_v_i[14] : 
                (N117)? tag_v_i[32] : 
                (N116)? tag_v_i[50] : 
                (N118)? tag_v_i[68] : 1'b0;
  assign N123 = (N115)? tag_v_i[13] : 
                (N117)? tag_v_i[31] : 
                (N116)? tag_v_i[49] : 
                (N118)? tag_v_i[67] : 1'b0;
  assign N124 = (N115)? tag_v_i[12] : 
                (N117)? tag_v_i[30] : 
                (N116)? tag_v_i[48] : 
                (N118)? tag_v_i[66] : 1'b0;
  assign N125 = (N115)? tag_v_i[11] : 
                (N117)? tag_v_i[29] : 
                (N116)? tag_v_i[47] : 
                (N118)? tag_v_i[65] : 1'b0;
  assign N126 = (N115)? tag_v_i[10] : 
                (N117)? tag_v_i[28] : 
                (N116)? tag_v_i[46] : 
                (N118)? tag_v_i[64] : 1'b0;
  assign N127 = (N115)? tag_v_i[9] : 
                (N117)? tag_v_i[27] : 
                (N116)? tag_v_i[45] : 
                (N118)? tag_v_i[63] : 1'b0;
  assign N128 = (N115)? tag_v_i[8] : 
                (N117)? tag_v_i[26] : 
                (N116)? tag_v_i[44] : 
                (N118)? tag_v_i[62] : 1'b0;
  assign N129 = (N115)? tag_v_i[7] : 
                (N117)? tag_v_i[25] : 
                (N116)? tag_v_i[43] : 
                (N118)? tag_v_i[61] : 1'b0;
  assign N130 = (N115)? tag_v_i[6] : 
                (N117)? tag_v_i[24] : 
                (N116)? tag_v_i[42] : 
                (N118)? tag_v_i[60] : 1'b0;
  assign N131 = (N115)? tag_v_i[5] : 
                (N117)? tag_v_i[23] : 
                (N116)? tag_v_i[41] : 
                (N118)? tag_v_i[59] : 1'b0;
  assign N132 = (N115)? tag_v_i[4] : 
                (N117)? tag_v_i[22] : 
                (N116)? tag_v_i[40] : 
                (N118)? tag_v_i[58] : 1'b0;
  assign N133 = (N115)? tag_v_i[3] : 
                (N117)? tag_v_i[21] : 
                (N116)? tag_v_i[39] : 
                (N118)? tag_v_i[57] : 1'b0;
  assign N134 = (N115)? tag_v_i[2] : 
                (N117)? tag_v_i[20] : 
                (N116)? tag_v_i[38] : 
                (N118)? tag_v_i[56] : 1'b0;
  assign N135 = (N115)? tag_v_i[1] : 
                (N117)? tag_v_i[19] : 
                (N116)? tag_v_i[37] : 
                (N118)? tag_v_i[55] : 1'b0;
  assign N136 = (N115)? tag_v_i[0] : 
                (N117)? tag_v_i[18] : 
                (N116)? tag_v_i[36] : 
                (N118)? tag_v_i[54] : 1'b0;
  assign N142 = (N138)? tag_v_i[17] : 
                (N140)? tag_v_i[35] : 
                (N139)? tag_v_i[53] : 
                (N141)? tag_v_i[71] : 1'b0;
  assign N143 = (N138)? tag_v_i[16] : 
                (N140)? tag_v_i[34] : 
                (N139)? tag_v_i[52] : 
                (N141)? tag_v_i[70] : 1'b0;
  assign N144 = (N138)? tag_v_i[15] : 
                (N140)? tag_v_i[33] : 
                (N139)? tag_v_i[51] : 
                (N141)? tag_v_i[69] : 1'b0;
  assign N145 = (N138)? tag_v_i[14] : 
                (N140)? tag_v_i[32] : 
                (N139)? tag_v_i[50] : 
                (N141)? tag_v_i[68] : 1'b0;
  assign N146 = (N138)? tag_v_i[13] : 
                (N140)? tag_v_i[31] : 
                (N139)? tag_v_i[49] : 
                (N141)? tag_v_i[67] : 1'b0;
  assign N147 = (N138)? tag_v_i[12] : 
                (N140)? tag_v_i[30] : 
                (N139)? tag_v_i[48] : 
                (N141)? tag_v_i[66] : 1'b0;
  assign N148 = (N138)? tag_v_i[11] : 
                (N140)? tag_v_i[29] : 
                (N139)? tag_v_i[47] : 
                (N141)? tag_v_i[65] : 1'b0;
  assign N149 = (N138)? tag_v_i[10] : 
                (N140)? tag_v_i[28] : 
                (N139)? tag_v_i[46] : 
                (N141)? tag_v_i[64] : 1'b0;
  assign N150 = (N138)? tag_v_i[9] : 
                (N140)? tag_v_i[27] : 
                (N139)? tag_v_i[45] : 
                (N141)? tag_v_i[63] : 1'b0;
  assign N151 = (N138)? tag_v_i[8] : 
                (N140)? tag_v_i[26] : 
                (N139)? tag_v_i[44] : 
                (N141)? tag_v_i[62] : 1'b0;
  assign N152 = (N138)? tag_v_i[7] : 
                (N140)? tag_v_i[25] : 
                (N139)? tag_v_i[43] : 
                (N141)? tag_v_i[61] : 1'b0;
  assign N153 = (N138)? tag_v_i[6] : 
                (N140)? tag_v_i[24] : 
                (N139)? tag_v_i[42] : 
                (N141)? tag_v_i[60] : 1'b0;
  assign N154 = (N138)? tag_v_i[5] : 
                (N140)? tag_v_i[23] : 
                (N139)? tag_v_i[41] : 
                (N141)? tag_v_i[59] : 1'b0;
  assign N155 = (N138)? tag_v_i[4] : 
                (N140)? tag_v_i[22] : 
                (N139)? tag_v_i[40] : 
                (N141)? tag_v_i[58] : 1'b0;
  assign N156 = (N138)? tag_v_i[3] : 
                (N140)? tag_v_i[21] : 
                (N139)? tag_v_i[39] : 
                (N141)? tag_v_i[57] : 1'b0;
  assign N157 = (N138)? tag_v_i[2] : 
                (N140)? tag_v_i[20] : 
                (N139)? tag_v_i[38] : 
                (N141)? tag_v_i[56] : 1'b0;
  assign N158 = (N138)? tag_v_i[1] : 
                (N140)? tag_v_i[19] : 
                (N139)? tag_v_i[37] : 
                (N141)? tag_v_i[55] : 1'b0;
  assign N159 = (N138)? tag_v_i[0] : 
                (N140)? tag_v_i[18] : 
                (N139)? tag_v_i[36] : 
                (N141)? tag_v_i[54] : 1'b0;
  assign { N65, N64, N63 } = (N0)? { 1'b0, 1'b0, 1'b1 } : 
                             (N169)? { 1'b0, 1'b1, 1'b0 } : 
                             (N62)? { 1'b1, 1'b0, 1'b0 } : 1'b0;
  assign N0 = goto_flush_op;
  assign { N68, N67, N66 } = (N1)? { N65, N64, N63 } : 
                             (N2)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = miss_v_i;
  assign N2 = N60;
  assign { N79, N78 } = (N3)? invalid_way_id : 
                        (N171)? backup_lru_way_id : 
                        (N77)? lru_way_id : 1'b0;
  assign N3 = invalid_exist;
  assign N89 = ~N88;
  assign { N91, N90 } = (N4)? { N89, N88 } : 
                        (N5)? { 1'b1, 1'b0 } : 1'b0;
  assign N4 = dma_done_i;
  assign N5 = N137;
  assign { N94, N93 } = (N6)? addr_v_i[11:10] : 
                        (N92)? tag_hit_way_id_i : 1'b0;
  assign N6 = decode_v_i[8];
  assign N112 = ~N111;
  assign N161 = (N4)? N160 : 
                (N5)? 1'b1 : 1'b0;
  assign stat_mem_v_o = (N7)? miss_v_i : 
                        (N8)? dma_done_i : 
                        (N9)? 1'b1 : 
                        (N10)? 1'b0 : 
                        (N11)? 1'b0 : 
                        (N12)? 1'b0 : 
                        (N13)? 1'b0 : 
                        (N14)? 1'b0 : 
                        (N15)? 1'b0 : 
                        (N16)? 1'b0 : 1'b0;
  assign N7 = N23;
  assign N8 = tag_mem_data_o[79];
  assign N9 = N31;
  assign N10 = N35;
  assign N11 = dma_cmd_o[1];
  assign N12 = N43;
  assign N13 = N47;
  assign N14 = N51;
  assign N15 = N55;
  assign N16 = N59;
  assign miss_state_n = (N7)? { 1'b0, N68, N67, N66 } : 
                        (N8)? { 1'b0, N91, dma_done_i, N90 } : 
                        (N9)? { 1'b0, N112, 1'b1, 1'b1 } : 
                        (N10)? { 1'b0, 1'b1, 1'b1, 1'b1 } : 
                        (N11)? { 1'b0, dma_done_i, N137, 1'b1 } : 
                        (N12)? { 1'b0, 1'b1, dma_done_i, N161 } : 
                        (N13)? { 1'b0, 1'b1, 1'b1, dma_done_i } : 
                        (N14)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                        (N15)? { N162, 1'b0, 1'b0, 1'b0 } : 
                        (N16)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign chosen_way_o = (N7)? dma_way_o : 
                        (N8)? { N79, N78 } : 
                        (N9)? { N94, N93 } : 
                        (N10)? tag_hit_way_id_i : 
                        (N11)? dma_way_o : 
                        (N12)? dma_way_o : 
                        (N13)? dma_way_o : 
                        (N14)? dma_way_o : 
                        (N15)? dma_way_o : 
                        (N16)? dma_way_o : 1'b0;
  assign dma_cmd_o[2] = (N13)? sbuf_empty_i : 
                        (N165)? 1'b0 : 1'b0;
  assign dma_cmd_o[3] = (N12)? sbuf_empty_i : 
                        (N166)? 1'b0 : 1'b0;
  assign dma_addr_o[3:2] = (N13)? addr_v_i[3:2] : 
                           (N165)? { 1'b0, 1'b0 } : 1'b0;
  assign dma_addr_o[27:4] = (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N8)? addr_v_i[27:4] : 
                            (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N11)? { N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, addr_v_i[9:4] } : 
                            (N12)? { N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, addr_v_i[9:4] } : 
                            (N13)? addr_v_i[27:4] : 
                            (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign stat_mem_w_o = (N7)? 1'b0 : 
                        (N8)? dma_done_i : 
                        (N9)? 1'b1 : 
                        (N10)? 1'b0 : 
                        (N11)? 1'b0 : 
                        (N12)? 1'b0 : 
                        (N13)? 1'b0 : 
                        (N14)? 1'b0 : 
                        (N15)? 1'b0 : 
                        (N16)? 1'b0 : 1'b0;
  assign stat_mem_data_o = (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N8)? { decode_v_i[10:10], decode_v_i[10:10], decode_v_i[10:10], decode_v_i[10:10], chosen_way_lru_data } : 
                           (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign stat_mem_w_mask_o = (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N8)? { chosen_way_decode, chosen_way_lru_mask } : 
                             (N9)? { chosen_way_decode, 1'b0, 1'b0, 1'b0 } : 
                             (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tag_mem_v_o = (N7)? 1'b0 : 
                       (N8)? dma_done_i : 
                       (N9)? 1'b1 : 
                       (N10)? 1'b1 : 
                       (N11)? 1'b0 : 
                       (N12)? 1'b0 : 
                       (N13)? 1'b0 : 
                       (N14)? 1'b0 : 
                       (N15)? 1'b0 : 
                       (N16)? 1'b0 : 1'b0;
  assign tag_mem_w_o = (N7)? 1'b0 : 
                       (N8)? dma_done_i : 
                       (N9)? 1'b1 : 
                       (N10)? 1'b1 : 
                       (N11)? 1'b0 : 
                       (N12)? 1'b0 : 
                       (N13)? 1'b0 : 
                       (N14)? 1'b0 : 
                       (N15)? 1'b0 : 
                       (N16)? 1'b0 : 1'b0;
  assign { tag_mem_w_mask_o[52:40], tag_mem_w_mask_o[37:20], tag_mem_w_mask_o[17:0] } = (N8)? { chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                                                                                        (N167)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { tag_mem_w_mask_o[79:78], tag_mem_w_mask_o[59:58], tag_mem_w_mask_o[39:38], tag_mem_w_mask_o[19:18] } = (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                  (N8)? { chosen_way_decode[3:3], chosen_way_decode[3:2], chosen_way_decode[2:1], chosen_way_decode[1:0], chosen_way_decode[0:0] } : 
                                                                                                                  (N9)? { N101, N102, N99, N100, N97, N98, N95, N96 } : 
                                                                                                                  (N10)? { 1'b0, chosen_way_decode[3:3], 1'b0, chosen_way_decode[2:2], 1'b0, chosen_way_decode[1:1], 1'b0, chosen_way_decode[0:0] } : 
                                                                                                                  (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                  (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                  (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                  (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                  (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                  (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { tag_mem_w_mask_o[77:60], tag_mem_w_mask_o[57:53] } = (N8)? { chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2] } : 
                                                                (N164)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { tag_mem_data_o[77:60], tag_mem_data_o[57:40], tag_mem_data_o[37:20], tag_mem_data_o[17:0] } = (N8)? { addr_v_i[27:10], addr_v_i[27:10], addr_v_i[27:10], addr_v_i[27:10] } : 
                                                                                                         (N164)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { tag_mem_data_o[78:78], tag_mem_data_o[58:58], tag_mem_data_o[38:38], tag_mem_data_o[18:18] } = (N7)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                          (N8)? { decode_v_i[2:2], decode_v_i[2:2], decode_v_i[2:2], decode_v_i[2:2] } : 
                                                                                                          (N9)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                          (N10)? { decode_v_i[2:2], decode_v_i[2:2], decode_v_i[2:2], decode_v_i[2:2] } : 
                                                                                                          (N11)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                          (N12)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                          (N13)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                          (N14)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                          (N15)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                          (N16)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign recover_o = (N7)? 1'b0 : 
                     (N8)? 1'b0 : 
                     (N9)? 1'b0 : 
                     (N10)? 1'b0 : 
                     (N11)? 1'b0 : 
                     (N12)? 1'b0 : 
                     (N13)? 1'b0 : 
                     (N14)? 1'b1 : 
                     (N15)? 1'b0 : 
                     (N16)? 1'b0 : 1'b0;
  assign done_o = (N7)? 1'b0 : 
                  (N8)? 1'b0 : 
                  (N9)? 1'b0 : 
                  (N10)? 1'b0 : 
                  (N11)? 1'b0 : 
                  (N12)? 1'b0 : 
                  (N13)? 1'b0 : 
                  (N14)? 1'b0 : 
                  (N15)? 1'b1 : 
                  (N16)? 1'b0 : 1'b0;
  assign n_0_net__3_ = N172 & N173;
  assign N172 = ~valid_v_i[3];
  assign N173 = ~lock_v_i[3];
  assign n_0_net__2_ = N174 & N175;
  assign N174 = ~valid_v_i[2];
  assign N175 = ~lock_v_i[2];
  assign n_0_net__1_ = N176 & N177;
  assign N176 = ~valid_v_i[1];
  assign N177 = ~lock_v_i[1];
  assign n_0_net__0_ = N178 & N179;
  assign N178 = ~valid_v_i[0];
  assign N179 = ~lock_v_i[0];
  assign goto_flush_op = N181 | decode_v_i[4];
  assign N181 = N180 | decode_v_i[5];
  assign N180 = decode_v_i[8] | decode_v_i[3];
  assign goto_lock_op = decode_v_i[1] | N182;
  assign N182 = decode_v_i[2] & tag_hit_found_i;
  assign n_2_net__3_ = ~lock_v_i[3];
  assign n_2_net__2_ = ~lock_v_i[2];
  assign n_2_net__1_ = ~lock_v_i[1];
  assign n_2_net__0_ = ~lock_v_i[0];
  assign N17 = ~miss_state_r[3];
  assign N18 = ~miss_state_r[2];
  assign N19 = ~miss_state_r[1];
  assign N20 = ~miss_state_r[0];
  assign N27 = ~N26;
  assign N31 = ~N30;
  assign N35 = ~N34;
  assign N39 = ~N38;
  assign N43 = ~N42;
  assign N47 = ~N46;
  assign N51 = ~N50;
  assign N55 = ~N54;
  assign N59 = N56 | N183;
  assign N183 = N57 | N58;
  assign tag_mem_data_o[79] = N27;
  assign dma_cmd_o[1] = N39;
  assign N60 = ~miss_v_i;
  assign N61 = goto_lock_op | goto_flush_op;
  assign N62 = ~N61;
  assign N69 = ~lru_way_id[0];
  assign N70 = ~lru_way_id[1];
  assign N71 = N69 & N70;
  assign N72 = N69 & lru_way_id[1];
  assign N73 = lru_way_id[0] & N70;
  assign N74 = lru_way_id[0] & lru_way_id[1];
  assign N76 = N75 | invalid_exist;
  assign N77 = ~N76;
  assign N80 = ~N78;
  assign N81 = ~N79;
  assign N82 = N80 & N81;
  assign N83 = N80 & N79;
  assign N84 = N78 & N81;
  assign N85 = N78 & N79;
  assign N88 = N86 & N87;
  assign N92 = ~decode_v_i[8];
  assign N95 = N184 & chosen_way_decode[0];
  assign N184 = decode_v_i[3] | decode_v_i[4];
  assign N96 = N185 & chosen_way_decode[0];
  assign N185 = decode_v_i[3] | decode_v_i[4];
  assign N97 = N186 & chosen_way_decode[1];
  assign N186 = decode_v_i[3] | decode_v_i[4];
  assign N98 = N187 & chosen_way_decode[1];
  assign N187 = decode_v_i[3] | decode_v_i[4];
  assign N99 = N188 & chosen_way_decode[2];
  assign N188 = decode_v_i[3] | decode_v_i[4];
  assign N100 = N189 & chosen_way_decode[2];
  assign N189 = decode_v_i[3] | decode_v_i[4];
  assign N101 = N190 & chosen_way_decode[3];
  assign N190 = decode_v_i[3] | decode_v_i[4];
  assign N102 = N191 & chosen_way_decode[3];
  assign N191 = decode_v_i[3] | decode_v_i[4];
  assign N103 = ~N93;
  assign N104 = ~N94;
  assign N105 = N103 & N104;
  assign N106 = N103 & N94;
  assign N107 = N93 & N104;
  assign N108 = N93 & N94;
  assign N111 = N193 & N110;
  assign N193 = N192 & N109;
  assign N192 = ~decode_v_i[3];
  assign N113 = ~dma_way_o[0];
  assign N114 = ~dma_way_o[1];
  assign N115 = N113 & N114;
  assign N116 = N113 & dma_way_o[1];
  assign N117 = dma_way_o[0] & N114;
  assign N118 = dma_way_o[0] & dma_way_o[1];
  assign N137 = ~dma_done_i;
  assign N138 = N113 & N114;
  assign N139 = N113 & dma_way_o[1];
  assign N140 = dma_way_o[0] & N114;
  assign N141 = dma_way_o[0] & dma_way_o[1];
  assign N160 = N194 | decode_v_i[5];
  assign N194 = decode_v_i[8] | decode_v_i[4];
  assign N162 = ~ack_i;
  assign N163 = ~tag_mem_data_o[79];
  assign N164 = N163;
  assign N165 = N46;
  assign N166 = N42;
  assign N167 = N163;
  assign N168 = ~goto_flush_op;
  assign N169 = goto_lock_op & N168;
  assign N170 = ~invalid_exist;
  assign N171 = N75 & N170;

  always @(posedge clk_i) begin
    if(reset_i) begin
      { dma_way_o[1:0] } <= { 1'b0, 1'b0 };
      { miss_state_r[3:0] } <= { 1'b0, 1'b0, 1'b0, 1'b0 };
    end else if(1'b1) begin
      { dma_way_o[1:0] } <= { chosen_way_o[1:0] };
      { miss_state_r[3:0] } <= { miss_state_n[3:0] };
    end 
  end


endmodule



module bsg_counter_clear_up_max_val_p4
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);

  output [2:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;
  reg [2:0] count_o;
  assign { N8, N7, N6 } = { N14, N13, N12 } + up_i;
  assign { N11, N10, N9 } = (N0)? { 1'b0, 1'b0, 1'b0 } : 
                            (N1)? { N8, N7, N6 } : 1'b0;
  assign N0 = reset_i;
  assign N1 = N2;
  assign { N14, N13, N12 } = count_o * N4;
  assign N2 = ~reset_i;
  assign N3 = N2;
  assign N4 = ~clear_i;
  assign N5 = N3 & N4;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { count_o[2:0] } <= { N11, N10, N9 };
    end 
  end


endmodule



module bsg_circular_ptr_slots_p4_max_add_p1
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [0:0] add_i;
  output [1:0] o;
  output [1:0] n_o;
  input clk;
  input reset_i;
  wire [1:0] n_o,genblk1_genblk1_ptr_r_p1;
  wire N0,N1,N2,N3,N4,N5,N6,N7;
  reg [1:0] o;
  assign genblk1_genblk1_ptr_r_p1 = o + 1'b1;
  assign { N6, N5 } = (N0)? { 1'b0, 1'b0 } : 
                      (N1)? n_o : 1'b0;
  assign N0 = reset_i;
  assign N1 = N4;
  assign n_o = (N2)? genblk1_genblk1_ptr_r_p1 : 
               (N3)? o : 1'b0;
  assign N2 = add_i[0];
  assign N3 = N7;
  assign N4 = ~reset_i;
  assign N7 = ~add_i[0];

  always @(posedge clk) begin
    if(1'b1) begin
      { o[1:0] } <= { N6, N5 };
    end 
  end


endmodule



module bsg_fifo_tracker_els_p4
(
  clk_i,
  reset_i,
  enq_i,
  deq_i,
  wptr_r_o,
  rptr_r_o,
  rptr_n_o,
  full_o,
  empty_o
);

  output [1:0] wptr_r_o;
  output [1:0] rptr_r_o;
  output [1:0] rptr_n_o;
  input clk_i;
  input reset_i;
  input enq_i;
  input deq_i;
  output full_o;
  output empty_o;
  wire [1:0] wptr_r_o,rptr_r_o,rptr_n_o;
  wire full_o,empty_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,equal_ptrs,SYNOPSYS_UNCONNECTED_1,
  SYNOPSYS_UNCONNECTED_2;
  reg deq_r,enq_r;

  bsg_circular_ptr_slots_p4_max_add_p1
  rptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(deq_i),
    .o(rptr_r_o),
    .n_o(rptr_n_o)
  );


  bsg_circular_ptr_slots_p4_max_add_p1
  wptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(enq_i),
    .o(wptr_r_o),
    .n_o({ SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2 })
  );

  assign equal_ptrs = rptr_r_o == wptr_r_o;
  assign N5 = (N0)? 1'b1 : 
              (N9)? 1'b1 : 
              (N4)? 1'b0 : 1'b0;
  assign N0 = N2;
  assign N6 = (N0)? 1'b0 : 
              (N9)? enq_i : 1'b0;
  assign N7 = (N0)? 1'b1 : 
              (N9)? deq_i : 1'b0;
  assign N1 = enq_i | deq_i;
  assign N2 = reset_i;
  assign N3 = N1 | N2;
  assign N4 = ~N3;
  assign N8 = ~N2;
  assign N9 = N1 & N8;
  assign empty_o = equal_ptrs & deq_r;
  assign full_o = equal_ptrs & enq_r;

  always @(posedge clk_i) begin
    if(N5) begin
      deq_r <= N7;
      enq_r <= N6;
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p32_els_p4_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [1:0] w_addr_i;
  input [31:0] w_data_i;
  input [1:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;
  reg [127:0] mem;
  assign r_data_o[31] = (N8)? mem[31] : 
                        (N10)? mem[63] : 
                        (N9)? mem[95] : 
                        (N11)? mem[127] : 1'b0;
  assign r_data_o[30] = (N8)? mem[30] : 
                        (N10)? mem[62] : 
                        (N9)? mem[94] : 
                        (N11)? mem[126] : 1'b0;
  assign r_data_o[29] = (N8)? mem[29] : 
                        (N10)? mem[61] : 
                        (N9)? mem[93] : 
                        (N11)? mem[125] : 1'b0;
  assign r_data_o[28] = (N8)? mem[28] : 
                        (N10)? mem[60] : 
                        (N9)? mem[92] : 
                        (N11)? mem[124] : 1'b0;
  assign r_data_o[27] = (N8)? mem[27] : 
                        (N10)? mem[59] : 
                        (N9)? mem[91] : 
                        (N11)? mem[123] : 1'b0;
  assign r_data_o[26] = (N8)? mem[26] : 
                        (N10)? mem[58] : 
                        (N9)? mem[90] : 
                        (N11)? mem[122] : 1'b0;
  assign r_data_o[25] = (N8)? mem[25] : 
                        (N10)? mem[57] : 
                        (N9)? mem[89] : 
                        (N11)? mem[121] : 1'b0;
  assign r_data_o[24] = (N8)? mem[24] : 
                        (N10)? mem[56] : 
                        (N9)? mem[88] : 
                        (N11)? mem[120] : 1'b0;
  assign r_data_o[23] = (N8)? mem[23] : 
                        (N10)? mem[55] : 
                        (N9)? mem[87] : 
                        (N11)? mem[119] : 1'b0;
  assign r_data_o[22] = (N8)? mem[22] : 
                        (N10)? mem[54] : 
                        (N9)? mem[86] : 
                        (N11)? mem[118] : 1'b0;
  assign r_data_o[21] = (N8)? mem[21] : 
                        (N10)? mem[53] : 
                        (N9)? mem[85] : 
                        (N11)? mem[117] : 1'b0;
  assign r_data_o[20] = (N8)? mem[20] : 
                        (N10)? mem[52] : 
                        (N9)? mem[84] : 
                        (N11)? mem[116] : 1'b0;
  assign r_data_o[19] = (N8)? mem[19] : 
                        (N10)? mem[51] : 
                        (N9)? mem[83] : 
                        (N11)? mem[115] : 1'b0;
  assign r_data_o[18] = (N8)? mem[18] : 
                        (N10)? mem[50] : 
                        (N9)? mem[82] : 
                        (N11)? mem[114] : 1'b0;
  assign r_data_o[17] = (N8)? mem[17] : 
                        (N10)? mem[49] : 
                        (N9)? mem[81] : 
                        (N11)? mem[113] : 1'b0;
  assign r_data_o[16] = (N8)? mem[16] : 
                        (N10)? mem[48] : 
                        (N9)? mem[80] : 
                        (N11)? mem[112] : 1'b0;
  assign r_data_o[15] = (N8)? mem[15] : 
                        (N10)? mem[47] : 
                        (N9)? mem[79] : 
                        (N11)? mem[111] : 1'b0;
  assign r_data_o[14] = (N8)? mem[14] : 
                        (N10)? mem[46] : 
                        (N9)? mem[78] : 
                        (N11)? mem[110] : 1'b0;
  assign r_data_o[13] = (N8)? mem[13] : 
                        (N10)? mem[45] : 
                        (N9)? mem[77] : 
                        (N11)? mem[109] : 1'b0;
  assign r_data_o[12] = (N8)? mem[12] : 
                        (N10)? mem[44] : 
                        (N9)? mem[76] : 
                        (N11)? mem[108] : 1'b0;
  assign r_data_o[11] = (N8)? mem[11] : 
                        (N10)? mem[43] : 
                        (N9)? mem[75] : 
                        (N11)? mem[107] : 1'b0;
  assign r_data_o[10] = (N8)? mem[10] : 
                        (N10)? mem[42] : 
                        (N9)? mem[74] : 
                        (N11)? mem[106] : 1'b0;
  assign r_data_o[9] = (N8)? mem[9] : 
                       (N10)? mem[41] : 
                       (N9)? mem[73] : 
                       (N11)? mem[105] : 1'b0;
  assign r_data_o[8] = (N8)? mem[8] : 
                       (N10)? mem[40] : 
                       (N9)? mem[72] : 
                       (N11)? mem[104] : 1'b0;
  assign r_data_o[7] = (N8)? mem[7] : 
                       (N10)? mem[39] : 
                       (N9)? mem[71] : 
                       (N11)? mem[103] : 1'b0;
  assign r_data_o[6] = (N8)? mem[6] : 
                       (N10)? mem[38] : 
                       (N9)? mem[70] : 
                       (N11)? mem[102] : 1'b0;
  assign r_data_o[5] = (N8)? mem[5] : 
                       (N10)? mem[37] : 
                       (N9)? mem[69] : 
                       (N11)? mem[101] : 1'b0;
  assign r_data_o[4] = (N8)? mem[4] : 
                       (N10)? mem[36] : 
                       (N9)? mem[68] : 
                       (N11)? mem[100] : 1'b0;
  assign r_data_o[3] = (N8)? mem[3] : 
                       (N10)? mem[35] : 
                       (N9)? mem[67] : 
                       (N11)? mem[99] : 1'b0;
  assign r_data_o[2] = (N8)? mem[2] : 
                       (N10)? mem[34] : 
                       (N9)? mem[66] : 
                       (N11)? mem[98] : 1'b0;
  assign r_data_o[1] = (N8)? mem[1] : 
                       (N10)? mem[33] : 
                       (N9)? mem[65] : 
                       (N11)? mem[97] : 1'b0;
  assign r_data_o[0] = (N8)? mem[0] : 
                       (N10)? mem[32] : 
                       (N9)? mem[64] : 
                       (N11)? mem[96] : 1'b0;
  assign N16 = w_addr_i[0] & w_addr_i[1];
  assign N15 = N0 & w_addr_i[1];
  assign N0 = ~w_addr_i[0];
  assign N14 = w_addr_i[0] & N1;
  assign N1 = ~w_addr_i[1];
  assign N13 = N2 & N3;
  assign N2 = ~w_addr_i[0];
  assign N3 = ~w_addr_i[1];
  assign { N20, N19, N18, N17 } = (N4)? { N16, N15, N14, N13 } : 
                                  (N5)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N4 = w_v_i;
  assign N5 = N12;
  assign N6 = ~r_addr_i[0];
  assign N7 = ~r_addr_i[1];
  assign N8 = N6 & N7;
  assign N9 = N6 & r_addr_i[1];
  assign N10 = r_addr_i[0] & N7;
  assign N11 = r_addr_i[0] & r_addr_i[1];
  assign N12 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N20) begin
      { mem[127:96] } <= { w_data_i[31:0] };
    end 
    if(N19) begin
      { mem[95:64] } <= { w_data_i[31:0] };
    end 
    if(N18) begin
      { mem[63:32] } <= { w_data_i[31:0] };
    end 
    if(N17) begin
      { mem[31:0] } <= { w_data_i[31:0] };
    end 
  end


endmodule



module bsg_mem_1r1w_width_p32_els_p4_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [1:0] w_addr_i;
  input [31:0] w_data_i;
  input [1:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;

  bsg_mem_1r1w_synth_width_p32_els_p4_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_fifo_1r1w_small_unhardened_width_p32_els_p4_ready_THEN_valid_p0
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,enque,full,empty,SYNOPSYS_UNCONNECTED_1,SYNOPSYS_UNCONNECTED_2;
  wire [1:0] wptr_r,rptr_r;

  bsg_fifo_tracker_els_p4
  ft
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .enq_i(enque),
    .deq_i(yumi_i),
    .wptr_r_o(wptr_r),
    .rptr_r_o(rptr_r),
    .rptr_n_o({ SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2 }),
    .full_o(full),
    .empty_o(empty)
  );


  bsg_mem_1r1w_width_p32_els_p4_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enque),
    .w_addr_i(wptr_r),
    .w_data_i(data_i),
    .r_v_i(v_o),
    .r_addr_i(rptr_r),
    .r_data_o(data_o)
  );

  assign enque = v_i & ready_o;
  assign ready_o = ~full;
  assign v_o = ~empty;

endmodule



module bsg_fifo_1r1w_small_width_p32_els_p4
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o;

  bsg_fifo_1r1w_small_unhardened_width_p32_els_p4_ready_THEN_valid_p0
  unhardened_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_o(ready_o),
    .data_i(data_i),
    .v_o(v_o),
    .data_o(data_o),
    .yumi_i(yumi_i)
  );


endmodule



module bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  reg [63:0] mem;
  assign r_data_o[31] = (N3)? mem[31] : 
                        (N0)? mem[63] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[30] = (N3)? mem[30] : 
                        (N0)? mem[62] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] : 
                        (N0)? mem[61] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] : 
                        (N0)? mem[60] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] : 
                        (N0)? mem[59] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] : 
                        (N0)? mem[58] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] : 
                        (N0)? mem[57] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] : 
                        (N0)? mem[56] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] : 
                        (N0)? mem[55] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] : 
                        (N0)? mem[54] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] : 
                        (N0)? mem[53] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] : 
                        (N0)? mem[52] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] : 
                        (N0)? mem[51] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] : 
                        (N0)? mem[50] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] : 
                        (N0)? mem[49] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] : 
                        (N0)? mem[48] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] : 
                        (N0)? mem[47] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] : 
                        (N0)? mem[46] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] : 
                        (N0)? mem[45] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] : 
                        (N0)? mem[44] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] : 
                        (N0)? mem[43] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] : 
                        (N0)? mem[42] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] : 
                       (N0)? mem[41] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] : 
                       (N0)? mem[40] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] : 
                       (N0)? mem[39] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] : 
                       (N0)? mem[38] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[37] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[36] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[35] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[34] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[33] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[32] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      { mem[63:32] } <= { w_data_i[31:0] };
    end 
    if(N7) begin
      { mem[31:0] } <= { w_data_i[31:0] };
    end 
  end


endmodule



module bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;

  bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p32
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 : 
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 : 
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 : 
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 : 
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 : 
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 : 
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end 
    if(N9) begin
      tail_r <= N10;
    end 
    if(N11) begin
      head_r <= N12;
    end 
  end


endmodule



module bsg_mux_width_p32_els_p4
(
  data_i,
  sel_i,
  data_o
);

  input [127:0] data_i;
  input [1:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[31] = (N2)? data_i[31] : 
                      (N4)? data_i[63] : 
                      (N3)? data_i[95] : 
                      (N5)? data_i[127] : 1'b0;
  assign data_o[30] = (N2)? data_i[30] : 
                      (N4)? data_i[62] : 
                      (N3)? data_i[94] : 
                      (N5)? data_i[126] : 1'b0;
  assign data_o[29] = (N2)? data_i[29] : 
                      (N4)? data_i[61] : 
                      (N3)? data_i[93] : 
                      (N5)? data_i[125] : 1'b0;
  assign data_o[28] = (N2)? data_i[28] : 
                      (N4)? data_i[60] : 
                      (N3)? data_i[92] : 
                      (N5)? data_i[124] : 1'b0;
  assign data_o[27] = (N2)? data_i[27] : 
                      (N4)? data_i[59] : 
                      (N3)? data_i[91] : 
                      (N5)? data_i[123] : 1'b0;
  assign data_o[26] = (N2)? data_i[26] : 
                      (N4)? data_i[58] : 
                      (N3)? data_i[90] : 
                      (N5)? data_i[122] : 1'b0;
  assign data_o[25] = (N2)? data_i[25] : 
                      (N4)? data_i[57] : 
                      (N3)? data_i[89] : 
                      (N5)? data_i[121] : 1'b0;
  assign data_o[24] = (N2)? data_i[24] : 
                      (N4)? data_i[56] : 
                      (N3)? data_i[88] : 
                      (N5)? data_i[120] : 1'b0;
  assign data_o[23] = (N2)? data_i[23] : 
                      (N4)? data_i[55] : 
                      (N3)? data_i[87] : 
                      (N5)? data_i[119] : 1'b0;
  assign data_o[22] = (N2)? data_i[22] : 
                      (N4)? data_i[54] : 
                      (N3)? data_i[86] : 
                      (N5)? data_i[118] : 1'b0;
  assign data_o[21] = (N2)? data_i[21] : 
                      (N4)? data_i[53] : 
                      (N3)? data_i[85] : 
                      (N5)? data_i[117] : 1'b0;
  assign data_o[20] = (N2)? data_i[20] : 
                      (N4)? data_i[52] : 
                      (N3)? data_i[84] : 
                      (N5)? data_i[116] : 1'b0;
  assign data_o[19] = (N2)? data_i[19] : 
                      (N4)? data_i[51] : 
                      (N3)? data_i[83] : 
                      (N5)? data_i[115] : 1'b0;
  assign data_o[18] = (N2)? data_i[18] : 
                      (N4)? data_i[50] : 
                      (N3)? data_i[82] : 
                      (N5)? data_i[114] : 1'b0;
  assign data_o[17] = (N2)? data_i[17] : 
                      (N4)? data_i[49] : 
                      (N3)? data_i[81] : 
                      (N5)? data_i[113] : 1'b0;
  assign data_o[16] = (N2)? data_i[16] : 
                      (N4)? data_i[48] : 
                      (N3)? data_i[80] : 
                      (N5)? data_i[112] : 1'b0;
  assign data_o[15] = (N2)? data_i[15] : 
                      (N4)? data_i[47] : 
                      (N3)? data_i[79] : 
                      (N5)? data_i[111] : 1'b0;
  assign data_o[14] = (N2)? data_i[14] : 
                      (N4)? data_i[46] : 
                      (N3)? data_i[78] : 
                      (N5)? data_i[110] : 1'b0;
  assign data_o[13] = (N2)? data_i[13] : 
                      (N4)? data_i[45] : 
                      (N3)? data_i[77] : 
                      (N5)? data_i[109] : 1'b0;
  assign data_o[12] = (N2)? data_i[12] : 
                      (N4)? data_i[44] : 
                      (N3)? data_i[76] : 
                      (N5)? data_i[108] : 1'b0;
  assign data_o[11] = (N2)? data_i[11] : 
                      (N4)? data_i[43] : 
                      (N3)? data_i[75] : 
                      (N5)? data_i[107] : 1'b0;
  assign data_o[10] = (N2)? data_i[10] : 
                      (N4)? data_i[42] : 
                      (N3)? data_i[74] : 
                      (N5)? data_i[106] : 1'b0;
  assign data_o[9] = (N2)? data_i[9] : 
                     (N4)? data_i[41] : 
                     (N3)? data_i[73] : 
                     (N5)? data_i[105] : 1'b0;
  assign data_o[8] = (N2)? data_i[8] : 
                     (N4)? data_i[40] : 
                     (N3)? data_i[72] : 
                     (N5)? data_i[104] : 1'b0;
  assign data_o[7] = (N2)? data_i[7] : 
                     (N4)? data_i[39] : 
                     (N3)? data_i[71] : 
                     (N5)? data_i[103] : 1'b0;
  assign data_o[6] = (N2)? data_i[6] : 
                     (N4)? data_i[38] : 
                     (N3)? data_i[70] : 
                     (N5)? data_i[102] : 1'b0;
  assign data_o[5] = (N2)? data_i[5] : 
                     (N4)? data_i[37] : 
                     (N3)? data_i[69] : 
                     (N5)? data_i[101] : 1'b0;
  assign data_o[4] = (N2)? data_i[4] : 
                     (N4)? data_i[36] : 
                     (N3)? data_i[68] : 
                     (N5)? data_i[100] : 1'b0;
  assign data_o[3] = (N2)? data_i[3] : 
                     (N4)? data_i[35] : 
                     (N3)? data_i[67] : 
                     (N5)? data_i[99] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] : 
                     (N4)? data_i[34] : 
                     (N3)? data_i[66] : 
                     (N5)? data_i[98] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N4)? data_i[33] : 
                     (N3)? data_i[65] : 
                     (N5)? data_i[97] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N4)? data_i[32] : 
                     (N3)? data_i[64] : 
                     (N5)? data_i[96] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_cache_dma_addr_width_p28_data_width_p32_block_size_in_words_p4_sets_p64_ways_p4_debug_p0
(
  clk_i,
  reset_i,
  dma_cmd_i,
  dma_way_i,
  dma_addr_i,
  done_o,
  snoop_word_o,
  dma_pkt_o,
  dma_pkt_v_o,
  dma_pkt_yumi_i,
  dma_data_i,
  dma_data_v_i,
  dma_data_ready_o,
  dma_data_o,
  dma_data_v_o,
  dma_data_yumi_i,
  data_mem_v_o,
  data_mem_w_o,
  data_mem_addr_o,
  data_mem_w_mask_o,
  data_mem_data_o,
  data_mem_data_i,
  dma_evict_o
);

  input [3:0] dma_cmd_i;
  input [1:0] dma_way_i;
  input [27:0] dma_addr_i;
  output [31:0] snoop_word_o;
  output [28:0] dma_pkt_o;
  input [31:0] dma_data_i;
  output [31:0] dma_data_o;
  output [7:0] data_mem_addr_o;
  output [15:0] data_mem_w_mask_o;
  output [127:0] data_mem_data_o;
  input [127:0] data_mem_data_i;
  input clk_i;
  input reset_i;
  input dma_pkt_yumi_i;
  input dma_data_v_i;
  input dma_data_yumi_i;
  output done_o;
  output dma_pkt_v_o;
  output dma_data_ready_o;
  output dma_data_v_o;
  output data_mem_v_o;
  output data_mem_w_o;
  output dma_evict_o;
  wire [28:0] dma_pkt_o;
  wire [31:0] dma_data_o,out_fifo_data_li;
  wire [7:0] data_mem_addr_o;
  wire [15:0] data_mem_w_mask_o;
  wire [127:0] data_mem_data_o;
  wire done_o,dma_pkt_v_o,dma_data_ready_o,dma_data_v_o,data_mem_v_o,data_mem_w_o,
  dma_evict_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,counter_clear,counter_up,in_fifo_v_lo,
  in_fifo_yumi_li,out_fifo_v_li,out_fifo_ready_lo,N11,N12,N13,N14,N15,N16,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,snoop_word_we,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,
  N75,N76;
  wire [2:2] counter_r;
  wire [1:0] dma_state_n;
  reg [31:0] snoop_word_o;
  reg [1:0] dma_state_r;
  assign dma_pkt_o[0] = 1'b0;
  assign dma_pkt_o[1] = 1'b0;
  assign dma_pkt_o[2] = 1'b0;
  assign dma_pkt_o[3] = 1'b0;
  assign dma_pkt_o[27] = dma_addr_i[27];
  assign dma_pkt_o[26] = dma_addr_i[26];
  assign dma_pkt_o[25] = dma_addr_i[25];
  assign dma_pkt_o[24] = dma_addr_i[24];
  assign dma_pkt_o[23] = dma_addr_i[23];
  assign dma_pkt_o[22] = dma_addr_i[22];
  assign dma_pkt_o[21] = dma_addr_i[21];
  assign dma_pkt_o[20] = dma_addr_i[20];
  assign dma_pkt_o[19] = dma_addr_i[19];
  assign dma_pkt_o[18] = dma_addr_i[18];
  assign dma_pkt_o[17] = dma_addr_i[17];
  assign dma_pkt_o[16] = dma_addr_i[16];
  assign dma_pkt_o[15] = dma_addr_i[15];
  assign dma_pkt_o[14] = dma_addr_i[14];
  assign dma_pkt_o[13] = dma_addr_i[13];
  assign dma_pkt_o[12] = dma_addr_i[12];
  assign dma_pkt_o[11] = dma_addr_i[11];
  assign dma_pkt_o[10] = dma_addr_i[10];
  assign dma_pkt_o[9] = dma_addr_i[9];
  assign data_mem_addr_o[7] = dma_addr_i[9];
  assign dma_pkt_o[8] = dma_addr_i[8];
  assign data_mem_addr_o[6] = dma_addr_i[8];
  assign dma_pkt_o[7] = dma_addr_i[7];
  assign data_mem_addr_o[5] = dma_addr_i[7];
  assign dma_pkt_o[6] = dma_addr_i[6];
  assign data_mem_addr_o[4] = dma_addr_i[6];
  assign dma_pkt_o[5] = dma_addr_i[5];
  assign data_mem_addr_o[3] = dma_addr_i[5];
  assign dma_pkt_o[4] = dma_addr_i[4];
  assign data_mem_addr_o[2] = dma_addr_i[4];
  assign data_mem_w_mask_o[12] = data_mem_w_mask_o[15];
  assign data_mem_w_mask_o[13] = data_mem_w_mask_o[15];
  assign data_mem_w_mask_o[14] = data_mem_w_mask_o[15];
  assign data_mem_w_mask_o[8] = data_mem_w_mask_o[11];
  assign data_mem_w_mask_o[9] = data_mem_w_mask_o[11];
  assign data_mem_w_mask_o[10] = data_mem_w_mask_o[11];
  assign data_mem_w_mask_o[4] = data_mem_w_mask_o[7];
  assign data_mem_w_mask_o[5] = data_mem_w_mask_o[7];
  assign data_mem_w_mask_o[6] = data_mem_w_mask_o[7];
  assign data_mem_w_mask_o[0] = data_mem_w_mask_o[3];
  assign data_mem_w_mask_o[1] = data_mem_w_mask_o[3];
  assign data_mem_w_mask_o[2] = data_mem_w_mask_o[3];
  assign data_mem_data_o[31] = data_mem_data_o[127];
  assign data_mem_data_o[63] = data_mem_data_o[127];
  assign data_mem_data_o[95] = data_mem_data_o[127];
  assign data_mem_data_o[30] = data_mem_data_o[126];
  assign data_mem_data_o[62] = data_mem_data_o[126];
  assign data_mem_data_o[94] = data_mem_data_o[126];
  assign data_mem_data_o[29] = data_mem_data_o[125];
  assign data_mem_data_o[61] = data_mem_data_o[125];
  assign data_mem_data_o[93] = data_mem_data_o[125];
  assign data_mem_data_o[28] = data_mem_data_o[124];
  assign data_mem_data_o[60] = data_mem_data_o[124];
  assign data_mem_data_o[92] = data_mem_data_o[124];
  assign data_mem_data_o[27] = data_mem_data_o[123];
  assign data_mem_data_o[59] = data_mem_data_o[123];
  assign data_mem_data_o[91] = data_mem_data_o[123];
  assign data_mem_data_o[26] = data_mem_data_o[122];
  assign data_mem_data_o[58] = data_mem_data_o[122];
  assign data_mem_data_o[90] = data_mem_data_o[122];
  assign data_mem_data_o[25] = data_mem_data_o[121];
  assign data_mem_data_o[57] = data_mem_data_o[121];
  assign data_mem_data_o[89] = data_mem_data_o[121];
  assign data_mem_data_o[24] = data_mem_data_o[120];
  assign data_mem_data_o[56] = data_mem_data_o[120];
  assign data_mem_data_o[88] = data_mem_data_o[120];
  assign data_mem_data_o[23] = data_mem_data_o[119];
  assign data_mem_data_o[55] = data_mem_data_o[119];
  assign data_mem_data_o[87] = data_mem_data_o[119];
  assign data_mem_data_o[22] = data_mem_data_o[118];
  assign data_mem_data_o[54] = data_mem_data_o[118];
  assign data_mem_data_o[86] = data_mem_data_o[118];
  assign data_mem_data_o[21] = data_mem_data_o[117];
  assign data_mem_data_o[53] = data_mem_data_o[117];
  assign data_mem_data_o[85] = data_mem_data_o[117];
  assign data_mem_data_o[20] = data_mem_data_o[116];
  assign data_mem_data_o[52] = data_mem_data_o[116];
  assign data_mem_data_o[84] = data_mem_data_o[116];
  assign data_mem_data_o[19] = data_mem_data_o[115];
  assign data_mem_data_o[51] = data_mem_data_o[115];
  assign data_mem_data_o[83] = data_mem_data_o[115];
  assign data_mem_data_o[18] = data_mem_data_o[114];
  assign data_mem_data_o[50] = data_mem_data_o[114];
  assign data_mem_data_o[82] = data_mem_data_o[114];
  assign data_mem_data_o[17] = data_mem_data_o[113];
  assign data_mem_data_o[49] = data_mem_data_o[113];
  assign data_mem_data_o[81] = data_mem_data_o[113];
  assign data_mem_data_o[16] = data_mem_data_o[112];
  assign data_mem_data_o[48] = data_mem_data_o[112];
  assign data_mem_data_o[80] = data_mem_data_o[112];
  assign data_mem_data_o[15] = data_mem_data_o[111];
  assign data_mem_data_o[47] = data_mem_data_o[111];
  assign data_mem_data_o[79] = data_mem_data_o[111];
  assign data_mem_data_o[14] = data_mem_data_o[110];
  assign data_mem_data_o[46] = data_mem_data_o[110];
  assign data_mem_data_o[78] = data_mem_data_o[110];
  assign data_mem_data_o[13] = data_mem_data_o[109];
  assign data_mem_data_o[45] = data_mem_data_o[109];
  assign data_mem_data_o[77] = data_mem_data_o[109];
  assign data_mem_data_o[12] = data_mem_data_o[108];
  assign data_mem_data_o[44] = data_mem_data_o[108];
  assign data_mem_data_o[76] = data_mem_data_o[108];
  assign data_mem_data_o[11] = data_mem_data_o[107];
  assign data_mem_data_o[43] = data_mem_data_o[107];
  assign data_mem_data_o[75] = data_mem_data_o[107];
  assign data_mem_data_o[10] = data_mem_data_o[106];
  assign data_mem_data_o[42] = data_mem_data_o[106];
  assign data_mem_data_o[74] = data_mem_data_o[106];
  assign data_mem_data_o[9] = data_mem_data_o[105];
  assign data_mem_data_o[41] = data_mem_data_o[105];
  assign data_mem_data_o[73] = data_mem_data_o[105];
  assign data_mem_data_o[8] = data_mem_data_o[104];
  assign data_mem_data_o[40] = data_mem_data_o[104];
  assign data_mem_data_o[72] = data_mem_data_o[104];
  assign data_mem_data_o[7] = data_mem_data_o[103];
  assign data_mem_data_o[39] = data_mem_data_o[103];
  assign data_mem_data_o[71] = data_mem_data_o[103];
  assign data_mem_data_o[6] = data_mem_data_o[102];
  assign data_mem_data_o[38] = data_mem_data_o[102];
  assign data_mem_data_o[70] = data_mem_data_o[102];
  assign data_mem_data_o[5] = data_mem_data_o[101];
  assign data_mem_data_o[37] = data_mem_data_o[101];
  assign data_mem_data_o[69] = data_mem_data_o[101];
  assign data_mem_data_o[4] = data_mem_data_o[100];
  assign data_mem_data_o[36] = data_mem_data_o[100];
  assign data_mem_data_o[68] = data_mem_data_o[100];
  assign data_mem_data_o[3] = data_mem_data_o[99];
  assign data_mem_data_o[35] = data_mem_data_o[99];
  assign data_mem_data_o[67] = data_mem_data_o[99];
  assign data_mem_data_o[2] = data_mem_data_o[98];
  assign data_mem_data_o[34] = data_mem_data_o[98];
  assign data_mem_data_o[66] = data_mem_data_o[98];
  assign data_mem_data_o[1] = data_mem_data_o[97];
  assign data_mem_data_o[33] = data_mem_data_o[97];
  assign data_mem_data_o[65] = data_mem_data_o[97];
  assign data_mem_data_o[0] = data_mem_data_o[96];
  assign data_mem_data_o[32] = data_mem_data_o[96];
  assign data_mem_data_o[64] = data_mem_data_o[96];

  bsg_counter_clear_up_max_val_p4
  dma_counter
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(counter_clear),
    .up_i(counter_up),
    .count_o({ counter_r[2:2], data_mem_addr_o[1:0] })
  );


  bsg_fifo_1r1w_small_width_p32_els_p4
  in_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(dma_data_v_i),
    .ready_o(dma_data_ready_o),
    .data_i(dma_data_i),
    .v_o(in_fifo_v_lo),
    .data_o(data_mem_data_o[127:96]),
    .yumi_i(in_fifo_yumi_li)
  );


  bsg_two_fifo_width_p32
  out_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(out_fifo_ready_lo),
    .data_i(out_fifo_data_li),
    .v_i(out_fifo_v_li),
    .v_o(dma_data_v_o),
    .data_o(dma_data_o),
    .yumi_i(dma_data_yumi_i)
  );


  bsg_decode_num_out_p4
  dma_way_demux
  (
    .i(dma_way_i),
    .o({ data_mem_w_mask_o[15:15], data_mem_w_mask_o[11:11], data_mem_w_mask_o[7:7], data_mem_w_mask_o[3:3] })
  );


  bsg_mux_width_p32_els_p4
  write_data_mux
  (
    .data_i(data_mem_data_i),
    .sel_i(dma_way_i),
    .data_o(out_fifo_data_li)
  );

  assign N12 = N11 & N64;
  assign N13 = dma_state_r[1] | N64;
  assign N15 = N11 | dma_state_r[0];
  assign N17 = dma_state_r[1] & dma_state_r[0];
  assign N18 = dma_cmd_i[1] | N35;
  assign N19 = N21 | N18;
  assign N21 = dma_cmd_i[3] | dma_cmd_i[2];
  assign N22 = N34 | dma_cmd_i[0];
  assign N23 = N21 | N22;
  assign N25 = dma_cmd_i[3] | N33;
  assign N26 = N25 | N29;
  assign N28 = N32 | dma_cmd_i[2];
  assign N29 = dma_cmd_i[1] | dma_cmd_i[0];
  assign N30 = N28 | N29;
  assign N36 = N32 & N33;
  assign N37 = N34 & N35;
  assign N38 = N36 & N37;
  assign N60 = dma_addr_i[3:2] == data_mem_addr_o[1:0];
  assign N64 = ~dma_state_r[0];
  assign N65 = N64 | dma_state_r[1];
  assign N66 = ~N65;
  assign N67 = ~counter_r[2];
  assign N68 = data_mem_addr_o[1] | N67;
  assign N69 = data_mem_addr_o[0] | N68;
  assign N70 = ~N69;
  assign N71 = ~data_mem_addr_o[1];
  assign N72 = ~data_mem_addr_o[0];
  assign N73 = N71 | counter_r[2];
  assign N74 = N72 | N73;
  assign N75 = ~N74;
  assign N44 = (N0)? 1'b1 : 
               (N1)? 1'b1 : 
               (N2)? 1'b0 : 
               (N3)? 1'b0 : 
               (N4)? 1'b0 : 
               (N43)? 1'b0 : 1'b0;
  assign N0 = N20;
  assign N1 = N24;
  assign N2 = N27;
  assign N3 = N31;
  assign N4 = N38;
  assign N45 = (N0)? 1'b0 : 
               (N1)? 1'b1 : 
               (N2)? 1'b0 : 
               (N3)? 1'b0 : 
               (N4)? 1'b0 : 
               (N43)? 1'b0 : 1'b0;
  assign N46 = (N0)? dma_pkt_yumi_i : 
               (N1)? dma_pkt_yumi_i : 
               (N2)? 1'b0 : 
               (N3)? 1'b0 : 
               (N4)? 1'b0 : 
               (N43)? 1'b0 : 1'b0;
  assign N47 = (N0)? 1'b0 : 
               (N1)? 1'b0 : 
               (N2)? 1'b1 : 
               (N3)? 1'b1 : 
               (N4)? 1'b0 : 
               (N43)? 1'b0 : 1'b0;
  assign N48 = (N0)? 1'b0 : 
               (N1)? 1'b0 : 
               (N2)? 1'b0 : 
               (N3)? 1'b1 : 
               (N4)? 1'b0 : 
               (N43)? 1'b0 : 1'b0;
  assign N50 = ~N49;
  assign N55 = ~N54;
  assign counter_clear = (N5)? N47 : 
                         (N6)? N52 : 
                         (N7)? N57 : 
                         (N8)? 1'b0 : 1'b0;
  assign N5 = N12;
  assign N6 = N14;
  assign N7 = N16;
  assign N8 = N17;
  assign counter_up = (N5)? N48 : 
                      (N6)? N51 : 
                      (N7)? N56 : 
                      (N8)? 1'b0 : 1'b0;
  assign data_mem_v_o = (N5)? N48 : 
                        (N6)? in_fifo_v_lo : 
                        (N7)? N58 : 
                        (N8)? 1'b0 : 1'b0;
  assign dma_pkt_v_o = (N5)? N44 : 
                       (N6)? 1'b0 : 
                       (N7)? 1'b0 : 
                       (N8)? 1'b0 : 1'b0;
  assign dma_pkt_o[28] = (N5)? N45 : 
                         (N6)? 1'b0 : 
                         (N7)? 1'b0 : 
                         (N8)? 1'b0 : 1'b0;
  assign done_o = (N5)? N46 : 
                  (N6)? N53 : 
                  (N7)? N59 : 
                  (N8)? 1'b0 : 1'b0;
  assign dma_state_n = (N5)? { N31, N27 } : 
                       (N6)? { 1'b0, N50 } : 
                       (N7)? { N55, 1'b0 } : 
                       (N8)? { 1'b0, 1'b0 } : 1'b0;
  assign data_mem_w_o = (N5)? 1'b0 : 
                        (N6)? in_fifo_v_lo : 
                        (N7)? 1'b0 : 
                        (N8)? 1'b0 : 1'b0;
  assign in_fifo_yumi_li = (N5)? 1'b0 : 
                           (N6)? in_fifo_v_lo : 
                           (N7)? 1'b0 : 
                           (N8)? 1'b0 : 1'b0;
  assign out_fifo_v_li = (N5)? 1'b0 : 
                         (N6)? 1'b0 : 
                         (N7)? 1'b1 : 
                         (N8)? 1'b0 : 1'b0;
  assign dma_evict_o = (N5)? 1'b0 : 
                       (N6)? 1'b0 : 
                       (N7)? 1'b1 : 
                       (N8)? 1'b0 : 1'b0;
  assign N63 = (N9)? 1'b0 : 
               (N10)? snoop_word_we : 1'b0;
  assign N9 = N62;
  assign N10 = N61;
  assign N11 = ~dma_state_r[1];
  assign N14 = ~N13;
  assign N16 = ~N15;
  assign N20 = ~N19;
  assign N24 = ~N23;
  assign N27 = ~N26;
  assign N31 = ~N30;
  assign N32 = ~dma_cmd_i[3];
  assign N33 = ~dma_cmd_i[2];
  assign N34 = ~dma_cmd_i[1];
  assign N35 = ~dma_cmd_i[0];
  assign N39 = N24 | N20;
  assign N40 = N27 | N39;
  assign N41 = N31 | N40;
  assign N42 = N38 | N41;
  assign N43 = ~N42;
  assign N49 = N75 & in_fifo_v_lo;
  assign N51 = in_fifo_v_lo & N74;
  assign N52 = in_fifo_v_lo & N75;
  assign N53 = N75 & in_fifo_v_lo;
  assign N54 = N70 & out_fifo_ready_lo;
  assign N56 = out_fifo_ready_lo & N69;
  assign N57 = out_fifo_ready_lo & N70;
  assign N58 = out_fifo_ready_lo & N69;
  assign N59 = N70 & out_fifo_ready_lo;
  assign snoop_word_we = N76 & in_fifo_v_lo;
  assign N76 = N66 & N60;
  assign N61 = ~reset_i;
  assign N62 = reset_i;

  always @(posedge clk_i) begin
    if(N63) begin
      { snoop_word_o[31:0] } <= { data_mem_data_o[127:96] };
    end 
    if(reset_i) begin
      { dma_state_r[1:0] } <= { 1'b0, 1'b0 };
    end else if(1'b1) begin
      { dma_state_r[1:0] } <= { dma_state_n[1:0] };
    end 
  end


endmodule



module bsg_cache_sbuf_queue_width_p66
(
  clk_i,
  data_i,
  el0_en_i,
  el1_en_i,
  mux0_sel_i,
  mux1_sel_i,
  el0_snoop_o,
  el1_snoop_o,
  data_o
);

  input [65:0] data_i;
  output [65:0] el0_snoop_o;
  output [65:0] el1_snoop_o;
  output [65:0] data_o;
  input clk_i;
  input el0_en_i;
  input el1_en_i;
  input mux0_sel_i;
  input mux1_sel_i;
  wire [65:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71;
  reg [65:0] el0_snoop_o,el1_snoop_o;
  assign { N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5 } = (N0)? el0_snoop_o : 
                                                                                                                                                                                                                                                                                                                                                   (N1)? data_i : 1'b0;
  assign N0 = mux0_sel_i;
  assign N1 = N4;
  assign data_o = (N2)? el1_snoop_o : 
                  (N3)? data_i : 1'b0;
  assign N2 = mux1_sel_i;
  assign N3 = N71;
  assign N4 = ~mux0_sel_i;
  assign N71 = ~mux1_sel_i;

  always @(posedge clk_i) begin
    if(el0_en_i) begin
      { el0_snoop_o[65:0] } <= { data_i[65:0] };
    end 
    if(el1_en_i) begin
      { el1_snoop_o[65:0] } <= { N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5 };
    end 
  end


endmodule



module bsg_mux_segmented_segments_p4_segment_width_p8
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [31:0] data0_i;
  input [31:0] data1_i;
  input [3:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7;
  assign data_o[7:0] = (N0)? data1_i[7:0] : 
                       (N4)? data0_i[7:0] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[15:8] = (N1)? data1_i[15:8] : 
                        (N5)? data0_i[15:8] : 1'b0;
  assign N1 = sel_i[1];
  assign data_o[23:16] = (N2)? data1_i[23:16] : 
                         (N6)? data0_i[23:16] : 1'b0;
  assign N2 = sel_i[2];
  assign data_o[31:24] = (N3)? data1_i[31:24] : 
                         (N7)? data0_i[31:24] : 1'b0;
  assign N3 = sel_i[3];
  assign N4 = ~sel_i[0];
  assign N5 = ~sel_i[1];
  assign N6 = ~sel_i[2];
  assign N7 = ~sel_i[3];

endmodule



module bsg_cache_sbuf_data_width_p32_addr_width_p28_ways_p4
(
  clk_i,
  reset_i,
  sbuf_entry_i,
  v_i,
  sbuf_entry_o,
  v_o,
  yumi_i,
  empty_o,
  bypass_addr_i,
  bypass_v_i,
  bypass_data_o,
  bypass_mask_o
);

  input [65:0] sbuf_entry_i;
  output [65:0] sbuf_entry_o;
  input [27:0] bypass_addr_i;
  output [31:0] bypass_data_o;
  output [3:0] bypass_mask_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  input bypass_v_i;
  output v_o;
  output empty_o;
  wire [65:0] sbuf_entry_o,el0,el1;
  wire v_o,empty_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,el0_valid,el1_valid,
  el0_enable,N14,el1_enable,mux0_sel,mux1_sel,N15,N16,N17,N18,N19,N20,N21,N22,N23,
  N24,N25,tag_hit0_n,tag_hit1_n,tag_hit2_n,n_2_net__3_,n_2_net__2_,n_2_net__1_,
  n_2_net__0_,n_4_net__3_,n_4_net__2_,n_4_net__1_,n_4_net__0_,N26,N27,N28,N29,N30,N31,
  N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,
  N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,
  N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83;
  wire [3:3] tag_hit0x4,tag_hit1x4,tag_hit2x4;
  wire [3:0] bypass_mask_n;
  wire [31:0] el0or1_data,bypass_data_n;
  reg [1:0] num_els_r;
  reg [31:0] bypass_data_o;
  reg [3:0] bypass_mask_o;
  assign N8 = N6 & N7;
  assign N9 = num_els_r[1] | N7;
  assign N11 = N6 | num_els_r[0];
  assign N13 = num_els_r[1] & num_els_r[0];

  bsg_cache_sbuf_queue_width_p66
  sbq
  (
    .clk_i(clk_i),
    .data_i(sbuf_entry_i),
    .el0_en_i(el0_enable),
    .el1_en_i(el1_enable),
    .mux0_sel_i(mux0_sel),
    .mux1_sel_i(mux1_sel),
    .el0_snoop_o(el0),
    .el1_snoop_o(el1),
    .data_o(sbuf_entry_o)
  );

  assign tag_hit0_n = bypass_addr_i[27:2] == el0[65:40];
  assign tag_hit1_n = bypass_addr_i[27:2] == el1[65:40];
  assign tag_hit2_n = bypass_addr_i[27:2] == sbuf_entry_i[65:40];

  bsg_mux_segmented_segments_p4_segment_width_p8
  mux_segmented_merge0
  (
    .data0_i(el1[37:6]),
    .data1_i(el0[37:6]),
    .sel_i({ n_2_net__3_, n_2_net__2_, n_2_net__1_, n_2_net__0_ }),
    .data_o(el0or1_data)
  );


  bsg_mux_segmented_segments_p4_segment_width_p8
  mux_segmented_merge1
  (
    .data0_i(el0or1_data),
    .data1_i(sbuf_entry_i[37:6]),
    .sel_i({ n_4_net__3_, n_4_net__2_, n_4_net__1_, n_4_net__0_ }),
    .data_o(bypass_data_n)
  );

  assign { N20, N19 } = num_els_r + v_i;
  assign { N23, N22 } = { N20, N19 } - N21;
  assign v_o = (N0)? v_i : 
               (N1)? 1'b1 : 
               (N2)? 1'b1 : 
               (N3)? 1'b0 : 1'b0;
  assign N0 = N8;
  assign N1 = N10;
  assign N2 = N12;
  assign N3 = N13;
  assign empty_o = (N0)? 1'b1 : 
                   (N1)? 1'b0 : 
                   (N2)? 1'b0 : 
                   (N3)? 1'b0 : 1'b0;
  assign el0_valid = (N0)? 1'b0 : 
                     (N1)? 1'b0 : 
                     (N2)? 1'b1 : 
                     (N3)? 1'b0 : 1'b0;
  assign el1_valid = (N0)? 1'b0 : 
                     (N1)? 1'b1 : 
                     (N2)? 1'b1 : 
                     (N3)? 1'b0 : 1'b0;
  assign el0_enable = (N0)? 1'b0 : 
                      (N1)? N15 : 
                      (N2)? N17 : 
                      (N3)? 1'b0 : 1'b0;
  assign el1_enable = (N0)? N14 : 
                      (N1)? N16 : 
                      (N2)? yumi_i : 
                      (N3)? 1'b0 : 1'b0;
  assign mux0_sel = (N0)? 1'b0 : 
                    (N1)? 1'b0 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b0 : 1'b0;
  assign mux1_sel = (N0)? 1'b0 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b0 : 1'b0;
  assign { N25, N24 } = (N4)? { 1'b0, 1'b0 } : 
                        (N5)? { N23, N22 } : 1'b0;
  assign N4 = reset_i;
  assign N5 = N18;
  assign N28 = (N4)? 1'b1 : 
               (N66)? 1'b1 : 
               (N27)? 1'b0 : 1'b0;
  assign { N32, N31, N30, N29 } = (N4)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N66)? bypass_mask_n : 1'b0;
  assign { N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33 } = (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                              (N66)? bypass_data_n : 1'b0;
  assign N6 = ~num_els_r[1];
  assign N7 = ~num_els_r[0];
  assign N10 = ~N9;
  assign N12 = ~N11;
  assign N14 = v_i & N67;
  assign N67 = ~yumi_i;
  assign N15 = v_i & N67;
  assign N16 = v_i & yumi_i;
  assign N17 = v_i & yumi_i;
  assign N18 = ~reset_i;
  assign N21 = v_o & yumi_i;
  assign tag_hit0x4[3] = tag_hit0_n & el0_valid;
  assign tag_hit1x4[3] = tag_hit1_n & el1_valid;
  assign tag_hit2x4[3] = tag_hit2_n & v_i;
  assign bypass_mask_n[3] = N70 | N71;
  assign N70 = N68 | N69;
  assign N68 = tag_hit0x4[3] & el0[5];
  assign N69 = tag_hit1x4[3] & el1[5];
  assign N71 = tag_hit2x4[3] & sbuf_entry_i[5];
  assign bypass_mask_n[2] = N74 | N75;
  assign N74 = N72 | N73;
  assign N72 = tag_hit0x4[3] & el0[4];
  assign N73 = tag_hit1x4[3] & el1[4];
  assign N75 = tag_hit2x4[3] & sbuf_entry_i[4];
  assign bypass_mask_n[1] = N78 | N79;
  assign N78 = N76 | N77;
  assign N76 = tag_hit0x4[3] & el0[3];
  assign N77 = tag_hit1x4[3] & el1[3];
  assign N79 = tag_hit2x4[3] & sbuf_entry_i[3];
  assign bypass_mask_n[0] = N82 | N83;
  assign N82 = N80 | N81;
  assign N80 = tag_hit0x4[3] & el0[2];
  assign N81 = tag_hit1x4[3] & el1[2];
  assign N83 = tag_hit2x4[3] & sbuf_entry_i[2];
  assign n_2_net__3_ = tag_hit0x4[3] & el0[5];
  assign n_2_net__2_ = tag_hit0x4[3] & el0[4];
  assign n_2_net__1_ = tag_hit0x4[3] & el0[3];
  assign n_2_net__0_ = tag_hit0x4[3] & el0[2];
  assign n_4_net__3_ = tag_hit2x4[3] & sbuf_entry_i[5];
  assign n_4_net__2_ = tag_hit2x4[3] & sbuf_entry_i[4];
  assign n_4_net__1_ = tag_hit2x4[3] & sbuf_entry_i[3];
  assign n_4_net__0_ = tag_hit2x4[3] & sbuf_entry_i[2];
  assign N26 = bypass_v_i | reset_i;
  assign N27 = ~N26;
  assign N65 = ~reset_i;
  assign N66 = bypass_v_i & N65;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { num_els_r[1:0] } <= { N25, N24 };
    end 
    if(N28) begin
      { bypass_data_o[31:0] } <= { N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33 };
      { bypass_mask_o[3:0] } <= { N32, N31, N30, N29 };
    end 
  end


endmodule



module bsg_mux_width_p32_els_p3
(
  data_i,
  sel_i,
  data_o
);

  input [95:0] data_i;
  input [1:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign N5 = N0 & N1;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign data_o[31] = (N2)? data_i[31] : 
                      (N3)? data_i[63] : 
                      (N4)? data_i[95] : 1'b0;
  assign N2 = N5;
  assign N3 = sel_i[0];
  assign N4 = sel_i[1];
  assign data_o[30] = (N2)? data_i[30] : 
                      (N3)? data_i[62] : 
                      (N4)? data_i[94] : 1'b0;
  assign data_o[29] = (N2)? data_i[29] : 
                      (N3)? data_i[61] : 
                      (N4)? data_i[93] : 1'b0;
  assign data_o[28] = (N2)? data_i[28] : 
                      (N3)? data_i[60] : 
                      (N4)? data_i[92] : 1'b0;
  assign data_o[27] = (N2)? data_i[27] : 
                      (N3)? data_i[59] : 
                      (N4)? data_i[91] : 1'b0;
  assign data_o[26] = (N2)? data_i[26] : 
                      (N3)? data_i[58] : 
                      (N4)? data_i[90] : 1'b0;
  assign data_o[25] = (N2)? data_i[25] : 
                      (N3)? data_i[57] : 
                      (N4)? data_i[89] : 1'b0;
  assign data_o[24] = (N2)? data_i[24] : 
                      (N3)? data_i[56] : 
                      (N4)? data_i[88] : 1'b0;
  assign data_o[23] = (N2)? data_i[23] : 
                      (N3)? data_i[55] : 
                      (N4)? data_i[87] : 1'b0;
  assign data_o[22] = (N2)? data_i[22] : 
                      (N3)? data_i[54] : 
                      (N4)? data_i[86] : 1'b0;
  assign data_o[21] = (N2)? data_i[21] : 
                      (N3)? data_i[53] : 
                      (N4)? data_i[85] : 1'b0;
  assign data_o[20] = (N2)? data_i[20] : 
                      (N3)? data_i[52] : 
                      (N4)? data_i[84] : 1'b0;
  assign data_o[19] = (N2)? data_i[19] : 
                      (N3)? data_i[51] : 
                      (N4)? data_i[83] : 1'b0;
  assign data_o[18] = (N2)? data_i[18] : 
                      (N3)? data_i[50] : 
                      (N4)? data_i[82] : 1'b0;
  assign data_o[17] = (N2)? data_i[17] : 
                      (N3)? data_i[49] : 
                      (N4)? data_i[81] : 1'b0;
  assign data_o[16] = (N2)? data_i[16] : 
                      (N3)? data_i[48] : 
                      (N4)? data_i[80] : 1'b0;
  assign data_o[15] = (N2)? data_i[15] : 
                      (N3)? data_i[47] : 
                      (N4)? data_i[79] : 1'b0;
  assign data_o[14] = (N2)? data_i[14] : 
                      (N3)? data_i[46] : 
                      (N4)? data_i[78] : 1'b0;
  assign data_o[13] = (N2)? data_i[13] : 
                      (N3)? data_i[45] : 
                      (N4)? data_i[77] : 1'b0;
  assign data_o[12] = (N2)? data_i[12] : 
                      (N3)? data_i[44] : 
                      (N4)? data_i[76] : 1'b0;
  assign data_o[11] = (N2)? data_i[11] : 
                      (N3)? data_i[43] : 
                      (N4)? data_i[75] : 1'b0;
  assign data_o[10] = (N2)? data_i[10] : 
                      (N3)? data_i[42] : 
                      (N4)? data_i[74] : 1'b0;
  assign data_o[9] = (N2)? data_i[9] : 
                     (N3)? data_i[41] : 
                     (N4)? data_i[73] : 1'b0;
  assign data_o[8] = (N2)? data_i[8] : 
                     (N3)? data_i[40] : 
                     (N4)? data_i[72] : 1'b0;
  assign data_o[7] = (N2)? data_i[7] : 
                     (N3)? data_i[39] : 
                     (N4)? data_i[71] : 1'b0;
  assign data_o[6] = (N2)? data_i[6] : 
                     (N3)? data_i[38] : 
                     (N4)? data_i[70] : 1'b0;
  assign data_o[5] = (N2)? data_i[5] : 
                     (N3)? data_i[37] : 
                     (N4)? data_i[69] : 1'b0;
  assign data_o[4] = (N2)? data_i[4] : 
                     (N3)? data_i[36] : 
                     (N4)? data_i[68] : 1'b0;
  assign data_o[3] = (N2)? data_i[3] : 
                     (N3)? data_i[35] : 
                     (N4)? data_i[67] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] : 
                     (N3)? data_i[34] : 
                     (N4)? data_i[66] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N3)? data_i[33] : 
                     (N4)? data_i[65] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N3)? data_i[32] : 
                     (N4)? data_i[64] : 1'b0;

endmodule



module bsg_mux_width_p4_els_p3
(
  data_i,
  sel_i,
  data_o
);

  input [11:0] data_i;
  input [1:0] sel_i;
  output [3:0] data_o;
  wire [3:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign N5 = N0 & N1;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign data_o[3] = (N2)? data_i[3] : 
                     (N3)? data_i[7] : 
                     (N4)? data_i[11] : 1'b0;
  assign N2 = N5;
  assign N3 = sel_i[0];
  assign N4 = sel_i[1];
  assign data_o[2] = (N2)? data_i[2] : 
                     (N3)? data_i[6] : 
                     (N4)? data_i[10] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N3)? data_i[5] : 
                     (N4)? data_i[9] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N3)? data_i[4] : 
                     (N4)? data_i[8] : 1'b0;

endmodule



module bsg_decode_num_out_p2
(
  i,
  o
);

  input [0:0] i;
  output [1:0] o;
  wire [1:0] o;
  assign o = { 1'b0, 1'b1 } << i[0];

endmodule



module bsg_mux_width_p8_els_p4
(
  data_i,
  sel_i,
  data_o
);

  input [31:0] data_i;
  input [1:0] sel_i;
  output [7:0] data_o;
  wire [7:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[7] = (N2)? data_i[7] : 
                     (N4)? data_i[15] : 
                     (N3)? data_i[23] : 
                     (N5)? data_i[31] : 1'b0;
  assign data_o[6] = (N2)? data_i[6] : 
                     (N4)? data_i[14] : 
                     (N3)? data_i[22] : 
                     (N5)? data_i[30] : 1'b0;
  assign data_o[5] = (N2)? data_i[5] : 
                     (N4)? data_i[13] : 
                     (N3)? data_i[21] : 
                     (N5)? data_i[29] : 1'b0;
  assign data_o[4] = (N2)? data_i[4] : 
                     (N4)? data_i[12] : 
                     (N3)? data_i[20] : 
                     (N5)? data_i[28] : 1'b0;
  assign data_o[3] = (N2)? data_i[3] : 
                     (N4)? data_i[11] : 
                     (N3)? data_i[19] : 
                     (N5)? data_i[27] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] : 
                     (N4)? data_i[10] : 
                     (N3)? data_i[18] : 
                     (N5)? data_i[26] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N4)? data_i[9] : 
                     (N3)? data_i[17] : 
                     (N5)? data_i[25] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N4)? data_i[8] : 
                     (N3)? data_i[16] : 
                     (N5)? data_i[24] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_mux_width_p16_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [31:0] data_i;
  input [0:0] sel_i;
  output [15:0] data_o;
  wire [15:0] data_o;
  wire N0,N1;
  assign data_o[15] = (N1)? data_i[15] : 
                      (N0)? data_i[31] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[14] = (N1)? data_i[14] : 
                      (N0)? data_i[30] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] : 
                      (N0)? data_i[29] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] : 
                      (N0)? data_i[28] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] : 
                      (N0)? data_i[27] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] : 
                      (N0)? data_i[26] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] : 
                     (N0)? data_i[25] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] : 
                     (N0)? data_i[24] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] : 
                     (N0)? data_i[23] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] : 
                     (N0)? data_i[22] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] : 
                     (N0)? data_i[21] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] : 
                     (N0)? data_i[20] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[19] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[18] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[17] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[16] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module bsg_cache
(
  clk_i,
  reset_i,
  cache_pkt_i,
  v_i,
  ready_o,
  data_o,
  v_o,
  yumi_i,
  dma_pkt_o,
  dma_pkt_v_o,
  dma_pkt_yumi_i,
  dma_data_i,
  dma_data_v_i,
  dma_data_ready_o,
  dma_data_o,
  dma_data_v_o,
  dma_data_yumi_i,
  v_we_o
);

  input [68:0] cache_pkt_i;
  output [31:0] data_o;
  output [28:0] dma_pkt_o;
  input [31:0] dma_data_i;
  output [31:0] dma_data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  input dma_pkt_yumi_i;
  input dma_data_v_i;
  input dma_data_yumi_i;
  output ready_o;
  output v_o;
  output dma_pkt_v_o;
  output dma_data_ready_o;
  output dma_data_v_o;
  output v_we_o;
  wire [31:0] data_o,dma_data_o,snoop_word_lo,bypass_data_lo,sbuf_data_in,ld_data_way_picked,
  bypass_data_masked,snoop_or_ld_data,expanded_mask_v,ld_data_masked,
  ld_data_final_lo;
  wire [28:0] dma_pkt_o;
  wire ready_o,v_o,dma_pkt_v_o,dma_data_ready_o,dma_data_v_o,v_we_o,N0,N1,N2,N3,N4,N5,
  N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,
  N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,
  N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
  N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,
  N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,
  N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,
  tag_mem_v_li,tag_mem_w_li,data_mem_v_li,data_mem_w_li,N121,N122,N123,N124,N125,N126,
  N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,
  N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,
  N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,
  N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,
  N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
  N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,
  N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,
  N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,
  N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,
  N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,tag_hit_found,ld_st_miss,N297,
  N298,N299,N300,N301,N302,N303,tagfl_hit,aflinv_hit,N304,N305,N306,N307,N308,
  N309,N310,N311,N312,N313,N314,alock_miss,N315,N316,N317,N318,N319,N320,N321,N322,
  N323,N324,aunlock_hit,miss_v,retval_op_v,stat_mem_v_li,stat_mem_w_li,sbuf_empty_li,
  dma_done_li,miss_stat_mem_v_lo,miss_stat_mem_w_lo,miss_tag_mem_v_lo,
  miss_tag_mem_w_lo,recover_lo,miss_done_lo,n_0_net_,dma_data_mem_v_lo,dma_data_mem_w_lo,
  dma_evict_lo,sbuf_entry_li_data__31_,sbuf_entry_li_data__30_,sbuf_entry_li_data__29_,
  sbuf_entry_li_data__28_,sbuf_entry_li_data__27_,sbuf_entry_li_data__26_,
  sbuf_entry_li_data__25_,sbuf_entry_li_data__24_,sbuf_entry_li_data__23_,
  sbuf_entry_li_data__22_,sbuf_entry_li_data__21_,sbuf_entry_li_data__20_,sbuf_entry_li_data__19_,
  sbuf_entry_li_data__18_,sbuf_entry_li_data__17_,sbuf_entry_li_data__16_,
  sbuf_entry_li_data__15_,sbuf_entry_li_data__14_,sbuf_entry_li_data__13_,
  sbuf_entry_li_data__12_,sbuf_entry_li_data__11_,sbuf_entry_li_data__10_,sbuf_entry_li_data__9_,
  sbuf_entry_li_data__8_,sbuf_entry_li_data__7_,sbuf_entry_li_data__6_,
  sbuf_entry_li_data__5_,sbuf_entry_li_data__4_,sbuf_entry_li_data__3_,sbuf_entry_li_data__2_,
  sbuf_entry_li_data__1_,sbuf_entry_li_data__0_,sbuf_entry_li_mask__3_,
  sbuf_entry_li_mask__2_,sbuf_entry_li_mask__1_,sbuf_entry_li_mask__0_,
  sbuf_entry_li_way_id__1_,sbuf_entry_li_way_id__0_,sbuf_v_li,sbuf_v_lo,sbuf_yumi_li,bypass_v_li,
  sbuf_mask_in_mux_li_1__3_,sbuf_mask_in_mux_li_1__2_,sbuf_mask_in_mux_li_1__1_,
  sbuf_mask_in_mux_li_1__0_,sbuf_mask_in_mux_li_0__3_,sbuf_mask_in_mux_li_0__2_,
  sbuf_mask_in_mux_li_0__1_,sbuf_mask_in_mux_li_0__0_,N325,N326,N327,N328,N329,N330,
  ld_data_final_li_1__31_,ld_data_final_li_1__30_,ld_data_final_li_1__29_,
  ld_data_final_li_1__28_,ld_data_final_li_1__27_,ld_data_final_li_1__26_,ld_data_final_li_1__25_,
  ld_data_final_li_1__24_,ld_data_final_li_1__23_,ld_data_final_li_1__22_,
  ld_data_final_li_1__21_,ld_data_final_li_1__20_,ld_data_final_li_1__19_,
  ld_data_final_li_1__18_,ld_data_final_li_1__17_,ld_data_final_li_1__16_,ld_data_final_li_0__31_,
  ld_data_final_li_0__30_,ld_data_final_li_0__29_,ld_data_final_li_0__28_,
  ld_data_final_li_0__27_,ld_data_final_li_0__26_,ld_data_final_li_0__25_,
  ld_data_final_li_0__24_,ld_data_final_li_0__23_,ld_data_final_li_0__22_,ld_data_final_li_0__21_,
  ld_data_final_li_0__20_,ld_data_final_li_0__19_,ld_data_final_li_0__18_,
  ld_data_final_li_0__17_,ld_data_final_li_0__16_,ld_data_final_li_0__15_,
  ld_data_final_li_0__14_,ld_data_final_li_0__13_,ld_data_final_li_0__12_,ld_data_final_li_0__11_,
  ld_data_final_li_0__10_,ld_data_final_li_0__9_,ld_data_final_li_0__8_,N331,N332,
  N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
  N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,
  N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,
  N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,
  N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,
  N413,N414,N415,N416,N417,N418,N419,N420,tl_ready,N421,N422,tagst_write_en,N423,
  N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,
  N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,
  N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,
  N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,
  N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,
  N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
  N520,N521;
  wire [15:0] decode,data_mem_w_mask_li,dma_data_mem_w_mask_lo,sbuf_data_mem_w_mask,
  ld_data_sel_1__non_max_size_byte_sel;
  wire [5:0] tag_mem_addr_li,stat_mem_addr_li,miss_stat_mem_addr_lo,miss_tag_mem_addr_lo;
  wire [79:0] tag_mem_data_li,tag_mem_w_mask_li,tag_mem_data_lo,miss_tag_mem_data_lo,
  miss_tag_mem_w_mask_lo;
  wire [7:0] data_mem_addr_li,dma_data_mem_addr_lo,ld_data_sel_0__non_max_size_byte_sel;
  wire [127:0] data_mem_data_li,data_mem_data_lo,dma_data_mem_data_lo;
  wire [3:0] tag_hit_v,dma_cmd_lo,bypass_mask_lo,sbuf_way_decode,sbuf_mask_in,
  sbuf_in_sel_0__non_max_size_decode_lo,addr_way_decode;
  wire [1:0] tag_hit_way_id,dma_way_lo,chosen_way_lo,sbuf_in_sel_1__non_max_size_decode_lo;
  wire [6:0] stat_mem_data_li,stat_mem_w_mask_li,stat_mem_data_lo,miss_stat_mem_data_lo,
  miss_stat_mem_w_mask_lo;
  wire [27:0] dma_addr_lo;
  wire [65:0] sbuf_entry_lo;
  wire [2:0] plru_decode_data_lo,plru_decode_mask_lo;
  reg [31:0] data_tl_r,data_v_r;
  reg v_tl_r,v_v_r;
  reg [15:0] decode_tl_r,decode_v_r;
  reg [3:0] mask_tl_r,mask_v_r,valid_v_r,lock_v_r;
  reg [27:0] addr_tl_r,addr_v_r;
  reg [127:0] ld_data_v_r;
  reg [71:0] tag_v_r;

  bsg_cache_pkt_decode_data_width_p32_addr_width_p28
  cache_pkt_decoder
  (
    .cache_pkt_i(cache_pkt_i),
    .decode_o(decode)
  );


  bsg_mem_1rw_sync_mask_write_bit_width_p80_els_p64_latch_last_read_p1
  tag_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(tag_mem_data_li),
    .addr_i(tag_mem_addr_li),
    .v_i(tag_mem_v_li),
    .w_mask_i(tag_mem_w_mask_li),
    .w_i(tag_mem_w_li),
    .data_o(tag_mem_data_lo)
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p256_data_width_p128_latch_last_read_p1
  data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li),
    .data_i(data_mem_data_li),
    .write_mask_i(data_mem_w_mask_li),
    .data_o(data_mem_data_lo)
  );

  assign N293 = addr_v_r[27:10] == tag_v_r[17:0];
  assign N294 = addr_v_r[27:10] == tag_v_r[35:18];
  assign N295 = addr_v_r[27:10] == tag_v_r[53:36];
  assign N296 = addr_v_r[27:10] == tag_v_r[71:54];

  bsg_priority_encode_width_p4_lo_to_hi_p1
  tag_hit_pe
  (
    .i(tag_hit_v),
    .addr_o(tag_hit_way_id),
    .v_o(tag_hit_found)
  );

  assign N303 = (N299)? valid_v_r[0] : 
                (N301)? valid_v_r[1] : 
                (N300)? valid_v_r[2] : 
                (N302)? valid_v_r[3] : 1'b0;
  assign N312 = (N308)? lock_v_r[0] : 
                (N310)? lock_v_r[1] : 
                (N309)? lock_v_r[2] : 
                (N311)? lock_v_r[3] : 1'b0;
  assign N323 = (N319)? lock_v_r[0] : 
                (N321)? lock_v_r[1] : 
                (N320)? lock_v_r[2] : 
                (N322)? lock_v_r[3] : 1'b0;

  bsg_mem_1rw_sync_mask_write_bit_width_p7_els_p64_latch_last_read_p1
  stat_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(stat_mem_data_li),
    .addr_i(stat_mem_addr_li),
    .v_i(stat_mem_v_li),
    .w_mask_i(stat_mem_w_mask_li),
    .w_i(stat_mem_w_li),
    .data_o(stat_mem_data_lo)
  );


  bsg_cache_miss_addr_width_p28_data_width_p32_block_size_in_words_p4_sets_p64_ways_p4
  miss
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .miss_v_i(miss_v),
    .decode_v_i(decode_v_r),
    .addr_v_i(addr_v_r),
    .tag_v_i(tag_v_r),
    .valid_v_i(valid_v_r),
    .lock_v_i(lock_v_r),
    .tag_hit_way_id_i(tag_hit_way_id),
    .tag_hit_found_i(tag_hit_found),
    .sbuf_empty_i(sbuf_empty_li),
    .dma_cmd_o(dma_cmd_lo),
    .dma_way_o(dma_way_lo),
    .dma_addr_o(dma_addr_lo),
    .dma_done_i(dma_done_li),
    .stat_info_i(stat_mem_data_lo),
    .stat_mem_v_o(miss_stat_mem_v_lo),
    .stat_mem_w_o(miss_stat_mem_w_lo),
    .stat_mem_addr_o(miss_stat_mem_addr_lo),
    .stat_mem_data_o(miss_stat_mem_data_lo),
    .stat_mem_w_mask_o(miss_stat_mem_w_mask_lo),
    .tag_mem_v_o(miss_tag_mem_v_lo),
    .tag_mem_w_o(miss_tag_mem_w_lo),
    .tag_mem_addr_o(miss_tag_mem_addr_lo),
    .tag_mem_data_o(miss_tag_mem_data_lo),
    .tag_mem_w_mask_o(miss_tag_mem_w_mask_lo),
    .done_o(miss_done_lo),
    .recover_o(recover_lo),
    .chosen_way_o(chosen_way_lo),
    .ack_i(n_0_net_)
  );


  bsg_cache_dma_addr_width_p28_data_width_p32_block_size_in_words_p4_sets_p64_ways_p4_debug_p0
  dma
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .dma_cmd_i(dma_cmd_lo),
    .dma_way_i(dma_way_lo),
    .dma_addr_i(dma_addr_lo),
    .done_o(dma_done_li),
    .snoop_word_o(snoop_word_lo),
    .dma_pkt_o(dma_pkt_o),
    .dma_pkt_v_o(dma_pkt_v_o),
    .dma_pkt_yumi_i(dma_pkt_yumi_i),
    .dma_data_i(dma_data_i),
    .dma_data_v_i(dma_data_v_i),
    .dma_data_ready_o(dma_data_ready_o),
    .dma_data_o(dma_data_o),
    .dma_data_v_o(dma_data_v_o),
    .dma_data_yumi_i(dma_data_yumi_i),
    .data_mem_v_o(dma_data_mem_v_lo),
    .data_mem_w_o(dma_data_mem_w_lo),
    .data_mem_addr_o(dma_data_mem_addr_lo),
    .data_mem_w_mask_o(dma_data_mem_w_mask_lo),
    .data_mem_data_o(dma_data_mem_data_lo),
    .data_mem_data_i(data_mem_data_lo),
    .dma_evict_o(dma_evict_lo)
  );


  bsg_cache_sbuf_data_width_p32_addr_width_p28_ways_p4
  sbuf
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .sbuf_entry_i({ addr_v_r, sbuf_entry_li_data__31_, sbuf_entry_li_data__30_, sbuf_entry_li_data__29_, sbuf_entry_li_data__28_, sbuf_entry_li_data__27_, sbuf_entry_li_data__26_, sbuf_entry_li_data__25_, sbuf_entry_li_data__24_, sbuf_entry_li_data__23_, sbuf_entry_li_data__22_, sbuf_entry_li_data__21_, sbuf_entry_li_data__20_, sbuf_entry_li_data__19_, sbuf_entry_li_data__18_, sbuf_entry_li_data__17_, sbuf_entry_li_data__16_, sbuf_entry_li_data__15_, sbuf_entry_li_data__14_, sbuf_entry_li_data__13_, sbuf_entry_li_data__12_, sbuf_entry_li_data__11_, sbuf_entry_li_data__10_, sbuf_entry_li_data__9_, sbuf_entry_li_data__8_, sbuf_entry_li_data__7_, sbuf_entry_li_data__6_, sbuf_entry_li_data__5_, sbuf_entry_li_data__4_, sbuf_entry_li_data__3_, sbuf_entry_li_data__2_, sbuf_entry_li_data__1_, sbuf_entry_li_data__0_, sbuf_entry_li_mask__3_, sbuf_entry_li_mask__2_, sbuf_entry_li_mask__1_, sbuf_entry_li_mask__0_, sbuf_entry_li_way_id__1_, sbuf_entry_li_way_id__0_ }),
    .v_i(sbuf_v_li),
    .sbuf_entry_o(sbuf_entry_lo),
    .v_o(sbuf_v_lo),
    .yumi_i(sbuf_yumi_li),
    .empty_o(sbuf_empty_li),
    .bypass_addr_i(addr_tl_r),
    .bypass_v_i(bypass_v_li),
    .bypass_data_o(bypass_data_lo),
    .bypass_mask_o(bypass_mask_lo)
  );


  bsg_decode_num_out_p4
  sbuf_way_demux
  (
    .i(sbuf_entry_lo[1:0]),
    .o(sbuf_way_decode)
  );


  bsg_mux_width_p32_els_p3
  sbuf_data_in_mux
  (
    .data_i({ data_v_r, data_v_r[15:0], data_v_r[15:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0] }),
    .sel_i(decode_v_r[15:14]),
    .data_o(sbuf_data_in)
  );


  bsg_mux_width_p4_els_p3
  sbuf_mask_in_mux
  (
    .data_i({ 1'b1, 1'b1, 1'b1, 1'b1, sbuf_mask_in_mux_li_1__3_, sbuf_mask_in_mux_li_1__2_, sbuf_mask_in_mux_li_1__1_, sbuf_mask_in_mux_li_1__0_, sbuf_mask_in_mux_li_0__3_, sbuf_mask_in_mux_li_0__2_, sbuf_mask_in_mux_li_0__1_, sbuf_mask_in_mux_li_0__0_ }),
    .sel_i(decode_v_r[15:14]),
    .data_o(sbuf_mask_in)
  );


  bsg_decode_num_out_p4
  sbuf_in_sel_0__non_max_size_dec
  (
    .i(addr_v_r[1:0]),
    .o(sbuf_in_sel_0__non_max_size_decode_lo)
  );


  bsg_expand_bitmask
  sbuf_in_sel_0__non_max_size_exp
  (
    .i(sbuf_in_sel_0__non_max_size_decode_lo),
    .o({ sbuf_mask_in_mux_li_0__3_, sbuf_mask_in_mux_li_0__2_, sbuf_mask_in_mux_li_0__1_, sbuf_mask_in_mux_li_0__0_ })
  );


  bsg_decode_num_out_p2
  sbuf_in_sel_1__non_max_size_dec
  (
    .i(addr_v_r[1]),
    .o(sbuf_in_sel_1__non_max_size_decode_lo)
  );


  bsg_expand_bitmask
  sbuf_in_sel_1__non_max_size_exp
  (
    .i(sbuf_in_sel_1__non_max_size_decode_lo),
    .o({ sbuf_mask_in_mux_li_1__3_, sbuf_mask_in_mux_li_1__2_, sbuf_mask_in_mux_li_1__1_, sbuf_mask_in_mux_li_1__0_ })
  );


  bsg_mux_width_p32_els_p4
  ld_data_mux
  (
    .data_i(ld_data_v_r),
    .sel_i(tag_hit_way_id),
    .data_o(ld_data_way_picked)
  );


  bsg_mux_segmented_segments_p4_segment_width_p8
  bypass_mux_segmented
  (
    .data0_i(ld_data_way_picked),
    .data1_i(bypass_data_lo),
    .sel_i(bypass_mask_lo),
    .data_o(bypass_data_masked)
  );


  bsg_expand_bitmask
  mask_v_expand
  (
    .i(mask_v_r),
    .o(expanded_mask_v)
  );


  bsg_mux_width_p8_els_p4
  ld_data_sel_0__non_max_size_byte_mux
  (
    .data_i(snoop_or_ld_data),
    .sel_i(addr_v_r[1:0]),
    .data_o(ld_data_sel_0__non_max_size_byte_sel)
  );


  bsg_mux_width_p16_els_p2
  ld_data_sel_1__non_max_size_byte_mux
  (
    .data_i(snoop_or_ld_data),
    .sel_i(addr_v_r[1]),
    .data_o(ld_data_sel_1__non_max_size_byte_sel)
  );


  bsg_mux_width_p32_els_p3
  ld_data_size_mux
  (
    .data_i({ snoop_or_ld_data, ld_data_final_li_1__31_, ld_data_final_li_1__30_, ld_data_final_li_1__29_, ld_data_final_li_1__28_, ld_data_final_li_1__27_, ld_data_final_li_1__26_, ld_data_final_li_1__25_, ld_data_final_li_1__24_, ld_data_final_li_1__23_, ld_data_final_li_1__22_, ld_data_final_li_1__21_, ld_data_final_li_1__20_, ld_data_final_li_1__19_, ld_data_final_li_1__18_, ld_data_final_li_1__17_, ld_data_final_li_1__16_, ld_data_sel_1__non_max_size_byte_sel, ld_data_final_li_0__31_, ld_data_final_li_0__30_, ld_data_final_li_0__29_, ld_data_final_li_0__28_, ld_data_final_li_0__27_, ld_data_final_li_0__26_, ld_data_final_li_0__25_, ld_data_final_li_0__24_, ld_data_final_li_0__23_, ld_data_final_li_0__22_, ld_data_final_li_0__21_, ld_data_final_li_0__20_, ld_data_final_li_0__19_, ld_data_final_li_0__18_, ld_data_final_li_0__17_, ld_data_final_li_0__16_, ld_data_final_li_0__15_, ld_data_final_li_0__14_, ld_data_final_li_0__13_, ld_data_final_li_0__12_, ld_data_final_li_0__11_, ld_data_final_li_0__10_, ld_data_final_li_0__9_, ld_data_final_li_0__8_, ld_data_sel_0__non_max_size_byte_sel }),
    .sel_i(decode_v_r[15:14]),
    .data_o(ld_data_final_lo)
  );

  assign N344 = (N340)? lock_v_r[0] : 
                (N342)? lock_v_r[1] : 
                (N341)? lock_v_r[2] : 
                (N343)? lock_v_r[3] : 1'b0;
  assign N351 = (N347)? valid_v_r[0] : 
                (N349)? valid_v_r[1] : 
                (N348)? valid_v_r[2] : 
                (N350)? valid_v_r[3] : 1'b0;
  assign N358 = (N354)? tag_v_r[17] : 
                (N356)? tag_v_r[35] : 
                (N355)? tag_v_r[53] : 
                (N357)? tag_v_r[71] : 1'b0;
  assign N359 = (N354)? tag_v_r[16] : 
                (N356)? tag_v_r[34] : 
                (N355)? tag_v_r[52] : 
                (N357)? tag_v_r[70] : 1'b0;
  assign N360 = (N354)? tag_v_r[15] : 
                (N356)? tag_v_r[33] : 
                (N355)? tag_v_r[51] : 
                (N357)? tag_v_r[69] : 1'b0;
  assign N361 = (N354)? tag_v_r[14] : 
                (N356)? tag_v_r[32] : 
                (N355)? tag_v_r[50] : 
                (N357)? tag_v_r[68] : 1'b0;
  assign N362 = (N354)? tag_v_r[13] : 
                (N356)? tag_v_r[31] : 
                (N355)? tag_v_r[49] : 
                (N357)? tag_v_r[67] : 1'b0;
  assign N363 = (N354)? tag_v_r[12] : 
                (N356)? tag_v_r[30] : 
                (N355)? tag_v_r[48] : 
                (N357)? tag_v_r[66] : 1'b0;
  assign N364 = (N354)? tag_v_r[11] : 
                (N356)? tag_v_r[29] : 
                (N355)? tag_v_r[47] : 
                (N357)? tag_v_r[65] : 1'b0;
  assign N365 = (N354)? tag_v_r[10] : 
                (N356)? tag_v_r[28] : 
                (N355)? tag_v_r[46] : 
                (N357)? tag_v_r[64] : 1'b0;
  assign N366 = (N354)? tag_v_r[9] : 
                (N356)? tag_v_r[27] : 
                (N355)? tag_v_r[45] : 
                (N357)? tag_v_r[63] : 1'b0;
  assign N367 = (N354)? tag_v_r[8] : 
                (N356)? tag_v_r[26] : 
                (N355)? tag_v_r[44] : 
                (N357)? tag_v_r[62] : 1'b0;
  assign N368 = (N354)? tag_v_r[7] : 
                (N356)? tag_v_r[25] : 
                (N355)? tag_v_r[43] : 
                (N357)? tag_v_r[61] : 1'b0;
  assign N369 = (N354)? tag_v_r[6] : 
                (N356)? tag_v_r[24] : 
                (N355)? tag_v_r[42] : 
                (N357)? tag_v_r[60] : 1'b0;
  assign N370 = (N354)? tag_v_r[5] : 
                (N356)? tag_v_r[23] : 
                (N355)? tag_v_r[41] : 
                (N357)? tag_v_r[59] : 1'b0;
  assign N371 = (N354)? tag_v_r[4] : 
                (N356)? tag_v_r[22] : 
                (N355)? tag_v_r[40] : 
                (N357)? tag_v_r[58] : 1'b0;
  assign N372 = (N354)? tag_v_r[3] : 
                (N356)? tag_v_r[21] : 
                (N355)? tag_v_r[39] : 
                (N357)? tag_v_r[57] : 1'b0;
  assign N373 = (N354)? tag_v_r[2] : 
                (N356)? tag_v_r[20] : 
                (N355)? tag_v_r[38] : 
                (N357)? tag_v_r[56] : 1'b0;
  assign N374 = (N354)? tag_v_r[1] : 
                (N356)? tag_v_r[19] : 
                (N355)? tag_v_r[37] : 
                (N357)? tag_v_r[55] : 1'b0;
  assign N375 = (N354)? tag_v_r[0] : 
                (N356)? tag_v_r[18] : 
                (N355)? tag_v_r[36] : 
                (N357)? tag_v_r[54] : 1'b0;

  bsg_decode_num_out_p4
  addr_way_demux
  (
    .i(cache_pkt_i[47:46]),
    .o(addr_way_decode)
  );


  bsg_lru_pseudo_tree_decode_ways_p4
  plru_decode
  (
    .way_id_i(tag_hit_way_id),
    .data_o(plru_decode_data_lo),
    .mask_o(plru_decode_mask_lo)
  );

  assign N36 = (N0)? 1'b1 : 
               (N120)? 1'b1 : 
               (N35)? 1'b0 : 1'b0;
  assign N0 = N33;
  assign N37 = (N0)? 1'b0 : 
               (N120)? v_i : 1'b0;
  assign N38 = (N0)? 1'b1 : 
               (N120)? v_i : 
               (N35)? 1'b0 : 1'b0;
  assign { N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                              (N120)? decode : 1'b0;
  assign { N58, N57, N56, N55 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N120)? cache_pkt_i[3:0] : 1'b0;
  assign { N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                          (N120)? cache_pkt_i[63:36] : 1'b0;
  assign { N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                 (N120)? cache_pkt_i[35:4] : 1'b0;
  assign N124 = (N1)? 1'b1 : 
                (N292)? 1'b1 : 
                (N123)? 1'b0 : 1'b0;
  assign N1 = N121;
  assign N125 = (N1)? 1'b0 : 
                (N292)? v_tl_r : 1'b0;
  assign { N133, N126 } = (N1)? { 1'b1, 1'b1 } : 
                          (N292)? { v_tl_r, v_tl_r } : 
                          (N123)? { 1'b0, 1'b0 } : 1'b0;
  assign { N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N132, N131, N130, N129, N128, N127 } = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N292)? { tag_mem_data_lo[77:60], tag_mem_data_lo[57:40], tag_mem_data_lo[37:20], tag_mem_data_lo[17:0] } : 1'b0;
  assign N200 = (N1)? 1'b1 : 
                (N292)? v_tl_r : 
                (N123)? 1'b0 : 1'b0;
  assign { N204, N203, N202, N201 } = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N292)? mask_tl_r : 1'b0;
  assign { N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205 } = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                              (N292)? decode_tl_r : 1'b0;
  assign { N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221 } = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                      (N292)? addr_tl_r : 1'b0;
  assign { N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249 } = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                              (N292)? data_tl_r : 1'b0;
  assign { N284, N283, N282, N281 } = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N292)? { tag_mem_data_lo[79:79], tag_mem_data_lo[59:59], tag_mem_data_lo[39:39], tag_mem_data_lo[19:19] } : 1'b0;
  assign { N288, N287, N286, N285 } = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N292)? { tag_mem_data_lo[78:78], tag_mem_data_lo[58:58], tag_mem_data_lo[38:38], tag_mem_data_lo[18:18] } : 1'b0;
  assign { N290, N289 } = (N1)? { 1'b0, 1'b0 } : 
                          (N292)? { v_tl_r, v_tl_r } : 
                          (N123)? { 1'b0, 1'b0 } : 1'b0;
  assign N314 = (N2)? N313 : 
                (N3)? 1'b1 : 1'b0;
  assign N2 = N305;
  assign N3 = N304;
  assign N324 = (N4)? N323 : 
                (N5)? 1'b0 : 1'b0;
  assign N4 = N316;
  assign N5 = N315;
  assign { sbuf_entry_li_data__31_, sbuf_entry_li_data__30_, sbuf_entry_li_data__29_, sbuf_entry_li_data__28_, sbuf_entry_li_data__27_, sbuf_entry_li_data__26_, sbuf_entry_li_data__25_, sbuf_entry_li_data__24_, sbuf_entry_li_data__23_, sbuf_entry_li_data__22_, sbuf_entry_li_data__21_, sbuf_entry_li_data__20_, sbuf_entry_li_data__19_, sbuf_entry_li_data__18_, sbuf_entry_li_data__17_, sbuf_entry_li_data__16_, sbuf_entry_li_data__15_, sbuf_entry_li_data__14_, sbuf_entry_li_data__13_, sbuf_entry_li_data__12_, sbuf_entry_li_data__11_, sbuf_entry_li_data__10_, sbuf_entry_li_data__9_, sbuf_entry_li_data__8_, sbuf_entry_li_data__7_, sbuf_entry_li_data__6_, sbuf_entry_li_data__5_, sbuf_entry_li_data__4_, sbuf_entry_li_data__3_, sbuf_entry_li_data__2_, sbuf_entry_li_data__1_, sbuf_entry_li_data__0_ } = (N6)? data_v_r : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N326)? sbuf_data_in : 1'b0;
  assign N6 = N325;
  assign { sbuf_entry_li_mask__3_, sbuf_entry_li_mask__2_, sbuf_entry_li_mask__1_, sbuf_entry_li_mask__0_ } = (N7)? mask_v_r : 
                                                                                                              (N328)? sbuf_mask_in : 1'b0;
  assign N7 = N327;
  assign snoop_or_ld_data = (N8)? snoop_word_lo : 
                            (N9)? bypass_data_masked : 1'b0;
  assign N8 = N330;
  assign N9 = N329;
  assign { N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376 } = (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N344, N351 } : 
                                                                                                                                                                                                              (N409)? { 1'b0, 1'b0, 1'b0, 1'b0, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, addr_v_r[9:4], 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                              (N412)? ld_data_masked : 
                                                                                                                                                                                                              (N337)? ld_data_final_lo : 1'b0;
  assign N10 = N332;
  assign data_o = (N11)? { N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376 } : 
                  (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = retval_op_v;
  assign N12 = N331;
  assign N415 = (N13)? miss_done_lo : 
                (N14)? 1'b1 : 1'b0;
  assign N13 = N414;
  assign N14 = N413;
  assign v_we_o = (N15)? N417 : 
                  (N16)? 1'b1 : 1'b0;
  assign N15 = v_v_r;
  assign N16 = N416;
  assign tl_ready = (N17)? N420 : 
                    (N18)? 1'b1 : 1'b0;
  assign N17 = N419;
  assign N18 = N418;
  assign ready_o = (N19)? N422 : 
                   (N20)? tl_ready : 1'b0;
  assign N19 = v_tl_r;
  assign N20 = N421;
  assign tag_mem_w_li = (N21)? miss_tag_mem_w_lo : 
                        (N22)? tagst_write_en : 1'b0;
  assign N21 = N424;
  assign N22 = N423;
  assign { N434, N433, N432, N431, N430, N429 } = (N23)? addr_tl_r[9:4] : 
                                                  (N436)? miss_tag_mem_addr_lo : 
                                                  (N428)? cache_pkt_i[45:40] : 1'b0;
  assign N23 = recover_lo;
  assign tag_mem_addr_li = (N24)? { N434, N433, N432, N431, N430, N429 } : 
                           (N25)? cache_pkt_i[45:40] : 1'b0;
  assign N24 = N426;
  assign N25 = N425;
  assign tag_mem_data_li = (N24)? miss_tag_mem_data_lo : 
                           (N25)? { cache_pkt_i[35:34], cache_pkt_i[21:4], cache_pkt_i[35:34], cache_pkt_i[21:4], cache_pkt_i[35:34], cache_pkt_i[21:4], cache_pkt_i[35:34], cache_pkt_i[21:4] } : 1'b0;
  assign tag_mem_w_mask_li = (N24)? miss_tag_mem_w_mask_lo : 
                             (N25)? { addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0] } : 1'b0;
  assign data_mem_data_li = (N26)? dma_data_mem_data_lo : 
                            (N27)? { sbuf_entry_lo[37:6], sbuf_entry_lo[37:6], sbuf_entry_lo[37:6], sbuf_entry_lo[37:6] } : 1'b0;
  assign N26 = dma_data_mem_w_lo;
  assign N27 = N437;
  assign data_mem_addr_li = (N23)? addr_tl_r[9:2] : 
                            (N442)? dma_data_mem_addr_lo : 
                            (N445)? cache_pkt_i[45:38] : 
                            (N441)? sbuf_entry_lo[47:40] : 1'b0;
  assign data_mem_w_mask_li = (N26)? dma_data_mem_w_mask_lo : 
                              (N27)? sbuf_data_mem_w_mask : 1'b0;
  assign { N462, N461, N460, N459, N458, N457, N456 } = (N28)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N451)? { decode_v_r[10:10], decode_v_r[10:10], decode_v_r[10:10], decode_v_r[10:10], plru_decode_data_lo } : 1'b0;
  assign N28 = N450;
  assign { N469, N468, N467, N466, N465, N464, N463 } = (N28)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                        (N451)? { N452, N453, N454, N455, plru_decode_mask_lo } : 1'b0;
  assign stat_mem_v_li = (N29)? miss_stat_mem_v_lo : 
                         (N30)? N448 : 1'b0;
  assign N29 = N447;
  assign N30 = N446;
  assign stat_mem_w_li = (N29)? miss_stat_mem_w_lo : 
                         (N30)? N449 : 1'b0;
  assign stat_mem_addr_li = (N29)? miss_stat_mem_addr_lo : 
                            (N30)? addr_v_r[9:4] : 1'b0;
  assign stat_mem_data_li = (N29)? miss_stat_mem_data_lo : 
                            (N30)? { N462, N461, N460, N459, N458, N457, N456 } : 1'b0;
  assign stat_mem_w_mask_li = (N29)? miss_stat_mem_w_mask_lo : 
                              (N30)? { N469, N468, N467, N466, N465, N464, N463 } : 1'b0;
  assign { sbuf_entry_li_way_id__1_, sbuf_entry_li_way_id__0_ } = (N31)? chosen_way_lo : 
                                                                  (N32)? tag_hit_way_id : 1'b0;
  assign N31 = N471;
  assign N32 = N470;
  assign N33 = reset_i;
  assign N34 = ready_o | N33;
  assign N35 = ~N34;
  assign N119 = ~N33;
  assign N120 = ready_o & N119;
  assign N121 = reset_i;
  assign N122 = v_we_o | N121;
  assign N123 = ~N122;
  assign N291 = ~N121;
  assign N292 = v_we_o & N291;
  assign tag_hit_v[0] = N293 & valid_v_r[0];
  assign tag_hit_v[1] = N294 & valid_v_r[1];
  assign tag_hit_v[2] = N295 & valid_v_r[2];
  assign tag_hit_v[3] = N296 & valid_v_r[3];
  assign ld_st_miss = N472 & N473;
  assign N472 = ~tag_hit_found;
  assign N473 = decode_v_r[11] | decode_v_r[10];
  assign N297 = ~addr_v_r[10];
  assign N298 = ~addr_v_r[11];
  assign N299 = N297 & N298;
  assign N300 = N297 & addr_v_r[11];
  assign N301 = addr_v_r[10] & N298;
  assign N302 = addr_v_r[10] & addr_v_r[11];
  assign tagfl_hit = decode_v_r[8] & N303;
  assign aflinv_hit = N475 & tag_hit_found;
  assign N475 = N474 | decode_v_r[3];
  assign N474 = decode_v_r[5] | decode_v_r[4];
  assign N304 = ~tag_hit_found;
  assign N305 = tag_hit_found;
  assign N306 = ~tag_hit_way_id[0];
  assign N307 = ~tag_hit_way_id[1];
  assign N308 = N306 & N307;
  assign N309 = N306 & tag_hit_way_id[1];
  assign N310 = tag_hit_way_id[0] & N307;
  assign N311 = tag_hit_way_id[0] & tag_hit_way_id[1];
  assign N313 = ~N312;
  assign alock_miss = decode_v_r[2] & N314;
  assign N315 = ~tag_hit_found;
  assign N316 = tag_hit_found;
  assign N317 = ~tag_hit_way_id[0];
  assign N318 = ~tag_hit_way_id[1];
  assign N319 = N317 & N318;
  assign N320 = N317 & tag_hit_way_id[1];
  assign N321 = tag_hit_way_id[0] & N318;
  assign N322 = tag_hit_way_id[0] & tag_hit_way_id[1];
  assign aunlock_hit = decode_v_r[1] & N324;
  assign miss_v = N477 & N481;
  assign N477 = N476 & v_v_r;
  assign N476 = ~decode_v_r[9];
  assign N481 = N480 | aunlock_hit;
  assign N480 = N479 | alock_miss;
  assign N479 = N478 | aflinv_hit;
  assign N478 = ld_st_miss | tagfl_hit;
  assign retval_op_v = N482 | decode_v_r[6];
  assign N482 = decode_v_r[11] | decode_v_r[7];
  assign n_0_net_ = v_o & yumi_i;
  assign sbuf_data_mem_w_mask[3] = sbuf_way_decode[0] & sbuf_entry_lo[5];
  assign sbuf_data_mem_w_mask[2] = sbuf_way_decode[0] & sbuf_entry_lo[4];
  assign sbuf_data_mem_w_mask[1] = sbuf_way_decode[0] & sbuf_entry_lo[3];
  assign sbuf_data_mem_w_mask[0] = sbuf_way_decode[0] & sbuf_entry_lo[2];
  assign sbuf_data_mem_w_mask[7] = sbuf_way_decode[1] & sbuf_entry_lo[5];
  assign sbuf_data_mem_w_mask[6] = sbuf_way_decode[1] & sbuf_entry_lo[4];
  assign sbuf_data_mem_w_mask[5] = sbuf_way_decode[1] & sbuf_entry_lo[3];
  assign sbuf_data_mem_w_mask[4] = sbuf_way_decode[1] & sbuf_entry_lo[2];
  assign sbuf_data_mem_w_mask[11] = sbuf_way_decode[2] & sbuf_entry_lo[5];
  assign sbuf_data_mem_w_mask[10] = sbuf_way_decode[2] & sbuf_entry_lo[4];
  assign sbuf_data_mem_w_mask[9] = sbuf_way_decode[2] & sbuf_entry_lo[3];
  assign sbuf_data_mem_w_mask[8] = sbuf_way_decode[2] & sbuf_entry_lo[2];
  assign sbuf_data_mem_w_mask[15] = sbuf_way_decode[3] & sbuf_entry_lo[5];
  assign sbuf_data_mem_w_mask[14] = sbuf_way_decode[3] & sbuf_entry_lo[4];
  assign sbuf_data_mem_w_mask[13] = sbuf_way_decode[3] & sbuf_entry_lo[3];
  assign sbuf_data_mem_w_mask[12] = sbuf_way_decode[3] & sbuf_entry_lo[2];
  assign N325 = decode_v_r[12];
  assign N326 = ~N325;
  assign N327 = decode_v_r[12];
  assign N328 = ~N327;
  assign N329 = ~miss_v;
  assign N330 = miss_v;
  assign ld_data_masked[31] = snoop_or_ld_data[31] & expanded_mask_v[31];
  assign ld_data_masked[30] = snoop_or_ld_data[30] & expanded_mask_v[30];
  assign ld_data_masked[29] = snoop_or_ld_data[29] & expanded_mask_v[29];
  assign ld_data_masked[28] = snoop_or_ld_data[28] & expanded_mask_v[28];
  assign ld_data_masked[27] = snoop_or_ld_data[27] & expanded_mask_v[27];
  assign ld_data_masked[26] = snoop_or_ld_data[26] & expanded_mask_v[26];
  assign ld_data_masked[25] = snoop_or_ld_data[25] & expanded_mask_v[25];
  assign ld_data_masked[24] = snoop_or_ld_data[24] & expanded_mask_v[24];
  assign ld_data_masked[23] = snoop_or_ld_data[23] & expanded_mask_v[23];
  assign ld_data_masked[22] = snoop_or_ld_data[22] & expanded_mask_v[22];
  assign ld_data_masked[21] = snoop_or_ld_data[21] & expanded_mask_v[21];
  assign ld_data_masked[20] = snoop_or_ld_data[20] & expanded_mask_v[20];
  assign ld_data_masked[19] = snoop_or_ld_data[19] & expanded_mask_v[19];
  assign ld_data_masked[18] = snoop_or_ld_data[18] & expanded_mask_v[18];
  assign ld_data_masked[17] = snoop_or_ld_data[17] & expanded_mask_v[17];
  assign ld_data_masked[16] = snoop_or_ld_data[16] & expanded_mask_v[16];
  assign ld_data_masked[15] = snoop_or_ld_data[15] & expanded_mask_v[15];
  assign ld_data_masked[14] = snoop_or_ld_data[14] & expanded_mask_v[14];
  assign ld_data_masked[13] = snoop_or_ld_data[13] & expanded_mask_v[13];
  assign ld_data_masked[12] = snoop_or_ld_data[12] & expanded_mask_v[12];
  assign ld_data_masked[11] = snoop_or_ld_data[11] & expanded_mask_v[11];
  assign ld_data_masked[10] = snoop_or_ld_data[10] & expanded_mask_v[10];
  assign ld_data_masked[9] = snoop_or_ld_data[9] & expanded_mask_v[9];
  assign ld_data_masked[8] = snoop_or_ld_data[8] & expanded_mask_v[8];
  assign ld_data_masked[7] = snoop_or_ld_data[7] & expanded_mask_v[7];
  assign ld_data_masked[6] = snoop_or_ld_data[6] & expanded_mask_v[6];
  assign ld_data_masked[5] = snoop_or_ld_data[5] & expanded_mask_v[5];
  assign ld_data_masked[4] = snoop_or_ld_data[4] & expanded_mask_v[4];
  assign ld_data_masked[3] = snoop_or_ld_data[3] & expanded_mask_v[3];
  assign ld_data_masked[2] = snoop_or_ld_data[2] & expanded_mask_v[2];
  assign ld_data_masked[1] = snoop_or_ld_data[1] & expanded_mask_v[1];
  assign ld_data_masked[0] = snoop_or_ld_data[0] & expanded_mask_v[0];
  assign ld_data_final_li_0__31_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__30_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__29_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__28_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__27_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__26_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__25_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__24_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__23_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__22_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__21_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__20_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__19_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__18_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__17_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__16_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__15_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__14_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__13_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__12_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__11_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__10_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__9_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__8_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_1__31_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__30_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__29_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__28_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__27_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__26_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__25_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__24_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__23_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__22_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__21_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__20_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__19_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__18_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__17_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__16_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign N331 = ~retval_op_v;
  assign N332 = decode_v_r[7];
  assign N333 = decode_v_r[6];
  assign N334 = decode_v_r[12];
  assign N335 = N333 | N332;
  assign N336 = N334 | N335;
  assign N337 = ~N336;
  assign N338 = ~addr_v_r[10];
  assign N339 = ~addr_v_r[11];
  assign N340 = N338 & N339;
  assign N341 = N338 & addr_v_r[11];
  assign N342 = addr_v_r[10] & N339;
  assign N343 = addr_v_r[10] & addr_v_r[11];
  assign N345 = ~addr_v_r[10];
  assign N346 = ~addr_v_r[11];
  assign N347 = N345 & N346;
  assign N348 = N345 & addr_v_r[11];
  assign N349 = addr_v_r[10] & N346;
  assign N350 = addr_v_r[10] & addr_v_r[11];
  assign N352 = ~addr_v_r[10];
  assign N353 = ~addr_v_r[11];
  assign N354 = N352 & N353;
  assign N355 = N352 & addr_v_r[11];
  assign N356 = addr_v_r[10] & N353;
  assign N357 = addr_v_r[10] & addr_v_r[11];
  assign N408 = ~N332;
  assign N409 = N333 & N408;
  assign N410 = ~N333;
  assign N411 = N408 & N410;
  assign N412 = N334 & N411;
  assign N413 = ~miss_v;
  assign N414 = miss_v;
  assign v_o = v_v_r & N415;
  assign N416 = ~v_v_r;
  assign N417 = v_o & yumi_i;
  assign N418 = ~miss_v;
  assign N419 = miss_v;
  assign N420 = N490 & N491;
  assign N490 = N488 & N489;
  assign N488 = N486 & N487;
  assign N486 = N484 & N485;
  assign N484 = ~N483;
  assign N483 = decode[9] & v_i;
  assign N485 = ~miss_tag_mem_v_lo;
  assign N487 = ~dma_data_mem_v_lo;
  assign N489 = ~recover_lo;
  assign N491 = ~dma_evict_lo;
  assign N421 = ~v_tl_r;
  assign N422 = v_we_o & tl_ready;
  assign tagst_write_en = N492 & v_i;
  assign N492 = decode[9] & ready_o;
  assign tag_mem_v_li = N498 | N500;
  assign N498 = N497 | miss_tag_mem_v_lo;
  assign N497 = N494 | N496;
  assign N494 = N493 & v_i;
  assign N493 = decode[0] & ready_o;
  assign N496 = N495 & v_tl_r;
  assign N495 = recover_lo & decode_tl_r[0];
  assign N500 = N499 & v_i;
  assign N499 = decode[9] & ready_o;
  assign N423 = ~miss_v;
  assign N424 = miss_v;
  assign N425 = ~miss_v;
  assign N426 = miss_v;
  assign N427 = miss_tag_mem_v_lo | recover_lo;
  assign N428 = ~N427;
  assign N435 = ~recover_lo;
  assign N436 = miss_tag_mem_v_lo & N435;
  assign data_mem_v_li = N506 | N507;
  assign N506 = N505 | dma_data_mem_v_lo;
  assign N505 = N502 | N504;
  assign N502 = N501 & ready_o;
  assign N501 = v_i & decode[11];
  assign N504 = N503 & decode_tl_r[11];
  assign N503 = v_tl_r & recover_lo;
  assign N507 = sbuf_v_lo & sbuf_yumi_li;
  assign data_mem_w_li = dma_data_mem_w_lo | N508;
  assign N508 = sbuf_v_lo & sbuf_yumi_li;
  assign N437 = ~dma_data_mem_w_lo;
  assign N438 = N509 & ready_o;
  assign N509 = decode[11] & v_i;
  assign N439 = dma_data_mem_v_lo | recover_lo;
  assign N440 = N438 | N439;
  assign N441 = ~N440;
  assign N442 = dma_data_mem_v_lo & N435;
  assign N443 = ~dma_data_mem_v_lo;
  assign N444 = N435 & N443;
  assign N445 = N438 & N444;
  assign N446 = ~miss_v;
  assign N447 = miss_v;
  assign N448 = N512 & yumi_i;
  assign N512 = N511 & v_o;
  assign N511 = N510 | decode_v_r[9];
  assign N510 = decode_v_r[10] | decode_v_r[11];
  assign N449 = N515 & yumi_i;
  assign N515 = N514 & v_o;
  assign N514 = N513 | decode_v_r[9];
  assign N513 = decode_v_r[10] | decode_v_r[11];
  assign N450 = decode_v_r[9];
  assign N451 = ~N450;
  assign N452 = decode_v_r[10] & tag_hit_v[3];
  assign N453 = decode_v_r[10] & tag_hit_v[2];
  assign N454 = decode_v_r[10] & tag_hit_v[1];
  assign N455 = decode_v_r[10] & tag_hit_v[0];
  assign sbuf_v_li = N516 & yumi_i;
  assign N516 = decode_v_r[10] & v_o;
  assign N470 = ~miss_v;
  assign N471 = miss_v;
  assign sbuf_yumi_li = N520 & N487;
  assign N520 = sbuf_v_lo & N519;
  assign N519 = ~N518;
  assign N518 = N517 & ready_o;
  assign N517 = decode[11] & v_i;
  assign bypass_v_li = N521 & v_we_o;
  assign N521 = decode_tl_r[11] & v_tl_r;

  always @(posedge clk_i) begin
    if(N38) begin
      { data_tl_r[31:0] } <= { N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87 };
      { decode_tl_r[15:0] } <= { N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39 };
      { mask_tl_r[3:0] } <= { N58, N57, N56, N55 };
      { addr_tl_r[27:0] } <= { N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59 };
    end 
    if(N36) begin
      v_tl_r <= N37;
    end 
    if(N290) begin
      { ld_data_v_r[127:29] } <= { data_mem_data_lo[127:29] };
    end 
    if(N289) begin
      { ld_data_v_r[28:0] } <= { data_mem_data_lo[28:0] };
    end 
    if(N124) begin
      v_v_r <= N125;
    end 
    if(N133) begin
      { tag_v_r[71:6] } <= { N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134 };
      { mask_v_r[1:1] } <= { N202 };
      { lock_v_r[3:0] } <= { N288, N287, N286, N285 };
    end 
    if(N126) begin
      { tag_v_r[5:0] } <= { N132, N131, N130, N129, N128, N127 };
      { mask_v_r[3:2] } <= { N204, N203 };
      { decode_v_r[15:0] } <= { N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205 };
      { addr_v_r[27:0] } <= { N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221 };
      { data_v_r[31:0] } <= { N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249 };
      { valid_v_r[3:0] } <= { N284, N283, N282, N281 };
    end 
    if(N200) begin
      { mask_v_r[0:0] } <= { N201 };
    end 
  end


endmodule

