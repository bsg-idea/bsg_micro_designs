

module top
(
  clk,
  reset,
  calibration_done_i,
  valid_i,
  data_i,
  yumi_o,
  in_top_channel_i,
  out_top_channel_i,
  valid_o,
  data_o,
  yumi_i
);

  input [9:0] valid_i;
  input [319:0] data_i;
  output [9:0] yumi_o;
  input [3:0] in_top_channel_i;
  input [2:0] out_top_channel_i;
  output [159:0] data_o;
  input clk;
  input reset;
  input calibration_done_i;
  input yumi_i;
  output valid_o;

  bsg_assembler_in
  wrapper
  (
    .valid_i(valid_i),
    .data_i(data_i),
    .yumi_o(yumi_o),
    .in_top_channel_i(in_top_channel_i),
    .out_top_channel_i(out_top_channel_i),
    .data_o(data_o),
    .clk(clk),
    .reset(reset),
    .calibration_done_i(calibration_done_i),
    .yumi_i(yumi_i),
    .valid_o(valid_o)
  );


endmodule



module bsg_make_2D_array_width_p32_items_p5
(
  i,
  o
);

  input [159:0] i;
  output [159:0] o;
  wire [159:0] o;
  assign o[159] = i[159];
  assign o[158] = i[158];
  assign o[157] = i[157];
  assign o[156] = i[156];
  assign o[155] = i[155];
  assign o[154] = i[154];
  assign o[153] = i[153];
  assign o[152] = i[152];
  assign o[151] = i[151];
  assign o[150] = i[150];
  assign o[149] = i[149];
  assign o[148] = i[148];
  assign o[147] = i[147];
  assign o[146] = i[146];
  assign o[145] = i[145];
  assign o[144] = i[144];
  assign o[143] = i[143];
  assign o[142] = i[142];
  assign o[141] = i[141];
  assign o[140] = i[140];
  assign o[139] = i[139];
  assign o[138] = i[138];
  assign o[137] = i[137];
  assign o[136] = i[136];
  assign o[135] = i[135];
  assign o[134] = i[134];
  assign o[133] = i[133];
  assign o[132] = i[132];
  assign o[131] = i[131];
  assign o[130] = i[130];
  assign o[129] = i[129];
  assign o[128] = i[128];
  assign o[127] = i[127];
  assign o[126] = i[126];
  assign o[125] = i[125];
  assign o[124] = i[124];
  assign o[123] = i[123];
  assign o[122] = i[122];
  assign o[121] = i[121];
  assign o[120] = i[120];
  assign o[119] = i[119];
  assign o[118] = i[118];
  assign o[117] = i[117];
  assign o[116] = i[116];
  assign o[115] = i[115];
  assign o[114] = i[114];
  assign o[113] = i[113];
  assign o[112] = i[112];
  assign o[111] = i[111];
  assign o[110] = i[110];
  assign o[109] = i[109];
  assign o[108] = i[108];
  assign o[107] = i[107];
  assign o[106] = i[106];
  assign o[105] = i[105];
  assign o[104] = i[104];
  assign o[103] = i[103];
  assign o[102] = i[102];
  assign o[101] = i[101];
  assign o[100] = i[100];
  assign o[99] = i[99];
  assign o[98] = i[98];
  assign o[97] = i[97];
  assign o[96] = i[96];
  assign o[95] = i[95];
  assign o[94] = i[94];
  assign o[93] = i[93];
  assign o[92] = i[92];
  assign o[91] = i[91];
  assign o[90] = i[90];
  assign o[89] = i[89];
  assign o[88] = i[88];
  assign o[87] = i[87];
  assign o[86] = i[86];
  assign o[85] = i[85];
  assign o[84] = i[84];
  assign o[83] = i[83];
  assign o[82] = i[82];
  assign o[81] = i[81];
  assign o[80] = i[80];
  assign o[79] = i[79];
  assign o[78] = i[78];
  assign o[77] = i[77];
  assign o[76] = i[76];
  assign o[75] = i[75];
  assign o[74] = i[74];
  assign o[73] = i[73];
  assign o[72] = i[72];
  assign o[71] = i[71];
  assign o[70] = i[70];
  assign o[69] = i[69];
  assign o[68] = i[68];
  assign o[67] = i[67];
  assign o[66] = i[66];
  assign o[65] = i[65];
  assign o[64] = i[64];
  assign o[63] = i[63];
  assign o[62] = i[62];
  assign o[61] = i[61];
  assign o[60] = i[60];
  assign o[59] = i[59];
  assign o[58] = i[58];
  assign o[57] = i[57];
  assign o[56] = i[56];
  assign o[55] = i[55];
  assign o[54] = i[54];
  assign o[53] = i[53];
  assign o[52] = i[52];
  assign o[51] = i[51];
  assign o[50] = i[50];
  assign o[49] = i[49];
  assign o[48] = i[48];
  assign o[47] = i[47];
  assign o[46] = i[46];
  assign o[45] = i[45];
  assign o[44] = i[44];
  assign o[43] = i[43];
  assign o[42] = i[42];
  assign o[41] = i[41];
  assign o[40] = i[40];
  assign o[39] = i[39];
  assign o[38] = i[38];
  assign o[37] = i[37];
  assign o[36] = i[36];
  assign o[35] = i[35];
  assign o[34] = i[34];
  assign o[33] = i[33];
  assign o[32] = i[32];
  assign o[31] = i[31];
  assign o[30] = i[30];
  assign o[29] = i[29];
  assign o[28] = i[28];
  assign o[27] = i[27];
  assign o[26] = i[26];
  assign o[25] = i[25];
  assign o[24] = i[24];
  assign o[23] = i[23];
  assign o[22] = i[22];
  assign o[21] = i[21];
  assign o[20] = i[20];
  assign o[19] = i[19];
  assign o[18] = i[18];
  assign o[17] = i[17];
  assign o[16] = i[16];
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_rotate_right_width_p10
(
  data_i,
  rot_i,
  o
);

  input [9:0] data_i;
  input [3:0] rot_i;
  output [9:0] o;
  wire [9:0] o;
  wire sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,
  sv2v_dc_9,sv2v_dc_10;
  assign { sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, o } = { data_i, data_i } >> rot_i;

endmodule



module bsg_circular_ptr_slots_p10_max_add_p5
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [2:0] add_i;
  output [3:0] o;
  output [3:0] n_o;
  input clk;
  input reset_i;
  wire [3:0] o,n_o,ptr_nowrap;
  wire N0,N1,N2,N3,N4,N5,N6,N7;
  wire [4:0] ptr_wrap;
  reg o_3_sv2v_reg,o_2_sv2v_reg,o_1_sv2v_reg,o_0_sv2v_reg;
  assign o[3] = o_3_sv2v_reg;
  assign o[2] = o_2_sv2v_reg;
  assign o[1] = o_1_sv2v_reg;
  assign o[0] = o_0_sv2v_reg;
  assign ptr_nowrap = o + add_i;
  assign { N6, N5, N4, N3, N2 } = o - { 1'b1, 1'b0, 1'b1, 1'b0 };
  assign ptr_wrap = { N6, N5, N4, N3, N2 } + add_i;
  assign n_o = (N0)? ptr_wrap[3:0] : 
               (N1)? ptr_nowrap : 1'b0;
  assign N0 = N7;
  assign N1 = ptr_wrap[4];
  assign N7 = ~ptr_wrap[4];

  always @(posedge clk) begin
    if(reset_i) begin
      o_3_sv2v_reg <= 1'b0;
      o_2_sv2v_reg <= 1'b0;
      o_1_sv2v_reg <= 1'b0;
      o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      o_3_sv2v_reg <= n_o[3];
      o_2_sv2v_reg <= n_o[2];
      o_1_sv2v_reg <= n_o[1];
      o_0_sv2v_reg <= n_o[0];
    end 
  end


endmodule



module bsg_rr_f2f_input_width_p32_num_in_p10_middle_meet_p5
(
  clk,
  reset,
  valid_i,
  data_i,
  data_head_o,
  valid_head_o,
  go_channels_i,
  go_cnt_i,
  yumi_o
);

  input [9:0] valid_i;
  input [319:0] data_i;
  output [159:0] data_head_o;
  output [4:0] valid_head_o;
  input [4:0] go_channels_i;
  input [2:0] go_cnt_i;
  output [9:0] yumi_o;
  input clk;
  input reset;
  wire [159:0] data_head_o,data_head_o_flat_pretrunc;
  wire [4:0] valid_head_o;
  wire [9:0] yumi_o;
  wire sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,
  sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,sv2v_dc_13,sv2v_dc_14,sv2v_dc_15,
  sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,sv2v_dc_20,sv2v_dc_21,sv2v_dc_22,
  sv2v_dc_23,sv2v_dc_24,sv2v_dc_25,sv2v_dc_26,sv2v_dc_27,sv2v_dc_28,sv2v_dc_29,
  sv2v_dc_30,sv2v_dc_31,sv2v_dc_32,sv2v_dc_33,sv2v_dc_34,sv2v_dc_35,sv2v_dc_36,sv2v_dc_37,
  sv2v_dc_38,sv2v_dc_39,sv2v_dc_40,sv2v_dc_41,sv2v_dc_42,sv2v_dc_43,sv2v_dc_44,
  sv2v_dc_45,sv2v_dc_46,sv2v_dc_47,sv2v_dc_48,sv2v_dc_49,sv2v_dc_50,sv2v_dc_51,
  sv2v_dc_52,sv2v_dc_53,sv2v_dc_54,sv2v_dc_55,sv2v_dc_56,sv2v_dc_57,sv2v_dc_58,sv2v_dc_59,
  sv2v_dc_60,sv2v_dc_61,sv2v_dc_62,sv2v_dc_63,sv2v_dc_64,sv2v_dc_65,sv2v_dc_66,
  sv2v_dc_67,sv2v_dc_68,sv2v_dc_69,sv2v_dc_70,sv2v_dc_71,sv2v_dc_72,sv2v_dc_73,
  sv2v_dc_74,sv2v_dc_75,sv2v_dc_76,sv2v_dc_77,sv2v_dc_78,sv2v_dc_79,sv2v_dc_80,
  sv2v_dc_81,sv2v_dc_82,sv2v_dc_83,sv2v_dc_84,sv2v_dc_85,sv2v_dc_86,sv2v_dc_87,sv2v_dc_88,
  sv2v_dc_89,sv2v_dc_90,sv2v_dc_91,sv2v_dc_92,sv2v_dc_93,sv2v_dc_94,sv2v_dc_95,
  sv2v_dc_96,sv2v_dc_97,sv2v_dc_98,sv2v_dc_99,sv2v_dc_100,sv2v_dc_101,sv2v_dc_102,
  sv2v_dc_103,sv2v_dc_104,sv2v_dc_105,sv2v_dc_106,sv2v_dc_107,sv2v_dc_108,sv2v_dc_109,
  sv2v_dc_110,sv2v_dc_111,sv2v_dc_112,sv2v_dc_113,sv2v_dc_114,sv2v_dc_115,
  sv2v_dc_116,sv2v_dc_117,sv2v_dc_118,sv2v_dc_119,sv2v_dc_120,sv2v_dc_121,sv2v_dc_122,
  sv2v_dc_123,sv2v_dc_124,sv2v_dc_125,sv2v_dc_126,sv2v_dc_127,sv2v_dc_128,sv2v_dc_129,
  sv2v_dc_130,sv2v_dc_131,sv2v_dc_132,sv2v_dc_133,sv2v_dc_134,sv2v_dc_135,
  sv2v_dc_136,sv2v_dc_137,sv2v_dc_138,sv2v_dc_139,sv2v_dc_140,sv2v_dc_141,sv2v_dc_142,
  sv2v_dc_143,sv2v_dc_144,sv2v_dc_145,sv2v_dc_146,sv2v_dc_147,sv2v_dc_148,sv2v_dc_149,
  sv2v_dc_150,sv2v_dc_151,sv2v_dc_152,sv2v_dc_153,sv2v_dc_154,sv2v_dc_155,
  sv2v_dc_156,sv2v_dc_157,sv2v_dc_158,sv2v_dc_159,sv2v_dc_160,sv2v_dc_161,sv2v_dc_162,
  sv2v_dc_163,sv2v_dc_164,sv2v_dc_165,sv2v_dc_166,sv2v_dc_167,sv2v_dc_168,sv2v_dc_169,
  sv2v_dc_170,sv2v_dc_171,sv2v_dc_172,sv2v_dc_173,sv2v_dc_174,sv2v_dc_175,
  sv2v_dc_176,sv2v_dc_177,sv2v_dc_178,sv2v_dc_179,sv2v_dc_180,sv2v_dc_181,sv2v_dc_182,
  sv2v_dc_183,sv2v_dc_184,sv2v_dc_185,sv2v_dc_186,sv2v_dc_187,sv2v_dc_188,sv2v_dc_189,
  sv2v_dc_190,sv2v_dc_191,sv2v_dc_192,sv2v_dc_193,sv2v_dc_194,sv2v_dc_195,
  sv2v_dc_196,sv2v_dc_197,sv2v_dc_198,sv2v_dc_199,sv2v_dc_200,sv2v_dc_201,sv2v_dc_202,
  sv2v_dc_203,sv2v_dc_204,sv2v_dc_205,sv2v_dc_206,sv2v_dc_207,sv2v_dc_208,sv2v_dc_209,
  sv2v_dc_210,sv2v_dc_211,sv2v_dc_212,sv2v_dc_213,sv2v_dc_214,sv2v_dc_215,
  sv2v_dc_216,sv2v_dc_217,sv2v_dc_218,sv2v_dc_219,sv2v_dc_220,sv2v_dc_221,sv2v_dc_222,
  sv2v_dc_223,sv2v_dc_224,sv2v_dc_225,sv2v_dc_226,sv2v_dc_227,sv2v_dc_228,sv2v_dc_229,
  sv2v_dc_230,sv2v_dc_231,sv2v_dc_232,sv2v_dc_233,sv2v_dc_234,sv2v_dc_235,
  sv2v_dc_236,sv2v_dc_237,sv2v_dc_238,sv2v_dc_239,sv2v_dc_240,sv2v_dc_241,sv2v_dc_242,
  sv2v_dc_243,sv2v_dc_244,sv2v_dc_245,sv2v_dc_246,sv2v_dc_247,sv2v_dc_248,sv2v_dc_249,
  sv2v_dc_250,sv2v_dc_251,sv2v_dc_252,sv2v_dc_253,sv2v_dc_254,sv2v_dc_255,
  sv2v_dc_256,sv2v_dc_257,sv2v_dc_258,sv2v_dc_259,sv2v_dc_260,sv2v_dc_261,sv2v_dc_262,
  sv2v_dc_263,sv2v_dc_264,sv2v_dc_265,sv2v_dc_266,sv2v_dc_267,sv2v_dc_268,sv2v_dc_269,
  sv2v_dc_270,sv2v_dc_271,sv2v_dc_272,sv2v_dc_273,sv2v_dc_274,sv2v_dc_275,
  sv2v_dc_276,sv2v_dc_277,sv2v_dc_278,sv2v_dc_279,sv2v_dc_280,sv2v_dc_281,sv2v_dc_282,
  sv2v_dc_283,sv2v_dc_284,sv2v_dc_285,sv2v_dc_286,sv2v_dc_287,sv2v_dc_288,sv2v_dc_289,
  sv2v_dc_290,sv2v_dc_291,sv2v_dc_292,sv2v_dc_293,sv2v_dc_294,sv2v_dc_295,
  sv2v_dc_296,sv2v_dc_297,sv2v_dc_298,sv2v_dc_299,sv2v_dc_300,sv2v_dc_301,sv2v_dc_302,
  sv2v_dc_303,sv2v_dc_304,sv2v_dc_305,sv2v_dc_306,sv2v_dc_307,sv2v_dc_308,sv2v_dc_309,
  sv2v_dc_310,sv2v_dc_311,sv2v_dc_312,sv2v_dc_313,sv2v_dc_314,sv2v_dc_315,
  sv2v_dc_316,sv2v_dc_317,sv2v_dc_318,sv2v_dc_319,sv2v_dc_320,sv2v_dc_321,sv2v_dc_322,
  sv2v_dc_323,sv2v_dc_324,sv2v_dc_325,sv2v_dc_326,sv2v_dc_327,sv2v_dc_328,sv2v_dc_329,
  sv2v_dc_330,sv2v_dc_331,sv2v_dc_332,sv2v_dc_333,sv2v_dc_334,sv2v_dc_335,
  sv2v_dc_336,sv2v_dc_337,sv2v_dc_338,sv2v_dc_339,sv2v_dc_340,sv2v_dc_341,sv2v_dc_342,
  sv2v_dc_343,sv2v_dc_344,sv2v_dc_345,sv2v_dc_346,sv2v_dc_347,sv2v_dc_348,sv2v_dc_349,
  sv2v_dc_350,sv2v_dc_351,sv2v_dc_352,sv2v_dc_353,sv2v_dc_354,sv2v_dc_355,
  sv2v_dc_356,sv2v_dc_357,sv2v_dc_358,sv2v_dc_359,sv2v_dc_360,sv2v_dc_361,sv2v_dc_362,
  sv2v_dc_363,sv2v_dc_364,sv2v_dc_365,sv2v_dc_366,sv2v_dc_367,sv2v_dc_368,sv2v_dc_369,
  sv2v_dc_370,sv2v_dc_371,sv2v_dc_372,sv2v_dc_373,sv2v_dc_374,sv2v_dc_375,
  sv2v_dc_376,sv2v_dc_377,sv2v_dc_378,sv2v_dc_379,sv2v_dc_380,sv2v_dc_381,sv2v_dc_382,
  sv2v_dc_383,sv2v_dc_384,sv2v_dc_385,sv2v_dc_386,sv2v_dc_387,sv2v_dc_388,sv2v_dc_389,
  sv2v_dc_390,sv2v_dc_391,sv2v_dc_392,sv2v_dc_393,sv2v_dc_394,sv2v_dc_395,
  sv2v_dc_396,sv2v_dc_397,sv2v_dc_398,sv2v_dc_399,sv2v_dc_400,sv2v_dc_401,sv2v_dc_402,
  sv2v_dc_403,sv2v_dc_404,sv2v_dc_405,sv2v_dc_406,sv2v_dc_407,sv2v_dc_408,sv2v_dc_409,
  sv2v_dc_410,sv2v_dc_411,sv2v_dc_412,sv2v_dc_413,sv2v_dc_414,sv2v_dc_415,
  sv2v_dc_416,sv2v_dc_417,sv2v_dc_418,sv2v_dc_419,sv2v_dc_420,sv2v_dc_421,sv2v_dc_422,
  sv2v_dc_423,sv2v_dc_424,sv2v_dc_425,sv2v_dc_426,sv2v_dc_427,sv2v_dc_428,sv2v_dc_429,
  sv2v_dc_430,sv2v_dc_431,sv2v_dc_432,sv2v_dc_433,sv2v_dc_434,sv2v_dc_435,
  sv2v_dc_436,sv2v_dc_437,sv2v_dc_438,sv2v_dc_439,sv2v_dc_440,sv2v_dc_441,sv2v_dc_442,
  sv2v_dc_443,sv2v_dc_444,sv2v_dc_445,sv2v_dc_446,sv2v_dc_447,sv2v_dc_448,sv2v_dc_449,
  sv2v_dc_450,sv2v_dc_451,sv2v_dc_452,sv2v_dc_453,sv2v_dc_454,sv2v_dc_455,
  sv2v_dc_456,sv2v_dc_457,sv2v_dc_458,sv2v_dc_459,sv2v_dc_460,sv2v_dc_461,sv2v_dc_462,
  sv2v_dc_463,sv2v_dc_464,sv2v_dc_465,sv2v_dc_466,sv2v_dc_467,sv2v_dc_468,sv2v_dc_469,
  sv2v_dc_470,sv2v_dc_471,sv2v_dc_472,sv2v_dc_473,sv2v_dc_474,sv2v_dc_475,
  sv2v_dc_476,sv2v_dc_477,sv2v_dc_478,sv2v_dc_479,sv2v_dc_480,sv2v_dc_481,sv2v_dc_482,
  sv2v_dc_483,sv2v_dc_484,sv2v_dc_485,sv2v_dc_486,sv2v_dc_487,sv2v_dc_488,sv2v_dc_489,
  sv2v_dc_490,sv2v_dc_491,sv2v_dc_492,sv2v_dc_493,sv2v_dc_494,sv2v_dc_495,
  sv2v_dc_496,sv2v_dc_497,sv2v_dc_498;
  wire [3:0] iptr_r,iptr_r_data;
  wire [9:5] valid_head_o_pretrunc;

  bsg_make_2D_array_width_p32_items_p5
  bm2Da
  (
    .i(data_head_o_flat_pretrunc),
    .o(data_head_o)
  );


  bsg_rotate_right_width_p10
  valid_rr
  (
    .data_i(valid_i),
    .rot_i(iptr_r),
    .o({ valid_head_o_pretrunc, valid_head_o })
  );

  assign { sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25, sv2v_dc_26, sv2v_dc_27, sv2v_dc_28, sv2v_dc_29, sv2v_dc_30, sv2v_dc_31, sv2v_dc_32, sv2v_dc_33, sv2v_dc_34, sv2v_dc_35, sv2v_dc_36, sv2v_dc_37, sv2v_dc_38, sv2v_dc_39, sv2v_dc_40, sv2v_dc_41, sv2v_dc_42, sv2v_dc_43, sv2v_dc_44, sv2v_dc_45, sv2v_dc_46, sv2v_dc_47, sv2v_dc_48, sv2v_dc_49, sv2v_dc_50, sv2v_dc_51, sv2v_dc_52, sv2v_dc_53, sv2v_dc_54, sv2v_dc_55, sv2v_dc_56, sv2v_dc_57, sv2v_dc_58, sv2v_dc_59, sv2v_dc_60, sv2v_dc_61, sv2v_dc_62, sv2v_dc_63, sv2v_dc_64, sv2v_dc_65, sv2v_dc_66, sv2v_dc_67, sv2v_dc_68, sv2v_dc_69, sv2v_dc_70, sv2v_dc_71, sv2v_dc_72, sv2v_dc_73, sv2v_dc_74, sv2v_dc_75, sv2v_dc_76, sv2v_dc_77, sv2v_dc_78, sv2v_dc_79, sv2v_dc_80, sv2v_dc_81, sv2v_dc_82, sv2v_dc_83, sv2v_dc_84, sv2v_dc_85, sv2v_dc_86, sv2v_dc_87, sv2v_dc_88, sv2v_dc_89, sv2v_dc_90, sv2v_dc_91, sv2v_dc_92, sv2v_dc_93, sv2v_dc_94, sv2v_dc_95, sv2v_dc_96, sv2v_dc_97, sv2v_dc_98, sv2v_dc_99, sv2v_dc_100, sv2v_dc_101, sv2v_dc_102, sv2v_dc_103, sv2v_dc_104, sv2v_dc_105, sv2v_dc_106, sv2v_dc_107, sv2v_dc_108, sv2v_dc_109, sv2v_dc_110, sv2v_dc_111, sv2v_dc_112, sv2v_dc_113, sv2v_dc_114, sv2v_dc_115, sv2v_dc_116, sv2v_dc_117, sv2v_dc_118, sv2v_dc_119, sv2v_dc_120, sv2v_dc_121, sv2v_dc_122, sv2v_dc_123, sv2v_dc_124, sv2v_dc_125, sv2v_dc_126, sv2v_dc_127, sv2v_dc_128, sv2v_dc_129, sv2v_dc_130, sv2v_dc_131, sv2v_dc_132, sv2v_dc_133, sv2v_dc_134, sv2v_dc_135, sv2v_dc_136, sv2v_dc_137, sv2v_dc_138, sv2v_dc_139, sv2v_dc_140, sv2v_dc_141, sv2v_dc_142, sv2v_dc_143, sv2v_dc_144, sv2v_dc_145, sv2v_dc_146, sv2v_dc_147, sv2v_dc_148, sv2v_dc_149, sv2v_dc_150, sv2v_dc_151, sv2v_dc_152, sv2v_dc_153, sv2v_dc_154, sv2v_dc_155, sv2v_dc_156, sv2v_dc_157, sv2v_dc_158, sv2v_dc_159, sv2v_dc_160, sv2v_dc_161, sv2v_dc_162, sv2v_dc_163, sv2v_dc_164, sv2v_dc_165, sv2v_dc_166, sv2v_dc_167, sv2v_dc_168, sv2v_dc_169, sv2v_dc_170, sv2v_dc_171, sv2v_dc_172, sv2v_dc_173, sv2v_dc_174, sv2v_dc_175, sv2v_dc_176, sv2v_dc_177, sv2v_dc_178, sv2v_dc_179, sv2v_dc_180, sv2v_dc_181, sv2v_dc_182, sv2v_dc_183, sv2v_dc_184, sv2v_dc_185, sv2v_dc_186, sv2v_dc_187, sv2v_dc_188, sv2v_dc_189, sv2v_dc_190, sv2v_dc_191, sv2v_dc_192, sv2v_dc_193, sv2v_dc_194, sv2v_dc_195, sv2v_dc_196, sv2v_dc_197, sv2v_dc_198, sv2v_dc_199, sv2v_dc_200, sv2v_dc_201, sv2v_dc_202, sv2v_dc_203, sv2v_dc_204, sv2v_dc_205, sv2v_dc_206, sv2v_dc_207, sv2v_dc_208, sv2v_dc_209, sv2v_dc_210, sv2v_dc_211, sv2v_dc_212, sv2v_dc_213, sv2v_dc_214, sv2v_dc_215, sv2v_dc_216, sv2v_dc_217, sv2v_dc_218, sv2v_dc_219, sv2v_dc_220, sv2v_dc_221, sv2v_dc_222, sv2v_dc_223, sv2v_dc_224, sv2v_dc_225, sv2v_dc_226, sv2v_dc_227, sv2v_dc_228, sv2v_dc_229, sv2v_dc_230, sv2v_dc_231, sv2v_dc_232, sv2v_dc_233, sv2v_dc_234, sv2v_dc_235, sv2v_dc_236, sv2v_dc_237, sv2v_dc_238, sv2v_dc_239, sv2v_dc_240, sv2v_dc_241, sv2v_dc_242, sv2v_dc_243, sv2v_dc_244, sv2v_dc_245, sv2v_dc_246, sv2v_dc_247, sv2v_dc_248, sv2v_dc_249, sv2v_dc_250, sv2v_dc_251, sv2v_dc_252, sv2v_dc_253, sv2v_dc_254, sv2v_dc_255, sv2v_dc_256, sv2v_dc_257, sv2v_dc_258, sv2v_dc_259, sv2v_dc_260, sv2v_dc_261, sv2v_dc_262, sv2v_dc_263, sv2v_dc_264, sv2v_dc_265, sv2v_dc_266, sv2v_dc_267, sv2v_dc_268, sv2v_dc_269, sv2v_dc_270, sv2v_dc_271, sv2v_dc_272, sv2v_dc_273, sv2v_dc_274, sv2v_dc_275, sv2v_dc_276, sv2v_dc_277, sv2v_dc_278, sv2v_dc_279, sv2v_dc_280, sv2v_dc_281, sv2v_dc_282, sv2v_dc_283, sv2v_dc_284, sv2v_dc_285, sv2v_dc_286, sv2v_dc_287, sv2v_dc_288, sv2v_dc_289, sv2v_dc_290, sv2v_dc_291, sv2v_dc_292, sv2v_dc_293, sv2v_dc_294, sv2v_dc_295, sv2v_dc_296, sv2v_dc_297, sv2v_dc_298, sv2v_dc_299, sv2v_dc_300, sv2v_dc_301, sv2v_dc_302, sv2v_dc_303, sv2v_dc_304, sv2v_dc_305, sv2v_dc_306, sv2v_dc_307, sv2v_dc_308, sv2v_dc_309, sv2v_dc_310, sv2v_dc_311, sv2v_dc_312, sv2v_dc_313, sv2v_dc_314, sv2v_dc_315, sv2v_dc_316, sv2v_dc_317, sv2v_dc_318, sv2v_dc_319, sv2v_dc_320, sv2v_dc_321, sv2v_dc_322, sv2v_dc_323, sv2v_dc_324, sv2v_dc_325, sv2v_dc_326, sv2v_dc_327, sv2v_dc_328, sv2v_dc_329, sv2v_dc_330, sv2v_dc_331, sv2v_dc_332, sv2v_dc_333, sv2v_dc_334, sv2v_dc_335, sv2v_dc_336, sv2v_dc_337, sv2v_dc_338, sv2v_dc_339, sv2v_dc_340, sv2v_dc_341, sv2v_dc_342, sv2v_dc_343, sv2v_dc_344, sv2v_dc_345, sv2v_dc_346, sv2v_dc_347, sv2v_dc_348, sv2v_dc_349, sv2v_dc_350, sv2v_dc_351, sv2v_dc_352, sv2v_dc_353, sv2v_dc_354, sv2v_dc_355, sv2v_dc_356, sv2v_dc_357, sv2v_dc_358, sv2v_dc_359, sv2v_dc_360, sv2v_dc_361, sv2v_dc_362, sv2v_dc_363, sv2v_dc_364, sv2v_dc_365, sv2v_dc_366, sv2v_dc_367, sv2v_dc_368, sv2v_dc_369, sv2v_dc_370, sv2v_dc_371, sv2v_dc_372, sv2v_dc_373, sv2v_dc_374, sv2v_dc_375, sv2v_dc_376, sv2v_dc_377, sv2v_dc_378, sv2v_dc_379, sv2v_dc_380, sv2v_dc_381, sv2v_dc_382, sv2v_dc_383, sv2v_dc_384, sv2v_dc_385, sv2v_dc_386, sv2v_dc_387, sv2v_dc_388, sv2v_dc_389, sv2v_dc_390, sv2v_dc_391, sv2v_dc_392, sv2v_dc_393, sv2v_dc_394, sv2v_dc_395, sv2v_dc_396, sv2v_dc_397, sv2v_dc_398, sv2v_dc_399, sv2v_dc_400, sv2v_dc_401, sv2v_dc_402, sv2v_dc_403, sv2v_dc_404, sv2v_dc_405, sv2v_dc_406, sv2v_dc_407, sv2v_dc_408, sv2v_dc_409, sv2v_dc_410, sv2v_dc_411, sv2v_dc_412, sv2v_dc_413, sv2v_dc_414, sv2v_dc_415, sv2v_dc_416, sv2v_dc_417, sv2v_dc_418, sv2v_dc_419, sv2v_dc_420, sv2v_dc_421, sv2v_dc_422, sv2v_dc_423, sv2v_dc_424, sv2v_dc_425, sv2v_dc_426, sv2v_dc_427, sv2v_dc_428, sv2v_dc_429, sv2v_dc_430, sv2v_dc_431, sv2v_dc_432, sv2v_dc_433, sv2v_dc_434, sv2v_dc_435, sv2v_dc_436, sv2v_dc_437, sv2v_dc_438, sv2v_dc_439, sv2v_dc_440, sv2v_dc_441, sv2v_dc_442, sv2v_dc_443, sv2v_dc_444, sv2v_dc_445, sv2v_dc_446, sv2v_dc_447, sv2v_dc_448, sv2v_dc_449, sv2v_dc_450, sv2v_dc_451, sv2v_dc_452, sv2v_dc_453, sv2v_dc_454, sv2v_dc_455, sv2v_dc_456, sv2v_dc_457, sv2v_dc_458, sv2v_dc_459, sv2v_dc_460, sv2v_dc_461, sv2v_dc_462, sv2v_dc_463, sv2v_dc_464, sv2v_dc_465, sv2v_dc_466, sv2v_dc_467, sv2v_dc_468, sv2v_dc_469, sv2v_dc_470, sv2v_dc_471, sv2v_dc_472, sv2v_dc_473, sv2v_dc_474, sv2v_dc_475, sv2v_dc_476, sv2v_dc_477, sv2v_dc_478, sv2v_dc_479, sv2v_dc_480, data_head_o_flat_pretrunc } = { data_i, data_i } >> { iptr_r_data, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign { yumi_o, sv2v_dc_481, sv2v_dc_482, sv2v_dc_483, sv2v_dc_484, sv2v_dc_485, sv2v_dc_486, sv2v_dc_487, sv2v_dc_488, sv2v_dc_489, sv2v_dc_490 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, go_channels_i, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, go_channels_i } << iptr_r;

  bsg_circular_ptr_slots_p10_max_add_p5
  c_ptr
  (
    .clk(clk),
    .reset_i(reset),
    .add_i(go_cnt_i),
    .o(iptr_r),
    .n_o({ sv2v_dc_491, sv2v_dc_492, sv2v_dc_493, sv2v_dc_494 })
  );


  bsg_circular_ptr_slots_p10_max_add_p5
  c_ptr_data
  (
    .clk(clk),
    .reset_i(reset),
    .add_i(go_cnt_i),
    .o(iptr_r_data),
    .n_o({ sv2v_dc_495, sv2v_dc_496, sv2v_dc_497, sv2v_dc_498 })
  );


endmodule



module bsg_scan_width_p5_and_p1_lo_to_hi_p1
(
  i,
  o
);

  input [4:0] i;
  output [4:0] o;
  wire [4:0] o;
  wire t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__4_ = i[0] & 1'b1;
  assign t_1__3_ = i[1] & i[0];
  assign t_1__2_ = i[2] & i[1];
  assign t_1__1_ = i[3] & i[2];
  assign t_1__0_ = i[4] & i[3];
  assign t_2__4_ = t_1__4_ & 1'b1;
  assign t_2__3_ = t_1__3_ & 1'b1;
  assign t_2__2_ = t_1__2_ & t_1__4_;
  assign t_2__1_ = t_1__1_ & t_1__3_;
  assign t_2__0_ = t_1__0_ & t_1__2_;
  assign o[0] = t_2__4_ & 1'b1;
  assign o[1] = t_2__3_ & 1'b1;
  assign o[2] = t_2__2_ & 1'b1;
  assign o[3] = t_2__1_ & 1'b1;
  assign o[4] = t_2__0_ & t_2__4_;

endmodule



module bsg_encode_one_hot_width_p1
(
  i,
  addr_o,
  v_o
);

  input [0:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  assign v_o = i[0];
  assign addr_o[0] = 1'b0;

endmodule



module bsg_encode_one_hot_width_p2
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o,\aligned.vs ;
  wire v_o;
  wire [1:0] \aligned.addrs ;

  bsg_encode_one_hot_width_p1
  \aligned.left 
  (
    .i(i[0]),
    .addr_o(\aligned.addrs [0]),
    .v_o(\aligned.vs [0])
  );


  bsg_encode_one_hot_width_p1
  \aligned.right 
  (
    .i(i[1]),
    .addr_o(\aligned.addrs [1]),
    .v_o(addr_o[0])
  );

  assign v_o = addr_o[0] | \aligned.vs [0];

endmodule



module bsg_encode_one_hot_width_p4
(
  i,
  addr_o,
  v_o
);

  input [3:0] i;
  output [1:0] addr_o;
  output v_o;
  wire [1:0] addr_o,\aligned.addrs ;
  wire v_o;
  wire [0:0] \aligned.vs ;

  bsg_encode_one_hot_width_p2
  \aligned.left 
  (
    .i(i[1:0]),
    .addr_o(\aligned.addrs [0]),
    .v_o(\aligned.vs [0])
  );


  bsg_encode_one_hot_width_p2
  \aligned.right 
  (
    .i(i[3:2]),
    .addr_o(\aligned.addrs [1]),
    .v_o(addr_o[1])
  );

  assign v_o = addr_o[1] | \aligned.vs [0];
  assign addr_o[0] = \aligned.addrs [0] | \aligned.addrs [1];

endmodule



module bsg_encode_one_hot_width_p8
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [3:0] \aligned.addrs ;
  wire [0:0] \aligned.vs ;

  bsg_encode_one_hot_width_p4
  \aligned.left 
  (
    .i(i[3:0]),
    .addr_o(\aligned.addrs [1:0]),
    .v_o(\aligned.vs [0])
  );


  bsg_encode_one_hot_width_p4
  \aligned.right 
  (
    .i(i[7:4]),
    .addr_o(\aligned.addrs [3:2]),
    .v_o(addr_o[2])
  );

  assign v_o = addr_o[2] | \aligned.vs [0];
  assign addr_o[1] = \aligned.addrs [1] | \aligned.addrs [3];
  assign addr_o[0] = \aligned.addrs [0] | \aligned.addrs [2];

endmodule



module bsg_encode_one_hot_width_p6
(
  i,
  addr_o,
  v_o
);

  input [5:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;

  bsg_encode_one_hot_width_p8
  \unaligned.align 
  (
    .i({ 1'b0, 1'b0, i }),
    .addr_o(addr_o),
    .v_o(v_o)
  );


endmodule



module bsg_thermometer_count_width_p5
(
  i,
  o
);

  input [4:0] i;
  output [2:0] o;
  wire [2:0] o;
  wire N0,N1,N2,N3;
  wire [4:0] \big.one_hot ;

  bsg_encode_one_hot_width_p6
  \big.encode_one_hot 
  (
    .i({ i[4:4], \big.one_hot  }),
    .addr_o(o)
  );

  assign \big.one_hot [4] = N0 & i[3];
  assign N0 = ~i[4];
  assign \big.one_hot [3] = N1 & i[2];
  assign N1 = ~i[3];
  assign \big.one_hot [2] = N2 & i[1];
  assign N2 = ~i[2];
  assign \big.one_hot [1] = N3 & i[0];
  assign N3 = ~i[1];
  assign \big.one_hot [0] = ~i[0];

endmodule



module bsg_rr_f2f_middle_width_p32_middle_meet_p5
(
  valid_head_i,
  ready_head_i,
  go_channels_o,
  go_cnt_o
);

  input [4:0] valid_head_i;
  input [4:0] ready_head_i;
  output [4:0] go_channels_o;
  output [2:0] go_cnt_o;
  wire [4:0] go_channels_o,happy_channels;
  wire [2:0] go_cnt_o;

  bsg_scan_width_p5_and_p1_lo_to_hi_p1
  and_scan
  (
    .i(happy_channels),
    .o(go_channels_o)
  );


  bsg_thermometer_count_width_p5
  \genblk1.genblk1.thermo 
  (
    .i(go_channels_o),
    .o(go_cnt_o)
  );

  assign happy_channels[4] = valid_head_i[4] & ready_head_i[4];
  assign happy_channels[3] = valid_head_i[3] & ready_head_i[3];
  assign happy_channels[2] = valid_head_i[2] & ready_head_i[2];
  assign happy_channels[1] = valid_head_i[1] & ready_head_i[1];
  assign happy_channels[0] = valid_head_i[0] & ready_head_i[0];

endmodule



module bsg_rotate_right_width_p5
(
  data_i,
  rot_i,
  o
);

  input [4:0] data_i;
  input [2:0] rot_i;
  output [4:0] o;
  wire [4:0] o;
  wire sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5;
  assign { sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, o } = { data_i, data_i } >> rot_i;

endmodule



module bsg_circular_ptr_slots_p5_max_add_p5
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [2:0] add_i;
  output [2:0] o;
  output [2:0] n_o;
  input clk;
  input reset_i;
  wire [2:0] o,n_o,ptr_nowrap;
  wire N0,N1,N2,N3,N4,N5,N6;
  wire [3:0] ptr_wrap;
  reg o_2_sv2v_reg,o_1_sv2v_reg,o_0_sv2v_reg;
  assign o[2] = o_2_sv2v_reg;
  assign o[1] = o_1_sv2v_reg;
  assign o[0] = o_0_sv2v_reg;
  assign ptr_nowrap = o + add_i;
  assign { N5, N4, N3, N2 } = o - { 1'b1, 1'b0, 1'b1 };
  assign ptr_wrap = { N5, N4, N3, N2 } + add_i;
  assign n_o = (N0)? ptr_wrap[2:0] : 
               (N1)? ptr_nowrap : 1'b0;
  assign N0 = N6;
  assign N1 = ptr_wrap[3];
  assign N6 = ~ptr_wrap[3];

  always @(posedge clk) begin
    if(reset_i) begin
      o_2_sv2v_reg <= 1'b0;
      o_1_sv2v_reg <= 1'b0;
      o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      o_2_sv2v_reg <= n_o[2];
      o_1_sv2v_reg <= n_o[1];
      o_0_sv2v_reg <= n_o[0];
    end 
  end


endmodule



module bsg_rr_f2f_output_width_p32_num_out_p5_middle_meet_p5
(
  clk,
  reset,
  ready_i,
  ready_head_o,
  go_channels_i,
  go_cnt_i,
  data_head_i,
  valid_o,
  data_o
);

  input [4:0] ready_i;
  output [4:0] ready_head_o;
  input [4:0] go_channels_i;
  input [2:0] go_cnt_i;
  input [159:0] data_head_i;
  output [4:0] valid_o;
  output [159:0] data_o;
  input clk;
  input reset;
  wire [4:0] ready_head_o,valid_o;
  wire [159:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,
  sv2v_dc_7,sv2v_dc_8,sv2v_dc_9,sv2v_dc_10,sv2v_dc_11;
  wire [2:0] optr_r,optr_r_data;

  bsg_rotate_right_width_p5
  ready_rr
  (
    .data_i(ready_i),
    .rot_i(optr_r),
    .o(ready_head_o)
  );

  assign { valid_o, sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5 } = { go_channels_i, go_channels_i } << optr_r;

  bsg_circular_ptr_slots_p5_max_add_p5
  c_ptr
  (
    .clk(clk),
    .reset_i(reset),
    .add_i(go_cnt_i),
    .o(optr_r),
    .n_o({ sv2v_dc_6, sv2v_dc_7, sv2v_dc_8 })
  );


  bsg_circular_ptr_slots_p5_max_add_p5
  c_ptr_data
  (
    .clk(clk),
    .reset_i(reset),
    .add_i(go_cnt_i),
    .o(optr_r_data),
    .n_o({ sv2v_dc_9, sv2v_dc_10, sv2v_dc_11 })
  );

  assign N133 = optr_r_data[0] & N0;
  assign N0 = ~optr_r_data[1];
  assign N101 = N133 & optr_r_data[2];
  assign N134 = N1 & N2;
  assign N1 = ~optr_r_data[0];
  assign N2 = ~optr_r_data[1];
  assign N100 = N134 & optr_r_data[2];
  assign N135 = optr_r_data[0] & optr_r_data[1];
  assign N99 = N135 & N3;
  assign N3 = ~optr_r_data[2];
  assign N136 = N4 & optr_r_data[1];
  assign N4 = ~optr_r_data[0];
  assign N98 = N136 & N5;
  assign N5 = ~optr_r_data[2];
  assign N137 = optr_r_data[0] & N6;
  assign N6 = ~optr_r_data[1];
  assign N97 = N137 & N7;
  assign N7 = ~optr_r_data[2];
  assign N138 = N8 & N9;
  assign N8 = ~optr_r_data[0];
  assign N9 = ~optr_r_data[1];
  assign N96 = N138 & N10;
  assign N10 = ~optr_r_data[2];
  assign N139 = N11 & optr_r_data[1];
  assign N11 = ~optr_r_data[0];
  assign N108 = N139 & optr_r_data[2];
  assign N140 = optr_r_data[0] & N12;
  assign N12 = ~optr_r_data[1];
  assign N107 = N140 & optr_r_data[2];
  assign N141 = N13 & N14;
  assign N13 = ~optr_r_data[0];
  assign N14 = ~optr_r_data[1];
  assign N106 = N141 & optr_r_data[2];
  assign N142 = optr_r_data[0] & optr_r_data[1];
  assign N105 = N142 & N15;
  assign N15 = ~optr_r_data[2];
  assign N143 = N16 & optr_r_data[1];
  assign N16 = ~optr_r_data[0];
  assign N104 = N143 & N17;
  assign N17 = ~optr_r_data[2];
  assign N144 = optr_r_data[0] & N18;
  assign N18 = ~optr_r_data[1];
  assign N103 = N144 & N19;
  assign N19 = ~optr_r_data[2];
  assign N145 = N20 & N21;
  assign N20 = ~optr_r_data[0];
  assign N21 = ~optr_r_data[1];
  assign N102 = N145 & N22;
  assign N22 = ~optr_r_data[2];
  assign N146 = optr_r_data[0] & optr_r_data[1];
  assign N116 = N146 & optr_r_data[2];
  assign N147 = N23 & optr_r_data[1];
  assign N23 = ~optr_r_data[0];
  assign N115 = N147 & optr_r_data[2];
  assign N148 = optr_r_data[0] & N24;
  assign N24 = ~optr_r_data[1];
  assign N114 = N148 & optr_r_data[2];
  assign N149 = N25 & N26;
  assign N25 = ~optr_r_data[0];
  assign N26 = ~optr_r_data[1];
  assign N113 = N149 & optr_r_data[2];
  assign N150 = optr_r_data[0] & optr_r_data[1];
  assign N112 = N150 & N27;
  assign N27 = ~optr_r_data[2];
  assign N151 = N28 & optr_r_data[1];
  assign N28 = ~optr_r_data[0];
  assign N111 = N151 & N29;
  assign N29 = ~optr_r_data[2];
  assign N152 = optr_r_data[0] & N30;
  assign N30 = ~optr_r_data[1];
  assign N110 = N152 & N31;
  assign N31 = ~optr_r_data[2];
  assign N153 = N32 & N33;
  assign N32 = ~optr_r_data[0];
  assign N33 = ~optr_r_data[1];
  assign N109 = N153 & N34;
  assign N34 = ~optr_r_data[2];
  assign N154 = optr_r_data[0] & optr_r_data[1];
  assign N124 = N154 & optr_r_data[2];
  assign N155 = N35 & optr_r_data[1];
  assign N35 = ~optr_r_data[0];
  assign N123 = N155 & optr_r_data[2];
  assign N156 = optr_r_data[0] & N36;
  assign N36 = ~optr_r_data[1];
  assign N122 = N156 & optr_r_data[2];
  assign N157 = N37 & N38;
  assign N37 = ~optr_r_data[0];
  assign N38 = ~optr_r_data[1];
  assign N121 = N157 & optr_r_data[2];
  assign N158 = optr_r_data[0] & optr_r_data[1];
  assign N120 = N158 & N39;
  assign N39 = ~optr_r_data[2];
  assign N159 = N40 & optr_r_data[1];
  assign N40 = ~optr_r_data[0];
  assign N119 = N159 & N41;
  assign N41 = ~optr_r_data[2];
  assign N160 = optr_r_data[0] & N42;
  assign N42 = ~optr_r_data[1];
  assign N118 = N160 & N43;
  assign N43 = ~optr_r_data[2];
  assign N161 = N44 & N45;
  assign N44 = ~optr_r_data[0];
  assign N45 = ~optr_r_data[1];
  assign N117 = N161 & N46;
  assign N46 = ~optr_r_data[2];
  assign N162 = optr_r_data[0] & optr_r_data[1];
  assign N132 = N162 & optr_r_data[2];
  assign N163 = N47 & optr_r_data[1];
  assign N47 = ~optr_r_data[0];
  assign N131 = N163 & optr_r_data[2];
  assign N164 = optr_r_data[0] & N48;
  assign N48 = ~optr_r_data[1];
  assign N130 = N164 & optr_r_data[2];
  assign N165 = N49 & N50;
  assign N49 = ~optr_r_data[0];
  assign N50 = ~optr_r_data[1];
  assign N129 = N165 & optr_r_data[2];
  assign N166 = optr_r_data[0] & optr_r_data[1];
  assign N128 = N166 & N51;
  assign N51 = ~optr_r_data[2];
  assign N167 = N52 & optr_r_data[1];
  assign N52 = ~optr_r_data[0];
  assign N127 = N167 & N53;
  assign N53 = ~optr_r_data[2];
  assign N168 = optr_r_data[0] & N54;
  assign N54 = ~optr_r_data[1];
  assign N126 = N168 & N55;
  assign N55 = ~optr_r_data[2];
  assign N169 = N56 & N57;
  assign N56 = ~optr_r_data[0];
  assign N57 = ~optr_r_data[1];
  assign N125 = N169 & N58;
  assign N58 = ~optr_r_data[2];
  assign data_o[31:0] = (N59)? data_head_i[31:0] : 
                        (N60)? data_head_i[63:32] : 
                        (N61)? data_head_i[95:64] : 
                        (N62)? data_head_i[127:96] : 
                        (N63)? data_head_i[159:128] : 
                        (N64)? data_head_i[31:0] : 1'b0;
  assign N59 = N101;
  assign N60 = N100;
  assign N61 = N99;
  assign N62 = N98;
  assign N63 = N97;
  assign N64 = N96;
  assign data_o[63:32] = (N65)? data_head_i[31:0] : 
                         (N66)? data_head_i[63:32] : 
                         (N67)? data_head_i[95:64] : 
                         (N68)? data_head_i[127:96] : 
                         (N69)? data_head_i[159:128] : 
                         (N70)? data_head_i[31:0] : 
                         (N71)? data_head_i[63:32] : 1'b0;
  assign N65 = N108;
  assign N66 = N107;
  assign N67 = N106;
  assign N68 = N105;
  assign N69 = N104;
  assign N70 = N103;
  assign N71 = N102;
  assign data_o[95:64] = (N72)? data_head_i[31:0] : 
                         (N73)? data_head_i[63:32] : 
                         (N74)? data_head_i[95:64] : 
                         (N75)? data_head_i[127:96] : 
                         (N76)? data_head_i[159:128] : 
                         (N77)? data_head_i[31:0] : 
                         (N78)? data_head_i[63:32] : 
                         (N79)? data_head_i[95:64] : 1'b0;
  assign N72 = N116;
  assign N73 = N115;
  assign N74 = N114;
  assign N75 = N113;
  assign N76 = N112;
  assign N77 = N111;
  assign N78 = N110;
  assign N79 = N109;
  assign data_o[127:96] = (N80)? data_head_i[63:32] : 
                          (N81)? data_head_i[95:64] : 
                          (N82)? data_head_i[127:96] : 
                          (N83)? data_head_i[159:128] : 
                          (N84)? data_head_i[31:0] : 
                          (N85)? data_head_i[63:32] : 
                          (N86)? data_head_i[95:64] : 
                          (N87)? data_head_i[127:96] : 1'b0;
  assign N80 = N124;
  assign N81 = N123;
  assign N82 = N122;
  assign N83 = N121;
  assign N84 = N120;
  assign N85 = N119;
  assign N86 = N118;
  assign N87 = N117;
  assign data_o[159:128] = (N88)? data_head_i[95:64] : 
                           (N89)? data_head_i[127:96] : 
                           (N90)? data_head_i[159:128] : 
                           (N91)? data_head_i[31:0] : 
                           (N92)? data_head_i[63:32] : 
                           (N93)? data_head_i[95:64] : 
                           (N94)? data_head_i[127:96] : 
                           (N95)? data_head_i[159:128] : 1'b0;
  assign N88 = N132;
  assign N89 = N131;
  assign N90 = N130;
  assign N91 = N129;
  assign N92 = N128;
  assign N93 = N127;
  assign N94 = N126;
  assign N95 = N125;

endmodule



module bsg_round_robin_fifo_to_fifo_width_p32_num_in_p10_num_out_p5_in_channel_count_mask_p512
(
  clk,
  reset,
  valid_i,
  data_i,
  yumi_o,
  in_top_channel_i,
  out_top_channel_i,
  valid_o,
  data_o,
  ready_i
);

  input [9:0] valid_i;
  input [319:0] data_i;
  output [9:0] yumi_o;
  input [3:0] in_top_channel_i;
  input [2:0] out_top_channel_i;
  output [4:0] valid_o;
  output [159:0] data_o;
  input [4:0] ready_i;
  input clk;
  input reset;
  wire [9:0] yumi_o;
  wire [4:0] valid_o,go_channels;
  wire [159:0] data_o,data_o_flat,\oc_4_.out_chan.data_head_array ;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,yumi_int_o_9__9_,yumi_int_o_9__8_,
  yumi_int_o_9__7_,yumi_int_o_9__6_,yumi_int_o_9__5_,yumi_int_o_9__4_,
  yumi_int_o_9__3_,yumi_int_o_9__2_,yumi_int_o_9__1_,yumi_int_o_9__0_,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,valid_int_o_4__4_,valid_int_o_4__3_,valid_int_o_4__2_,
  valid_int_o_4__1_,valid_int_o_4__0_,N104,N105,N106,N107,data_int_o_4__159_,
  data_int_o_4__158_,data_int_o_4__157_,data_int_o_4__156_,data_int_o_4__155_,
  data_int_o_4__154_,data_int_o_4__153_,data_int_o_4__152_,data_int_o_4__151_,data_int_o_4__150_,
  data_int_o_4__149_,data_int_o_4__148_,data_int_o_4__147_,data_int_o_4__146_,
  data_int_o_4__145_,data_int_o_4__144_,data_int_o_4__143_,data_int_o_4__142_,
  data_int_o_4__141_,data_int_o_4__140_,data_int_o_4__139_,data_int_o_4__138_,
  data_int_o_4__137_,data_int_o_4__136_,data_int_o_4__135_,data_int_o_4__134_,
  data_int_o_4__133_,data_int_o_4__132_,data_int_o_4__131_,data_int_o_4__130_,data_int_o_4__129_,
  data_int_o_4__128_,data_int_o_4__127_,data_int_o_4__126_,data_int_o_4__125_,
  data_int_o_4__124_,data_int_o_4__123_,data_int_o_4__122_,data_int_o_4__121_,
  data_int_o_4__120_,data_int_o_4__119_,data_int_o_4__118_,data_int_o_4__117_,
  data_int_o_4__116_,data_int_o_4__115_,data_int_o_4__114_,data_int_o_4__113_,
  data_int_o_4__112_,data_int_o_4__111_,data_int_o_4__110_,data_int_o_4__109_,data_int_o_4__108_,
  data_int_o_4__107_,data_int_o_4__106_,data_int_o_4__105_,data_int_o_4__104_,
  data_int_o_4__103_,data_int_o_4__102_,data_int_o_4__101_,data_int_o_4__100_,
  data_int_o_4__99_,data_int_o_4__98_,data_int_o_4__97_,data_int_o_4__96_,data_int_o_4__95_,
  data_int_o_4__94_,data_int_o_4__93_,data_int_o_4__92_,data_int_o_4__91_,
  data_int_o_4__90_,data_int_o_4__89_,data_int_o_4__88_,data_int_o_4__87_,
  data_int_o_4__86_,data_int_o_4__85_,data_int_o_4__84_,data_int_o_4__83_,data_int_o_4__82_,
  data_int_o_4__81_,data_int_o_4__80_,data_int_o_4__79_,data_int_o_4__78_,
  data_int_o_4__77_,data_int_o_4__76_,data_int_o_4__75_,data_int_o_4__74_,data_int_o_4__73_,
  data_int_o_4__72_,data_int_o_4__71_,data_int_o_4__70_,data_int_o_4__69_,
  data_int_o_4__68_,data_int_o_4__67_,data_int_o_4__66_,data_int_o_4__65_,data_int_o_4__64_,
  data_int_o_4__63_,data_int_o_4__62_,data_int_o_4__61_,data_int_o_4__60_,
  data_int_o_4__59_,data_int_o_4__58_,data_int_o_4__57_,data_int_o_4__56_,data_int_o_4__55_,
  data_int_o_4__54_,data_int_o_4__53_,data_int_o_4__52_,data_int_o_4__51_,
  data_int_o_4__50_,data_int_o_4__49_,data_int_o_4__48_,data_int_o_4__47_,
  data_int_o_4__46_,data_int_o_4__45_,data_int_o_4__44_,data_int_o_4__43_,data_int_o_4__42_,
  data_int_o_4__41_,data_int_o_4__40_,data_int_o_4__39_,data_int_o_4__38_,
  data_int_o_4__37_,data_int_o_4__36_,data_int_o_4__35_,data_int_o_4__34_,data_int_o_4__33_,
  data_int_o_4__32_,data_int_o_4__31_,data_int_o_4__30_,data_int_o_4__29_,
  data_int_o_4__28_,data_int_o_4__27_,data_int_o_4__26_,data_int_o_4__25_,data_int_o_4__24_,
  data_int_o_4__23_,data_int_o_4__22_,data_int_o_4__21_,data_int_o_4__20_,
  data_int_o_4__19_,data_int_o_4__18_,data_int_o_4__17_,data_int_o_4__16_,data_int_o_4__15_,
  data_int_o_4__14_,data_int_o_4__13_,data_int_o_4__12_,data_int_o_4__11_,
  data_int_o_4__10_,data_int_o_4__9_,data_int_o_4__8_,data_int_o_4__7_,data_int_o_4__6_,
  data_int_o_4__5_,data_int_o_4__4_,data_int_o_4__3_,data_int_o_4__2_,
  data_int_o_4__1_,data_int_o_4__0_,N108,N109,N110,N111,data_head_9__159_,data_head_9__158_,
  data_head_9__157_,data_head_9__156_,data_head_9__155_,data_head_9__154_,
  data_head_9__153_,data_head_9__152_,data_head_9__151_,data_head_9__150_,data_head_9__149_,
  data_head_9__148_,data_head_9__147_,data_head_9__146_,data_head_9__145_,
  data_head_9__144_,data_head_9__143_,data_head_9__142_,data_head_9__141_,data_head_9__140_,
  data_head_9__139_,data_head_9__138_,data_head_9__137_,data_head_9__136_,
  data_head_9__135_,data_head_9__134_,data_head_9__133_,data_head_9__132_,
  data_head_9__131_,data_head_9__130_,data_head_9__129_,data_head_9__128_,data_head_9__127_,
  data_head_9__126_,data_head_9__125_,data_head_9__124_,data_head_9__123_,
  data_head_9__122_,data_head_9__121_,data_head_9__120_,data_head_9__119_,data_head_9__118_,
  data_head_9__117_,data_head_9__116_,data_head_9__115_,data_head_9__114_,
  data_head_9__113_,data_head_9__112_,data_head_9__111_,data_head_9__110_,data_head_9__109_,
  data_head_9__108_,data_head_9__107_,data_head_9__106_,data_head_9__105_,
  data_head_9__104_,data_head_9__103_,data_head_9__102_,data_head_9__101_,data_head_9__100_,
  data_head_9__99_,data_head_9__98_,data_head_9__97_,data_head_9__96_,
  data_head_9__95_,data_head_9__94_,data_head_9__93_,data_head_9__92_,data_head_9__91_,
  data_head_9__90_,data_head_9__89_,data_head_9__88_,data_head_9__87_,data_head_9__86_,
  data_head_9__85_,data_head_9__84_,data_head_9__83_,data_head_9__82_,
  data_head_9__81_,data_head_9__80_,data_head_9__79_,data_head_9__78_,data_head_9__77_,
  data_head_9__76_,data_head_9__75_,data_head_9__74_,data_head_9__73_,data_head_9__72_,
  data_head_9__71_,data_head_9__70_,data_head_9__69_,data_head_9__68_,
  data_head_9__67_,data_head_9__66_,data_head_9__65_,data_head_9__64_,data_head_9__63_,
  data_head_9__62_,data_head_9__61_,data_head_9__60_,data_head_9__59_,data_head_9__58_,
  data_head_9__57_,data_head_9__56_,data_head_9__55_,data_head_9__54_,data_head_9__53_,
  data_head_9__52_,data_head_9__51_,data_head_9__50_,data_head_9__49_,
  data_head_9__48_,data_head_9__47_,data_head_9__46_,data_head_9__45_,data_head_9__44_,
  data_head_9__43_,data_head_9__42_,data_head_9__41_,data_head_9__40_,data_head_9__39_,
  data_head_9__38_,data_head_9__37_,data_head_9__36_,data_head_9__35_,
  data_head_9__34_,data_head_9__33_,data_head_9__32_,data_head_9__31_,data_head_9__30_,
  data_head_9__29_,data_head_9__28_,data_head_9__27_,data_head_9__26_,data_head_9__25_,
  data_head_9__24_,data_head_9__23_,data_head_9__22_,data_head_9__21_,data_head_9__20_,
  data_head_9__19_,data_head_9__18_,data_head_9__17_,data_head_9__16_,
  data_head_9__15_,data_head_9__14_,data_head_9__13_,data_head_9__12_,data_head_9__11_,
  data_head_9__10_,data_head_9__9_,data_head_9__8_,data_head_9__7_,data_head_9__6_,
  data_head_9__5_,data_head_9__4_,data_head_9__3_,data_head_9__2_,data_head_9__1_,
  data_head_9__0_,_0_net_,valid_head_9__4_,valid_head_9__3_,valid_head_9__2_,
  valid_head_9__1_,valid_head_9__0_,_2_net__4_,_2_net__3_,_2_net__2_,_2_net__1_,_2_net__0_,
  _3_net__4_,_3_net__3_,_3_net__2_,_3_net__1_,_3_net__0_,ready_head_4__4_,
  ready_head_4__3_,ready_head_4__2_,ready_head_4__1_,ready_head_4__0_,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,_4_net__159_,_4_net__158_,_4_net__157_,_4_net__156_,
  _4_net__155_,_4_net__154_,_4_net__153_,_4_net__152_,_4_net__151_,_4_net__150_,
  _4_net__149_,_4_net__148_,_4_net__147_,_4_net__146_,_4_net__145_,_4_net__144_,
  _4_net__143_,_4_net__142_,_4_net__141_,_4_net__140_,_4_net__139_,_4_net__138_,
  _4_net__137_,_4_net__136_,_4_net__135_,_4_net__134_,_4_net__133_,_4_net__132_,
  _4_net__131_,_4_net__130_,_4_net__129_,_4_net__128_,_4_net__127_,_4_net__126_,
  _4_net__125_,_4_net__124_,_4_net__123_,_4_net__122_,_4_net__121_,_4_net__120_,
  _4_net__119_,_4_net__118_,_4_net__117_,_4_net__116_,_4_net__115_,_4_net__114_,_4_net__113_,
  _4_net__112_,_4_net__111_,_4_net__110_,_4_net__109_,_4_net__108_,_4_net__107_,
  _4_net__106_,_4_net__105_,_4_net__104_,_4_net__103_,_4_net__102_,_4_net__101_,
  _4_net__100_,_4_net__99_,_4_net__98_,_4_net__97_,_4_net__96_,_4_net__95_,_4_net__94_,
  _4_net__93_,_4_net__92_,_4_net__91_,_4_net__90_,_4_net__89_,_4_net__88_,
  _4_net__87_,_4_net__86_,_4_net__85_,_4_net__84_,_4_net__83_,_4_net__82_,_4_net__81_,
  _4_net__80_,_4_net__79_,_4_net__78_,_4_net__77_,_4_net__76_,_4_net__75_,_4_net__74_,
  _4_net__73_,_4_net__72_,_4_net__71_,_4_net__70_,_4_net__69_,_4_net__68_,
  _4_net__67_,_4_net__66_,_4_net__65_,_4_net__64_,_4_net__63_,_4_net__62_,_4_net__61_,
  _4_net__60_,_4_net__59_,_4_net__58_,_4_net__57_,_4_net__56_,_4_net__55_,_4_net__54_,
  _4_net__53_,_4_net__52_,_4_net__51_,_4_net__50_,_4_net__49_,_4_net__48_,
  _4_net__47_,_4_net__46_,_4_net__45_,_4_net__44_,_4_net__43_,_4_net__42_,_4_net__41_,
  _4_net__40_,_4_net__39_,_4_net__38_,_4_net__37_,_4_net__36_,_4_net__35_,_4_net__34_,
  _4_net__33_,_4_net__32_,_4_net__31_,_4_net__30_,_4_net__29_,_4_net__28_,
  _4_net__27_,_4_net__26_,_4_net__25_,_4_net__24_,_4_net__23_,_4_net__22_,_4_net__21_,
  _4_net__20_,_4_net__19_,_4_net__18_,_4_net__17_,_4_net__16_,_4_net__15_,_4_net__14_,
  _4_net__13_,_4_net__12_,_4_net__11_,_4_net__10_,_4_net__9_,_4_net__8_,
  _4_net__7_,_4_net__6_,_4_net__5_,_4_net__4_,_4_net__3_,_4_net__2_,_4_net__1_,_4_net__0_,
  N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,_5_net_,N132,N133,N134,N135,
  N136,N137,N138,N139;
  wire [2:0] go_cnt;

  bsg_make_2D_array_width_p32_items_p5
  bm2Da
  (
    .i(data_o_flat),
    .o(data_o)
  );


  bsg_rr_f2f_input_width_p32_num_in_p10_middle_meet_p5
  \ic_9_.in_chan.bsg_rr_ff_in 
  (
    .clk(clk),
    .reset(_0_net_),
    .valid_i(valid_i),
    .data_i(data_i),
    .data_head_o({ data_head_9__159_, data_head_9__158_, data_head_9__157_, data_head_9__156_, data_head_9__155_, data_head_9__154_, data_head_9__153_, data_head_9__152_, data_head_9__151_, data_head_9__150_, data_head_9__149_, data_head_9__148_, data_head_9__147_, data_head_9__146_, data_head_9__145_, data_head_9__144_, data_head_9__143_, data_head_9__142_, data_head_9__141_, data_head_9__140_, data_head_9__139_, data_head_9__138_, data_head_9__137_, data_head_9__136_, data_head_9__135_, data_head_9__134_, data_head_9__133_, data_head_9__132_, data_head_9__131_, data_head_9__130_, data_head_9__129_, data_head_9__128_, data_head_9__127_, data_head_9__126_, data_head_9__125_, data_head_9__124_, data_head_9__123_, data_head_9__122_, data_head_9__121_, data_head_9__120_, data_head_9__119_, data_head_9__118_, data_head_9__117_, data_head_9__116_, data_head_9__115_, data_head_9__114_, data_head_9__113_, data_head_9__112_, data_head_9__111_, data_head_9__110_, data_head_9__109_, data_head_9__108_, data_head_9__107_, data_head_9__106_, data_head_9__105_, data_head_9__104_, data_head_9__103_, data_head_9__102_, data_head_9__101_, data_head_9__100_, data_head_9__99_, data_head_9__98_, data_head_9__97_, data_head_9__96_, data_head_9__95_, data_head_9__94_, data_head_9__93_, data_head_9__92_, data_head_9__91_, data_head_9__90_, data_head_9__89_, data_head_9__88_, data_head_9__87_, data_head_9__86_, data_head_9__85_, data_head_9__84_, data_head_9__83_, data_head_9__82_, data_head_9__81_, data_head_9__80_, data_head_9__79_, data_head_9__78_, data_head_9__77_, data_head_9__76_, data_head_9__75_, data_head_9__74_, data_head_9__73_, data_head_9__72_, data_head_9__71_, data_head_9__70_, data_head_9__69_, data_head_9__68_, data_head_9__67_, data_head_9__66_, data_head_9__65_, data_head_9__64_, data_head_9__63_, data_head_9__62_, data_head_9__61_, data_head_9__60_, data_head_9__59_, data_head_9__58_, data_head_9__57_, data_head_9__56_, data_head_9__55_, data_head_9__54_, data_head_9__53_, data_head_9__52_, data_head_9__51_, data_head_9__50_, data_head_9__49_, data_head_9__48_, data_head_9__47_, data_head_9__46_, data_head_9__45_, data_head_9__44_, data_head_9__43_, data_head_9__42_, data_head_9__41_, data_head_9__40_, data_head_9__39_, data_head_9__38_, data_head_9__37_, data_head_9__36_, data_head_9__35_, data_head_9__34_, data_head_9__33_, data_head_9__32_, data_head_9__31_, data_head_9__30_, data_head_9__29_, data_head_9__28_, data_head_9__27_, data_head_9__26_, data_head_9__25_, data_head_9__24_, data_head_9__23_, data_head_9__22_, data_head_9__21_, data_head_9__20_, data_head_9__19_, data_head_9__18_, data_head_9__17_, data_head_9__16_, data_head_9__15_, data_head_9__14_, data_head_9__13_, data_head_9__12_, data_head_9__11_, data_head_9__10_, data_head_9__9_, data_head_9__8_, data_head_9__7_, data_head_9__6_, data_head_9__5_, data_head_9__4_, data_head_9__3_, data_head_9__2_, data_head_9__1_, data_head_9__0_ }),
    .valid_head_o({ valid_head_9__4_, valid_head_9__3_, valid_head_9__2_, valid_head_9__1_, valid_head_9__0_ }),
    .go_channels_i(go_channels),
    .go_cnt_i(go_cnt),
    .yumi_o({ yumi_int_o_9__9_, yumi_int_o_9__8_, yumi_int_o_9__7_, yumi_int_o_9__6_, yumi_int_o_9__5_, yumi_int_o_9__4_, yumi_int_o_9__3_, yumi_int_o_9__2_, yumi_int_o_9__1_, yumi_int_o_9__0_ })
  );


  bsg_rr_f2f_middle_width_p32_middle_meet_p5
  brrf2fm
  (
    .valid_head_i({ _2_net__4_, _2_net__3_, _2_net__2_, _2_net__1_, _2_net__0_ }),
    .ready_head_i({ _3_net__4_, _3_net__3_, _3_net__2_, _3_net__1_, _3_net__0_ }),
    .go_channels_o(go_channels),
    .go_cnt_o(go_cnt)
  );


  bsg_make_2D_array_width_p32_items_p5
  \oc_4_.out_chan.bm2Da 
  (
    .i({ _4_net__159_, _4_net__158_, _4_net__157_, _4_net__156_, _4_net__155_, _4_net__154_, _4_net__153_, _4_net__152_, _4_net__151_, _4_net__150_, _4_net__149_, _4_net__148_, _4_net__147_, _4_net__146_, _4_net__145_, _4_net__144_, _4_net__143_, _4_net__142_, _4_net__141_, _4_net__140_, _4_net__139_, _4_net__138_, _4_net__137_, _4_net__136_, _4_net__135_, _4_net__134_, _4_net__133_, _4_net__132_, _4_net__131_, _4_net__130_, _4_net__129_, _4_net__128_, _4_net__127_, _4_net__126_, _4_net__125_, _4_net__124_, _4_net__123_, _4_net__122_, _4_net__121_, _4_net__120_, _4_net__119_, _4_net__118_, _4_net__117_, _4_net__116_, _4_net__115_, _4_net__114_, _4_net__113_, _4_net__112_, _4_net__111_, _4_net__110_, _4_net__109_, _4_net__108_, _4_net__107_, _4_net__106_, _4_net__105_, _4_net__104_, _4_net__103_, _4_net__102_, _4_net__101_, _4_net__100_, _4_net__99_, _4_net__98_, _4_net__97_, _4_net__96_, _4_net__95_, _4_net__94_, _4_net__93_, _4_net__92_, _4_net__91_, _4_net__90_, _4_net__89_, _4_net__88_, _4_net__87_, _4_net__86_, _4_net__85_, _4_net__84_, _4_net__83_, _4_net__82_, _4_net__81_, _4_net__80_, _4_net__79_, _4_net__78_, _4_net__77_, _4_net__76_, _4_net__75_, _4_net__74_, _4_net__73_, _4_net__72_, _4_net__71_, _4_net__70_, _4_net__69_, _4_net__68_, _4_net__67_, _4_net__66_, _4_net__65_, _4_net__64_, _4_net__63_, _4_net__62_, _4_net__61_, _4_net__60_, _4_net__59_, _4_net__58_, _4_net__57_, _4_net__56_, _4_net__55_, _4_net__54_, _4_net__53_, _4_net__52_, _4_net__51_, _4_net__50_, _4_net__49_, _4_net__48_, _4_net__47_, _4_net__46_, _4_net__45_, _4_net__44_, _4_net__43_, _4_net__42_, _4_net__41_, _4_net__40_, _4_net__39_, _4_net__38_, _4_net__37_, _4_net__36_, _4_net__35_, _4_net__34_, _4_net__33_, _4_net__32_, _4_net__31_, _4_net__30_, _4_net__29_, _4_net__28_, _4_net__27_, _4_net__26_, _4_net__25_, _4_net__24_, _4_net__23_, _4_net__22_, _4_net__21_, _4_net__20_, _4_net__19_, _4_net__18_, _4_net__17_, _4_net__16_, _4_net__15_, _4_net__14_, _4_net__13_, _4_net__12_, _4_net__11_, _4_net__10_, _4_net__9_, _4_net__8_, _4_net__7_, _4_net__6_, _4_net__5_, _4_net__4_, _4_net__3_, _4_net__2_, _4_net__1_, _4_net__0_ }),
    .o(\oc_4_.out_chan.data_head_array )
  );


  bsg_rr_f2f_output_width_p32_num_out_p5_middle_meet_p5
  \oc_4_.out_chan.bsg_rr_ff_out 
  (
    .clk(clk),
    .reset(_5_net_),
    .ready_i(ready_i),
    .ready_head_o({ ready_head_4__4_, ready_head_4__3_, ready_head_4__2_, ready_head_4__1_, ready_head_4__0_ }),
    .go_channels_i(go_channels),
    .go_cnt_i(go_cnt),
    .data_head_i(\oc_4_.out_chan.data_head_array ),
    .valid_o({ valid_int_o_4__4_, valid_int_o_4__3_, valid_int_o_4__2_, valid_int_o_4__1_, valid_int_o_4__0_ }),
    .data_o({ data_int_o_4__159_, data_int_o_4__158_, data_int_o_4__157_, data_int_o_4__156_, data_int_o_4__155_, data_int_o_4__154_, data_int_o_4__153_, data_int_o_4__152_, data_int_o_4__151_, data_int_o_4__150_, data_int_o_4__149_, data_int_o_4__148_, data_int_o_4__147_, data_int_o_4__146_, data_int_o_4__145_, data_int_o_4__144_, data_int_o_4__143_, data_int_o_4__142_, data_int_o_4__141_, data_int_o_4__140_, data_int_o_4__139_, data_int_o_4__138_, data_int_o_4__137_, data_int_o_4__136_, data_int_o_4__135_, data_int_o_4__134_, data_int_o_4__133_, data_int_o_4__132_, data_int_o_4__131_, data_int_o_4__130_, data_int_o_4__129_, data_int_o_4__128_, data_int_o_4__127_, data_int_o_4__126_, data_int_o_4__125_, data_int_o_4__124_, data_int_o_4__123_, data_int_o_4__122_, data_int_o_4__121_, data_int_o_4__120_, data_int_o_4__119_, data_int_o_4__118_, data_int_o_4__117_, data_int_o_4__116_, data_int_o_4__115_, data_int_o_4__114_, data_int_o_4__113_, data_int_o_4__112_, data_int_o_4__111_, data_int_o_4__110_, data_int_o_4__109_, data_int_o_4__108_, data_int_o_4__107_, data_int_o_4__106_, data_int_o_4__105_, data_int_o_4__104_, data_int_o_4__103_, data_int_o_4__102_, data_int_o_4__101_, data_int_o_4__100_, data_int_o_4__99_, data_int_o_4__98_, data_int_o_4__97_, data_int_o_4__96_, data_int_o_4__95_, data_int_o_4__94_, data_int_o_4__93_, data_int_o_4__92_, data_int_o_4__91_, data_int_o_4__90_, data_int_o_4__89_, data_int_o_4__88_, data_int_o_4__87_, data_int_o_4__86_, data_int_o_4__85_, data_int_o_4__84_, data_int_o_4__83_, data_int_o_4__82_, data_int_o_4__81_, data_int_o_4__80_, data_int_o_4__79_, data_int_o_4__78_, data_int_o_4__77_, data_int_o_4__76_, data_int_o_4__75_, data_int_o_4__74_, data_int_o_4__73_, data_int_o_4__72_, data_int_o_4__71_, data_int_o_4__70_, data_int_o_4__69_, data_int_o_4__68_, data_int_o_4__67_, data_int_o_4__66_, data_int_o_4__65_, data_int_o_4__64_, data_int_o_4__63_, data_int_o_4__62_, data_int_o_4__61_, data_int_o_4__60_, data_int_o_4__59_, data_int_o_4__58_, data_int_o_4__57_, data_int_o_4__56_, data_int_o_4__55_, data_int_o_4__54_, data_int_o_4__53_, data_int_o_4__52_, data_int_o_4__51_, data_int_o_4__50_, data_int_o_4__49_, data_int_o_4__48_, data_int_o_4__47_, data_int_o_4__46_, data_int_o_4__45_, data_int_o_4__44_, data_int_o_4__43_, data_int_o_4__42_, data_int_o_4__41_, data_int_o_4__40_, data_int_o_4__39_, data_int_o_4__38_, data_int_o_4__37_, data_int_o_4__36_, data_int_o_4__35_, data_int_o_4__34_, data_int_o_4__33_, data_int_o_4__32_, data_int_o_4__31_, data_int_o_4__30_, data_int_o_4__29_, data_int_o_4__28_, data_int_o_4__27_, data_int_o_4__26_, data_int_o_4__25_, data_int_o_4__24_, data_int_o_4__23_, data_int_o_4__22_, data_int_o_4__21_, data_int_o_4__20_, data_int_o_4__19_, data_int_o_4__18_, data_int_o_4__17_, data_int_o_4__16_, data_int_o_4__15_, data_int_o_4__14_, data_int_o_4__13_, data_int_o_4__12_, data_int_o_4__11_, data_int_o_4__10_, data_int_o_4__9_, data_int_o_4__8_, data_int_o_4__7_, data_int_o_4__6_, data_int_o_4__5_, data_int_o_4__4_, data_int_o_4__3_, data_int_o_4__2_, data_int_o_4__1_, data_int_o_4__0_ })
  );

  assign N132 = ~in_top_channel_i[3];
  assign N133 = ~in_top_channel_i[0];
  assign N134 = in_top_channel_i[2] | N132;
  assign N135 = in_top_channel_i[1] | N134;
  assign N136 = N133 | N135;
  assign N137 = ~out_top_channel_i[2];
  assign N138 = out_top_channel_i[1] | N137;
  assign N139 = out_top_channel_i[0] | N138;
  assign N104 = N0 & N1 & N2;
  assign N0 = ~out_top_channel_i[2];
  assign N1 = ~out_top_channel_i[0];
  assign N2 = ~out_top_channel_i[1];
  assign N105 = out_top_channel_i[0] & N3;
  assign N3 = ~out_top_channel_i[1];
  assign N106 = N4 & out_top_channel_i[1];
  assign N4 = ~out_top_channel_i[0];
  assign N107 = out_top_channel_i[0] & out_top_channel_i[1];
  assign N108 = N5 & N6 & N7;
  assign N5 = ~out_top_channel_i[2];
  assign N6 = ~out_top_channel_i[0];
  assign N7 = ~out_top_channel_i[1];
  assign N109 = out_top_channel_i[0] & N8;
  assign N8 = ~out_top_channel_i[1];
  assign N110 = N9 & out_top_channel_i[1];
  assign N9 = ~out_top_channel_i[0];
  assign N111 = out_top_channel_i[0] & out_top_channel_i[1];
  assign N94 = N10 & N11 & (N12 & N13);
  assign N10 = ~in_top_channel_i[3];
  assign N11 = ~in_top_channel_i[2];
  assign N12 = ~in_top_channel_i[0];
  assign N13 = ~in_top_channel_i[1];
  assign N95 = in_top_channel_i[3] & N14;
  assign N14 = ~in_top_channel_i[0];
  assign N96 = N15 & N16 & (in_top_channel_i[0] & N17);
  assign N15 = ~in_top_channel_i[3];
  assign N16 = ~in_top_channel_i[2];
  assign N17 = ~in_top_channel_i[1];
  assign N98 = N18 & N19 & in_top_channel_i[1];
  assign N18 = ~in_top_channel_i[2];
  assign N19 = ~in_top_channel_i[0];
  assign N99 = N20 & in_top_channel_i[0] & in_top_channel_i[1];
  assign N20 = ~in_top_channel_i[2];
  assign N100 = in_top_channel_i[2] & N21 & N22;
  assign N21 = ~in_top_channel_i[0];
  assign N22 = ~in_top_channel_i[1];
  assign N101 = in_top_channel_i[2] & in_top_channel_i[0] & N23;
  assign N23 = ~in_top_channel_i[1];
  assign N102 = in_top_channel_i[2] & N24 & in_top_channel_i[1];
  assign N24 = ~in_top_channel_i[0];
  assign N103 = in_top_channel_i[2] & in_top_channel_i[0] & in_top_channel_i[1];
  assign N97 = in_top_channel_i[3] & in_top_channel_i[0];
  assign N112 = N25 & N26 & (N27 & N28);
  assign N25 = ~in_top_channel_i[3];
  assign N26 = ~in_top_channel_i[2];
  assign N27 = ~in_top_channel_i[0];
  assign N28 = ~in_top_channel_i[1];
  assign N113 = in_top_channel_i[3] & N29;
  assign N29 = ~in_top_channel_i[0];
  assign N114 = N30 & N31 & (in_top_channel_i[0] & N32);
  assign N30 = ~in_top_channel_i[3];
  assign N31 = ~in_top_channel_i[2];
  assign N32 = ~in_top_channel_i[1];
  assign N116 = N33 & N34 & in_top_channel_i[1];
  assign N33 = ~in_top_channel_i[2];
  assign N34 = ~in_top_channel_i[0];
  assign N117 = N35 & in_top_channel_i[0] & in_top_channel_i[1];
  assign N35 = ~in_top_channel_i[2];
  assign N118 = in_top_channel_i[2] & N36 & N37;
  assign N36 = ~in_top_channel_i[0];
  assign N37 = ~in_top_channel_i[1];
  assign N119 = in_top_channel_i[2] & in_top_channel_i[0] & N38;
  assign N38 = ~in_top_channel_i[1];
  assign N120 = in_top_channel_i[2] & N39 & in_top_channel_i[1];
  assign N39 = ~in_top_channel_i[0];
  assign N121 = in_top_channel_i[2] & in_top_channel_i[0] & in_top_channel_i[1];
  assign N115 = in_top_channel_i[3] & in_top_channel_i[0];
  assign N122 = N40 & N41 & (N42 & N43);
  assign N40 = ~in_top_channel_i[3];
  assign N41 = ~in_top_channel_i[2];
  assign N42 = ~in_top_channel_i[0];
  assign N43 = ~in_top_channel_i[1];
  assign N123 = in_top_channel_i[3] & N44;
  assign N44 = ~in_top_channel_i[0];
  assign N124 = N45 & N46 & (in_top_channel_i[0] & N47);
  assign N45 = ~in_top_channel_i[3];
  assign N46 = ~in_top_channel_i[2];
  assign N47 = ~in_top_channel_i[1];
  assign N126 = N48 & N49 & in_top_channel_i[1];
  assign N48 = ~in_top_channel_i[2];
  assign N49 = ~in_top_channel_i[0];
  assign N127 = N50 & in_top_channel_i[0] & in_top_channel_i[1];
  assign N50 = ~in_top_channel_i[2];
  assign N128 = in_top_channel_i[2] & N51 & N52;
  assign N51 = ~in_top_channel_i[0];
  assign N52 = ~in_top_channel_i[1];
  assign N129 = in_top_channel_i[2] & in_top_channel_i[0] & N53;
  assign N53 = ~in_top_channel_i[1];
  assign N130 = in_top_channel_i[2] & N54 & in_top_channel_i[1];
  assign N54 = ~in_top_channel_i[0];
  assign N131 = in_top_channel_i[2] & in_top_channel_i[0] & in_top_channel_i[1];
  assign N125 = in_top_channel_i[3] & in_top_channel_i[0];
  assign valid_o[4] = (N55)? 1'b0 : 
                      (N56)? 1'b0 : 
                      (N57)? 1'b0 : 
                      (N58)? 1'b0 : 
                      (N59)? valid_int_o_4__4_ : 1'b0;
  assign N55 = N104;
  assign N56 = N105;
  assign N57 = N106;
  assign N58 = N107;
  assign N59 = out_top_channel_i[2];
  assign valid_o[3] = (N55)? 1'b0 : 
                      (N56)? 1'b0 : 
                      (N57)? 1'b0 : 
                      (N58)? 1'b0 : 
                      (N59)? valid_int_o_4__3_ : 1'b0;
  assign valid_o[2] = (N55)? 1'b0 : 
                      (N56)? 1'b0 : 
                      (N57)? 1'b0 : 
                      (N58)? 1'b0 : 
                      (N59)? valid_int_o_4__2_ : 1'b0;
  assign valid_o[1] = (N55)? 1'b0 : 
                      (N56)? 1'b0 : 
                      (N57)? 1'b0 : 
                      (N58)? 1'b0 : 
                      (N59)? valid_int_o_4__1_ : 1'b0;
  assign valid_o[0] = (N55)? 1'b0 : 
                      (N56)? 1'b0 : 
                      (N57)? 1'b0 : 
                      (N58)? 1'b0 : 
                      (N59)? valid_int_o_4__0_ : 1'b0;
  assign data_o_flat[159] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__159_ : 1'b0;
  assign N60 = N108;
  assign N61 = N109;
  assign N62 = N110;
  assign N63 = N111;
  assign data_o_flat[158] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__158_ : 1'b0;
  assign data_o_flat[157] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__157_ : 1'b0;
  assign data_o_flat[156] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__156_ : 1'b0;
  assign data_o_flat[155] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__155_ : 1'b0;
  assign data_o_flat[154] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__154_ : 1'b0;
  assign data_o_flat[153] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__153_ : 1'b0;
  assign data_o_flat[152] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__152_ : 1'b0;
  assign data_o_flat[151] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__151_ : 1'b0;
  assign data_o_flat[150] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__150_ : 1'b0;
  assign data_o_flat[149] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__149_ : 1'b0;
  assign data_o_flat[148] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__148_ : 1'b0;
  assign data_o_flat[147] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__147_ : 1'b0;
  assign data_o_flat[146] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__146_ : 1'b0;
  assign data_o_flat[145] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__145_ : 1'b0;
  assign data_o_flat[144] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__144_ : 1'b0;
  assign data_o_flat[143] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__143_ : 1'b0;
  assign data_o_flat[142] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__142_ : 1'b0;
  assign data_o_flat[141] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__141_ : 1'b0;
  assign data_o_flat[140] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__140_ : 1'b0;
  assign data_o_flat[139] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__139_ : 1'b0;
  assign data_o_flat[138] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__138_ : 1'b0;
  assign data_o_flat[137] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__137_ : 1'b0;
  assign data_o_flat[136] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__136_ : 1'b0;
  assign data_o_flat[135] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__135_ : 1'b0;
  assign data_o_flat[134] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__134_ : 1'b0;
  assign data_o_flat[133] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__133_ : 1'b0;
  assign data_o_flat[132] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__132_ : 1'b0;
  assign data_o_flat[131] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__131_ : 1'b0;
  assign data_o_flat[130] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__130_ : 1'b0;
  assign data_o_flat[129] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__129_ : 1'b0;
  assign data_o_flat[128] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__128_ : 1'b0;
  assign data_o_flat[127] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__127_ : 1'b0;
  assign data_o_flat[126] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__126_ : 1'b0;
  assign data_o_flat[125] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__125_ : 1'b0;
  assign data_o_flat[124] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__124_ : 1'b0;
  assign data_o_flat[123] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__123_ : 1'b0;
  assign data_o_flat[122] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__122_ : 1'b0;
  assign data_o_flat[121] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__121_ : 1'b0;
  assign data_o_flat[120] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__120_ : 1'b0;
  assign data_o_flat[119] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__119_ : 1'b0;
  assign data_o_flat[118] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__118_ : 1'b0;
  assign data_o_flat[117] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__117_ : 1'b0;
  assign data_o_flat[116] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__116_ : 1'b0;
  assign data_o_flat[115] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__115_ : 1'b0;
  assign data_o_flat[114] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__114_ : 1'b0;
  assign data_o_flat[113] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__113_ : 1'b0;
  assign data_o_flat[112] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__112_ : 1'b0;
  assign data_o_flat[111] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__111_ : 1'b0;
  assign data_o_flat[110] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__110_ : 1'b0;
  assign data_o_flat[109] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__109_ : 1'b0;
  assign data_o_flat[108] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__108_ : 1'b0;
  assign data_o_flat[107] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__107_ : 1'b0;
  assign data_o_flat[106] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__106_ : 1'b0;
  assign data_o_flat[105] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__105_ : 1'b0;
  assign data_o_flat[104] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__104_ : 1'b0;
  assign data_o_flat[103] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__103_ : 1'b0;
  assign data_o_flat[102] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__102_ : 1'b0;
  assign data_o_flat[101] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__101_ : 1'b0;
  assign data_o_flat[100] = (N60)? 1'b0 : 
                            (N61)? 1'b0 : 
                            (N62)? 1'b0 : 
                            (N63)? 1'b0 : 
                            (N59)? data_int_o_4__100_ : 1'b0;
  assign data_o_flat[99] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__99_ : 1'b0;
  assign data_o_flat[98] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__98_ : 1'b0;
  assign data_o_flat[97] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__97_ : 1'b0;
  assign data_o_flat[96] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__96_ : 1'b0;
  assign data_o_flat[95] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__95_ : 1'b0;
  assign data_o_flat[94] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__94_ : 1'b0;
  assign data_o_flat[93] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__93_ : 1'b0;
  assign data_o_flat[92] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__92_ : 1'b0;
  assign data_o_flat[91] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__91_ : 1'b0;
  assign data_o_flat[90] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__90_ : 1'b0;
  assign data_o_flat[89] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__89_ : 1'b0;
  assign data_o_flat[88] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__88_ : 1'b0;
  assign data_o_flat[87] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__87_ : 1'b0;
  assign data_o_flat[86] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__86_ : 1'b0;
  assign data_o_flat[85] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__85_ : 1'b0;
  assign data_o_flat[84] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__84_ : 1'b0;
  assign data_o_flat[83] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__83_ : 1'b0;
  assign data_o_flat[82] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__82_ : 1'b0;
  assign data_o_flat[81] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__81_ : 1'b0;
  assign data_o_flat[80] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__80_ : 1'b0;
  assign data_o_flat[79] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__79_ : 1'b0;
  assign data_o_flat[78] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__78_ : 1'b0;
  assign data_o_flat[77] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__77_ : 1'b0;
  assign data_o_flat[76] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__76_ : 1'b0;
  assign data_o_flat[75] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__75_ : 1'b0;
  assign data_o_flat[74] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__74_ : 1'b0;
  assign data_o_flat[73] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__73_ : 1'b0;
  assign data_o_flat[72] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__72_ : 1'b0;
  assign data_o_flat[71] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__71_ : 1'b0;
  assign data_o_flat[70] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__70_ : 1'b0;
  assign data_o_flat[69] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__69_ : 1'b0;
  assign data_o_flat[68] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__68_ : 1'b0;
  assign data_o_flat[67] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__67_ : 1'b0;
  assign data_o_flat[66] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__66_ : 1'b0;
  assign data_o_flat[65] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__65_ : 1'b0;
  assign data_o_flat[64] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__64_ : 1'b0;
  assign data_o_flat[63] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__63_ : 1'b0;
  assign data_o_flat[62] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__62_ : 1'b0;
  assign data_o_flat[61] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__61_ : 1'b0;
  assign data_o_flat[60] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__60_ : 1'b0;
  assign data_o_flat[59] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__59_ : 1'b0;
  assign data_o_flat[58] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__58_ : 1'b0;
  assign data_o_flat[57] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__57_ : 1'b0;
  assign data_o_flat[56] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__56_ : 1'b0;
  assign data_o_flat[55] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__55_ : 1'b0;
  assign data_o_flat[54] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__54_ : 1'b0;
  assign data_o_flat[53] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__53_ : 1'b0;
  assign data_o_flat[52] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__52_ : 1'b0;
  assign data_o_flat[51] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__51_ : 1'b0;
  assign data_o_flat[50] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__50_ : 1'b0;
  assign data_o_flat[49] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__49_ : 1'b0;
  assign data_o_flat[48] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__48_ : 1'b0;
  assign data_o_flat[47] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__47_ : 1'b0;
  assign data_o_flat[46] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__46_ : 1'b0;
  assign data_o_flat[45] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__45_ : 1'b0;
  assign data_o_flat[44] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__44_ : 1'b0;
  assign data_o_flat[43] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__43_ : 1'b0;
  assign data_o_flat[42] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__42_ : 1'b0;
  assign data_o_flat[41] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__41_ : 1'b0;
  assign data_o_flat[40] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__40_ : 1'b0;
  assign data_o_flat[39] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__39_ : 1'b0;
  assign data_o_flat[38] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__38_ : 1'b0;
  assign data_o_flat[37] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__37_ : 1'b0;
  assign data_o_flat[36] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__36_ : 1'b0;
  assign data_o_flat[35] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__35_ : 1'b0;
  assign data_o_flat[34] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__34_ : 1'b0;
  assign data_o_flat[33] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__33_ : 1'b0;
  assign data_o_flat[32] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__32_ : 1'b0;
  assign data_o_flat[31] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__31_ : 1'b0;
  assign data_o_flat[30] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__30_ : 1'b0;
  assign data_o_flat[29] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__29_ : 1'b0;
  assign data_o_flat[28] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__28_ : 1'b0;
  assign data_o_flat[27] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__27_ : 1'b0;
  assign data_o_flat[26] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__26_ : 1'b0;
  assign data_o_flat[25] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__25_ : 1'b0;
  assign data_o_flat[24] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__24_ : 1'b0;
  assign data_o_flat[23] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__23_ : 1'b0;
  assign data_o_flat[22] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__22_ : 1'b0;
  assign data_o_flat[21] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__21_ : 1'b0;
  assign data_o_flat[20] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__20_ : 1'b0;
  assign data_o_flat[19] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__19_ : 1'b0;
  assign data_o_flat[18] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__18_ : 1'b0;
  assign data_o_flat[17] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__17_ : 1'b0;
  assign data_o_flat[16] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__16_ : 1'b0;
  assign data_o_flat[15] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__15_ : 1'b0;
  assign data_o_flat[14] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__14_ : 1'b0;
  assign data_o_flat[13] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__13_ : 1'b0;
  assign data_o_flat[12] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__12_ : 1'b0;
  assign data_o_flat[11] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__11_ : 1'b0;
  assign data_o_flat[10] = (N60)? 1'b0 : 
                           (N61)? 1'b0 : 
                           (N62)? 1'b0 : 
                           (N63)? 1'b0 : 
                           (N59)? data_int_o_4__10_ : 1'b0;
  assign data_o_flat[9] = (N60)? 1'b0 : 
                          (N61)? 1'b0 : 
                          (N62)? 1'b0 : 
                          (N63)? 1'b0 : 
                          (N59)? data_int_o_4__9_ : 1'b0;
  assign data_o_flat[8] = (N60)? 1'b0 : 
                          (N61)? 1'b0 : 
                          (N62)? 1'b0 : 
                          (N63)? 1'b0 : 
                          (N59)? data_int_o_4__8_ : 1'b0;
  assign data_o_flat[7] = (N60)? 1'b0 : 
                          (N61)? 1'b0 : 
                          (N62)? 1'b0 : 
                          (N63)? 1'b0 : 
                          (N59)? data_int_o_4__7_ : 1'b0;
  assign data_o_flat[6] = (N60)? 1'b0 : 
                          (N61)? 1'b0 : 
                          (N62)? 1'b0 : 
                          (N63)? 1'b0 : 
                          (N59)? data_int_o_4__6_ : 1'b0;
  assign data_o_flat[5] = (N60)? 1'b0 : 
                          (N61)? 1'b0 : 
                          (N62)? 1'b0 : 
                          (N63)? 1'b0 : 
                          (N59)? data_int_o_4__5_ : 1'b0;
  assign data_o_flat[4] = (N60)? 1'b0 : 
                          (N61)? 1'b0 : 
                          (N62)? 1'b0 : 
                          (N63)? 1'b0 : 
                          (N59)? data_int_o_4__4_ : 1'b0;
  assign data_o_flat[3] = (N60)? 1'b0 : 
                          (N61)? 1'b0 : 
                          (N62)? 1'b0 : 
                          (N63)? 1'b0 : 
                          (N59)? data_int_o_4__3_ : 1'b0;
  assign data_o_flat[2] = (N60)? 1'b0 : 
                          (N61)? 1'b0 : 
                          (N62)? 1'b0 : 
                          (N63)? 1'b0 : 
                          (N59)? data_int_o_4__2_ : 1'b0;
  assign data_o_flat[1] = (N60)? 1'b0 : 
                          (N61)? 1'b0 : 
                          (N62)? 1'b0 : 
                          (N63)? 1'b0 : 
                          (N59)? data_int_o_4__1_ : 1'b0;
  assign data_o_flat[0] = (N60)? 1'b0 : 
                          (N61)? 1'b0 : 
                          (N62)? 1'b0 : 
                          (N63)? 1'b0 : 
                          (N59)? data_int_o_4__0_ : 1'b0;
  assign _3_net__4_ = (N55)? 1'b0 : 
                      (N56)? 1'b0 : 
                      (N57)? 1'b0 : 
                      (N58)? 1'b0 : 
                      (N59)? ready_head_4__4_ : 1'b0;
  assign _3_net__3_ = (N55)? 1'b0 : 
                      (N56)? 1'b0 : 
                      (N57)? 1'b0 : 
                      (N58)? 1'b0 : 
                      (N59)? ready_head_4__3_ : 1'b0;
  assign _3_net__2_ = (N55)? 1'b0 : 
                      (N56)? 1'b0 : 
                      (N57)? 1'b0 : 
                      (N58)? 1'b0 : 
                      (N59)? ready_head_4__2_ : 1'b0;
  assign _3_net__1_ = (N55)? 1'b0 : 
                      (N56)? 1'b0 : 
                      (N57)? 1'b0 : 
                      (N58)? 1'b0 : 
                      (N59)? ready_head_4__1_ : 1'b0;
  assign _3_net__0_ = (N55)? 1'b0 : 
                      (N56)? 1'b0 : 
                      (N57)? 1'b0 : 
                      (N58)? 1'b0 : 
                      (N59)? ready_head_4__0_ : 1'b0;
  assign yumi_o[9] = (N64)? 1'b0 : 
                     (N65)? 1'b0 : 
                     (N66)? 1'b0 : 
                     (N67)? 1'b0 : 
                     (N68)? 1'b0 : 
                     (N69)? 1'b0 : 
                     (N70)? 1'b0 : 
                     (N71)? 1'b0 : 
                     (N72)? 1'b0 : 
                     (N73)? yumi_int_o_9__9_ : 1'b0;
  assign N64 = N94;
  assign N65 = N96;
  assign N66 = N98;
  assign N67 = N99;
  assign N68 = N100;
  assign N69 = N101;
  assign N70 = N102;
  assign N71 = N103;
  assign N72 = N95;
  assign N73 = N97;
  assign yumi_o[8] = (N64)? 1'b0 : 
                     (N65)? 1'b0 : 
                     (N66)? 1'b0 : 
                     (N67)? 1'b0 : 
                     (N68)? 1'b0 : 
                     (N69)? 1'b0 : 
                     (N70)? 1'b0 : 
                     (N71)? 1'b0 : 
                     (N72)? 1'b0 : 
                     (N73)? yumi_int_o_9__8_ : 1'b0;
  assign yumi_o[7] = (N64)? 1'b0 : 
                     (N65)? 1'b0 : 
                     (N66)? 1'b0 : 
                     (N67)? 1'b0 : 
                     (N68)? 1'b0 : 
                     (N69)? 1'b0 : 
                     (N70)? 1'b0 : 
                     (N71)? 1'b0 : 
                     (N72)? 1'b0 : 
                     (N73)? yumi_int_o_9__7_ : 1'b0;
  assign yumi_o[6] = (N64)? 1'b0 : 
                     (N65)? 1'b0 : 
                     (N66)? 1'b0 : 
                     (N67)? 1'b0 : 
                     (N68)? 1'b0 : 
                     (N69)? 1'b0 : 
                     (N70)? 1'b0 : 
                     (N71)? 1'b0 : 
                     (N72)? 1'b0 : 
                     (N73)? yumi_int_o_9__6_ : 1'b0;
  assign yumi_o[5] = (N64)? 1'b0 : 
                     (N65)? 1'b0 : 
                     (N66)? 1'b0 : 
                     (N67)? 1'b0 : 
                     (N68)? 1'b0 : 
                     (N69)? 1'b0 : 
                     (N70)? 1'b0 : 
                     (N71)? 1'b0 : 
                     (N72)? 1'b0 : 
                     (N73)? yumi_int_o_9__5_ : 1'b0;
  assign yumi_o[4] = (N64)? 1'b0 : 
                     (N65)? 1'b0 : 
                     (N66)? 1'b0 : 
                     (N67)? 1'b0 : 
                     (N68)? 1'b0 : 
                     (N69)? 1'b0 : 
                     (N70)? 1'b0 : 
                     (N71)? 1'b0 : 
                     (N72)? 1'b0 : 
                     (N73)? yumi_int_o_9__4_ : 1'b0;
  assign yumi_o[3] = (N64)? 1'b0 : 
                     (N65)? 1'b0 : 
                     (N66)? 1'b0 : 
                     (N67)? 1'b0 : 
                     (N68)? 1'b0 : 
                     (N69)? 1'b0 : 
                     (N70)? 1'b0 : 
                     (N71)? 1'b0 : 
                     (N72)? 1'b0 : 
                     (N73)? yumi_int_o_9__3_ : 1'b0;
  assign yumi_o[2] = (N64)? 1'b0 : 
                     (N65)? 1'b0 : 
                     (N66)? 1'b0 : 
                     (N67)? 1'b0 : 
                     (N68)? 1'b0 : 
                     (N69)? 1'b0 : 
                     (N70)? 1'b0 : 
                     (N71)? 1'b0 : 
                     (N72)? 1'b0 : 
                     (N73)? yumi_int_o_9__2_ : 1'b0;
  assign yumi_o[1] = (N64)? 1'b0 : 
                     (N65)? 1'b0 : 
                     (N66)? 1'b0 : 
                     (N67)? 1'b0 : 
                     (N68)? 1'b0 : 
                     (N69)? 1'b0 : 
                     (N70)? 1'b0 : 
                     (N71)? 1'b0 : 
                     (N72)? 1'b0 : 
                     (N73)? yumi_int_o_9__1_ : 1'b0;
  assign yumi_o[0] = (N64)? 1'b0 : 
                     (N65)? 1'b0 : 
                     (N66)? 1'b0 : 
                     (N67)? 1'b0 : 
                     (N68)? 1'b0 : 
                     (N69)? 1'b0 : 
                     (N70)? 1'b0 : 
                     (N71)? 1'b0 : 
                     (N72)? 1'b0 : 
                     (N73)? yumi_int_o_9__0_ : 1'b0;
  assign _2_net__4_ = (N74)? 1'b0 : 
                      (N75)? 1'b0 : 
                      (N76)? 1'b0 : 
                      (N77)? 1'b0 : 
                      (N78)? 1'b0 : 
                      (N79)? 1'b0 : 
                      (N80)? 1'b0 : 
                      (N81)? 1'b0 : 
                      (N82)? 1'b0 : 
                      (N83)? valid_head_9__4_ : 1'b0;
  assign N74 = N112;
  assign N75 = N114;
  assign N76 = N116;
  assign N77 = N117;
  assign N78 = N118;
  assign N79 = N119;
  assign N80 = N120;
  assign N81 = N121;
  assign N82 = N113;
  assign N83 = N115;
  assign _2_net__3_ = (N74)? 1'b0 : 
                      (N75)? 1'b0 : 
                      (N76)? 1'b0 : 
                      (N77)? 1'b0 : 
                      (N78)? 1'b0 : 
                      (N79)? 1'b0 : 
                      (N80)? 1'b0 : 
                      (N81)? 1'b0 : 
                      (N82)? 1'b0 : 
                      (N83)? valid_head_9__3_ : 1'b0;
  assign _2_net__2_ = (N74)? 1'b0 : 
                      (N75)? 1'b0 : 
                      (N76)? 1'b0 : 
                      (N77)? 1'b0 : 
                      (N78)? 1'b0 : 
                      (N79)? 1'b0 : 
                      (N80)? 1'b0 : 
                      (N81)? 1'b0 : 
                      (N82)? 1'b0 : 
                      (N83)? valid_head_9__2_ : 1'b0;
  assign _2_net__1_ = (N74)? 1'b0 : 
                      (N75)? 1'b0 : 
                      (N76)? 1'b0 : 
                      (N77)? 1'b0 : 
                      (N78)? 1'b0 : 
                      (N79)? 1'b0 : 
                      (N80)? 1'b0 : 
                      (N81)? 1'b0 : 
                      (N82)? 1'b0 : 
                      (N83)? valid_head_9__1_ : 1'b0;
  assign _2_net__0_ = (N74)? 1'b0 : 
                      (N75)? 1'b0 : 
                      (N76)? 1'b0 : 
                      (N77)? 1'b0 : 
                      (N78)? 1'b0 : 
                      (N79)? 1'b0 : 
                      (N80)? 1'b0 : 
                      (N81)? 1'b0 : 
                      (N82)? 1'b0 : 
                      (N83)? valid_head_9__0_ : 1'b0;
  assign _4_net__159_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__159_ : 1'b0;
  assign N84 = N122;
  assign N85 = N124;
  assign N86 = N126;
  assign N87 = N127;
  assign N88 = N128;
  assign N89 = N129;
  assign N90 = N130;
  assign N91 = N131;
  assign N92 = N123;
  assign N93 = N125;
  assign _4_net__158_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__158_ : 1'b0;
  assign _4_net__157_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__157_ : 1'b0;
  assign _4_net__156_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__156_ : 1'b0;
  assign _4_net__155_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__155_ : 1'b0;
  assign _4_net__154_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__154_ : 1'b0;
  assign _4_net__153_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__153_ : 1'b0;
  assign _4_net__152_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__152_ : 1'b0;
  assign _4_net__151_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__151_ : 1'b0;
  assign _4_net__150_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__150_ : 1'b0;
  assign _4_net__149_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__149_ : 1'b0;
  assign _4_net__148_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__148_ : 1'b0;
  assign _4_net__147_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__147_ : 1'b0;
  assign _4_net__146_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__146_ : 1'b0;
  assign _4_net__145_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__145_ : 1'b0;
  assign _4_net__144_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__144_ : 1'b0;
  assign _4_net__143_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__143_ : 1'b0;
  assign _4_net__142_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__142_ : 1'b0;
  assign _4_net__141_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__141_ : 1'b0;
  assign _4_net__140_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__140_ : 1'b0;
  assign _4_net__139_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__139_ : 1'b0;
  assign _4_net__138_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__138_ : 1'b0;
  assign _4_net__137_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__137_ : 1'b0;
  assign _4_net__136_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__136_ : 1'b0;
  assign _4_net__135_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__135_ : 1'b0;
  assign _4_net__134_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__134_ : 1'b0;
  assign _4_net__133_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__133_ : 1'b0;
  assign _4_net__132_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__132_ : 1'b0;
  assign _4_net__131_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__131_ : 1'b0;
  assign _4_net__130_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__130_ : 1'b0;
  assign _4_net__129_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__129_ : 1'b0;
  assign _4_net__128_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__128_ : 1'b0;
  assign _4_net__127_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__127_ : 1'b0;
  assign _4_net__126_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__126_ : 1'b0;
  assign _4_net__125_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__125_ : 1'b0;
  assign _4_net__124_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__124_ : 1'b0;
  assign _4_net__123_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__123_ : 1'b0;
  assign _4_net__122_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__122_ : 1'b0;
  assign _4_net__121_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__121_ : 1'b0;
  assign _4_net__120_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__120_ : 1'b0;
  assign _4_net__119_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__119_ : 1'b0;
  assign _4_net__118_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__118_ : 1'b0;
  assign _4_net__117_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__117_ : 1'b0;
  assign _4_net__116_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__116_ : 1'b0;
  assign _4_net__115_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__115_ : 1'b0;
  assign _4_net__114_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__114_ : 1'b0;
  assign _4_net__113_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__113_ : 1'b0;
  assign _4_net__112_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__112_ : 1'b0;
  assign _4_net__111_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__111_ : 1'b0;
  assign _4_net__110_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__110_ : 1'b0;
  assign _4_net__109_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__109_ : 1'b0;
  assign _4_net__108_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__108_ : 1'b0;
  assign _4_net__107_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__107_ : 1'b0;
  assign _4_net__106_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__106_ : 1'b0;
  assign _4_net__105_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__105_ : 1'b0;
  assign _4_net__104_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__104_ : 1'b0;
  assign _4_net__103_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__103_ : 1'b0;
  assign _4_net__102_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__102_ : 1'b0;
  assign _4_net__101_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__101_ : 1'b0;
  assign _4_net__100_ = (N84)? 1'b0 : 
                        (N85)? 1'b0 : 
                        (N86)? 1'b0 : 
                        (N87)? 1'b0 : 
                        (N88)? 1'b0 : 
                        (N89)? 1'b0 : 
                        (N90)? 1'b0 : 
                        (N91)? 1'b0 : 
                        (N92)? 1'b0 : 
                        (N93)? data_head_9__100_ : 1'b0;
  assign _4_net__99_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__99_ : 1'b0;
  assign _4_net__98_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__98_ : 1'b0;
  assign _4_net__97_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__97_ : 1'b0;
  assign _4_net__96_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__96_ : 1'b0;
  assign _4_net__95_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__95_ : 1'b0;
  assign _4_net__94_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__94_ : 1'b0;
  assign _4_net__93_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__93_ : 1'b0;
  assign _4_net__92_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__92_ : 1'b0;
  assign _4_net__91_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__91_ : 1'b0;
  assign _4_net__90_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__90_ : 1'b0;
  assign _4_net__89_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__89_ : 1'b0;
  assign _4_net__88_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__88_ : 1'b0;
  assign _4_net__87_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__87_ : 1'b0;
  assign _4_net__86_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__86_ : 1'b0;
  assign _4_net__85_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__85_ : 1'b0;
  assign _4_net__84_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__84_ : 1'b0;
  assign _4_net__83_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__83_ : 1'b0;
  assign _4_net__82_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__82_ : 1'b0;
  assign _4_net__81_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__81_ : 1'b0;
  assign _4_net__80_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__80_ : 1'b0;
  assign _4_net__79_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__79_ : 1'b0;
  assign _4_net__78_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__78_ : 1'b0;
  assign _4_net__77_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__77_ : 1'b0;
  assign _4_net__76_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__76_ : 1'b0;
  assign _4_net__75_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__75_ : 1'b0;
  assign _4_net__74_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__74_ : 1'b0;
  assign _4_net__73_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__73_ : 1'b0;
  assign _4_net__72_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__72_ : 1'b0;
  assign _4_net__71_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__71_ : 1'b0;
  assign _4_net__70_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__70_ : 1'b0;
  assign _4_net__69_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__69_ : 1'b0;
  assign _4_net__68_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__68_ : 1'b0;
  assign _4_net__67_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__67_ : 1'b0;
  assign _4_net__66_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__66_ : 1'b0;
  assign _4_net__65_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__65_ : 1'b0;
  assign _4_net__64_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__64_ : 1'b0;
  assign _4_net__63_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__63_ : 1'b0;
  assign _4_net__62_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__62_ : 1'b0;
  assign _4_net__61_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__61_ : 1'b0;
  assign _4_net__60_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__60_ : 1'b0;
  assign _4_net__59_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__59_ : 1'b0;
  assign _4_net__58_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__58_ : 1'b0;
  assign _4_net__57_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__57_ : 1'b0;
  assign _4_net__56_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__56_ : 1'b0;
  assign _4_net__55_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__55_ : 1'b0;
  assign _4_net__54_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__54_ : 1'b0;
  assign _4_net__53_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__53_ : 1'b0;
  assign _4_net__52_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__52_ : 1'b0;
  assign _4_net__51_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__51_ : 1'b0;
  assign _4_net__50_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__50_ : 1'b0;
  assign _4_net__49_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__49_ : 1'b0;
  assign _4_net__48_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__48_ : 1'b0;
  assign _4_net__47_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__47_ : 1'b0;
  assign _4_net__46_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__46_ : 1'b0;
  assign _4_net__45_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__45_ : 1'b0;
  assign _4_net__44_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__44_ : 1'b0;
  assign _4_net__43_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__43_ : 1'b0;
  assign _4_net__42_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__42_ : 1'b0;
  assign _4_net__41_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__41_ : 1'b0;
  assign _4_net__40_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__40_ : 1'b0;
  assign _4_net__39_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__39_ : 1'b0;
  assign _4_net__38_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__38_ : 1'b0;
  assign _4_net__37_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__37_ : 1'b0;
  assign _4_net__36_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__36_ : 1'b0;
  assign _4_net__35_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__35_ : 1'b0;
  assign _4_net__34_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__34_ : 1'b0;
  assign _4_net__33_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__33_ : 1'b0;
  assign _4_net__32_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__32_ : 1'b0;
  assign _4_net__31_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__31_ : 1'b0;
  assign _4_net__30_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__30_ : 1'b0;
  assign _4_net__29_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__29_ : 1'b0;
  assign _4_net__28_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__28_ : 1'b0;
  assign _4_net__27_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__27_ : 1'b0;
  assign _4_net__26_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__26_ : 1'b0;
  assign _4_net__25_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__25_ : 1'b0;
  assign _4_net__24_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__24_ : 1'b0;
  assign _4_net__23_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__23_ : 1'b0;
  assign _4_net__22_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__22_ : 1'b0;
  assign _4_net__21_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__21_ : 1'b0;
  assign _4_net__20_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__20_ : 1'b0;
  assign _4_net__19_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__19_ : 1'b0;
  assign _4_net__18_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__18_ : 1'b0;
  assign _4_net__17_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__17_ : 1'b0;
  assign _4_net__16_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__16_ : 1'b0;
  assign _4_net__15_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__15_ : 1'b0;
  assign _4_net__14_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__14_ : 1'b0;
  assign _4_net__13_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__13_ : 1'b0;
  assign _4_net__12_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__12_ : 1'b0;
  assign _4_net__11_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__11_ : 1'b0;
  assign _4_net__10_ = (N84)? 1'b0 : 
                       (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? data_head_9__10_ : 1'b0;
  assign _4_net__9_ = (N84)? 1'b0 : 
                      (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? data_head_9__9_ : 1'b0;
  assign _4_net__8_ = (N84)? 1'b0 : 
                      (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? data_head_9__8_ : 1'b0;
  assign _4_net__7_ = (N84)? 1'b0 : 
                      (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? data_head_9__7_ : 1'b0;
  assign _4_net__6_ = (N84)? 1'b0 : 
                      (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? data_head_9__6_ : 1'b0;
  assign _4_net__5_ = (N84)? 1'b0 : 
                      (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? data_head_9__5_ : 1'b0;
  assign _4_net__4_ = (N84)? 1'b0 : 
                      (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? data_head_9__4_ : 1'b0;
  assign _4_net__3_ = (N84)? 1'b0 : 
                      (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? data_head_9__3_ : 1'b0;
  assign _4_net__2_ = (N84)? 1'b0 : 
                      (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? data_head_9__2_ : 1'b0;
  assign _4_net__1_ = (N84)? 1'b0 : 
                      (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? data_head_9__1_ : 1'b0;
  assign _4_net__0_ = (N84)? 1'b0 : 
                      (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? data_head_9__0_ : 1'b0;
  assign _0_net_ = reset | N136;
  assign _5_net_ = reset | N139;

endmodule



module bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  wire [63:0] mem;
  reg mem_63_sv2v_reg,mem_62_sv2v_reg,mem_61_sv2v_reg,mem_60_sv2v_reg,mem_59_sv2v_reg,
  mem_58_sv2v_reg,mem_57_sv2v_reg,mem_56_sv2v_reg,mem_55_sv2v_reg,mem_54_sv2v_reg,
  mem_53_sv2v_reg,mem_52_sv2v_reg,mem_51_sv2v_reg,mem_50_sv2v_reg,mem_49_sv2v_reg,
  mem_48_sv2v_reg,mem_47_sv2v_reg,mem_46_sv2v_reg,mem_45_sv2v_reg,mem_44_sv2v_reg,
  mem_43_sv2v_reg,mem_42_sv2v_reg,mem_41_sv2v_reg,mem_40_sv2v_reg,mem_39_sv2v_reg,
  mem_38_sv2v_reg,mem_37_sv2v_reg,mem_36_sv2v_reg,mem_35_sv2v_reg,mem_34_sv2v_reg,
  mem_33_sv2v_reg,mem_32_sv2v_reg,mem_31_sv2v_reg,mem_30_sv2v_reg,mem_29_sv2v_reg,
  mem_28_sv2v_reg,mem_27_sv2v_reg,mem_26_sv2v_reg,mem_25_sv2v_reg,mem_24_sv2v_reg,
  mem_23_sv2v_reg,mem_22_sv2v_reg,mem_21_sv2v_reg,mem_20_sv2v_reg,mem_19_sv2v_reg,
  mem_18_sv2v_reg,mem_17_sv2v_reg,mem_16_sv2v_reg,mem_15_sv2v_reg,mem_14_sv2v_reg,
  mem_13_sv2v_reg,mem_12_sv2v_reg,mem_11_sv2v_reg,mem_10_sv2v_reg,mem_9_sv2v_reg,
  mem_8_sv2v_reg,mem_7_sv2v_reg,mem_6_sv2v_reg,mem_5_sv2v_reg,mem_4_sv2v_reg,
  mem_3_sv2v_reg,mem_2_sv2v_reg,mem_1_sv2v_reg,mem_0_sv2v_reg;
  assign mem[63] = mem_63_sv2v_reg;
  assign mem[62] = mem_62_sv2v_reg;
  assign mem[61] = mem_61_sv2v_reg;
  assign mem[60] = mem_60_sv2v_reg;
  assign mem[59] = mem_59_sv2v_reg;
  assign mem[58] = mem_58_sv2v_reg;
  assign mem[57] = mem_57_sv2v_reg;
  assign mem[56] = mem_56_sv2v_reg;
  assign mem[55] = mem_55_sv2v_reg;
  assign mem[54] = mem_54_sv2v_reg;
  assign mem[53] = mem_53_sv2v_reg;
  assign mem[52] = mem_52_sv2v_reg;
  assign mem[51] = mem_51_sv2v_reg;
  assign mem[50] = mem_50_sv2v_reg;
  assign mem[49] = mem_49_sv2v_reg;
  assign mem[48] = mem_48_sv2v_reg;
  assign mem[47] = mem_47_sv2v_reg;
  assign mem[46] = mem_46_sv2v_reg;
  assign mem[45] = mem_45_sv2v_reg;
  assign mem[44] = mem_44_sv2v_reg;
  assign mem[43] = mem_43_sv2v_reg;
  assign mem[42] = mem_42_sv2v_reg;
  assign mem[41] = mem_41_sv2v_reg;
  assign mem[40] = mem_40_sv2v_reg;
  assign mem[39] = mem_39_sv2v_reg;
  assign mem[38] = mem_38_sv2v_reg;
  assign mem[37] = mem_37_sv2v_reg;
  assign mem[36] = mem_36_sv2v_reg;
  assign mem[35] = mem_35_sv2v_reg;
  assign mem[34] = mem_34_sv2v_reg;
  assign mem[33] = mem_33_sv2v_reg;
  assign mem[32] = mem_32_sv2v_reg;
  assign mem[31] = mem_31_sv2v_reg;
  assign mem[30] = mem_30_sv2v_reg;
  assign mem[29] = mem_29_sv2v_reg;
  assign mem[28] = mem_28_sv2v_reg;
  assign mem[27] = mem_27_sv2v_reg;
  assign mem[26] = mem_26_sv2v_reg;
  assign mem[25] = mem_25_sv2v_reg;
  assign mem[24] = mem_24_sv2v_reg;
  assign mem[23] = mem_23_sv2v_reg;
  assign mem[22] = mem_22_sv2v_reg;
  assign mem[21] = mem_21_sv2v_reg;
  assign mem[20] = mem_20_sv2v_reg;
  assign mem[19] = mem_19_sv2v_reg;
  assign mem[18] = mem_18_sv2v_reg;
  assign mem[17] = mem_17_sv2v_reg;
  assign mem[16] = mem_16_sv2v_reg;
  assign mem[15] = mem_15_sv2v_reg;
  assign mem[14] = mem_14_sv2v_reg;
  assign mem[13] = mem_13_sv2v_reg;
  assign mem[12] = mem_12_sv2v_reg;
  assign mem[11] = mem_11_sv2v_reg;
  assign mem[10] = mem_10_sv2v_reg;
  assign mem[9] = mem_9_sv2v_reg;
  assign mem[8] = mem_8_sv2v_reg;
  assign mem[7] = mem_7_sv2v_reg;
  assign mem[6] = mem_6_sv2v_reg;
  assign mem[5] = mem_5_sv2v_reg;
  assign mem[4] = mem_4_sv2v_reg;
  assign mem[3] = mem_3_sv2v_reg;
  assign mem[2] = mem_2_sv2v_reg;
  assign mem[1] = mem_1_sv2v_reg;
  assign mem[0] = mem_0_sv2v_reg;
  assign r_data_o[31] = (N3)? mem[31] : 
                        (N0)? mem[63] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[30] = (N3)? mem[30] : 
                        (N0)? mem[62] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] : 
                        (N0)? mem[61] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] : 
                        (N0)? mem[60] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] : 
                        (N0)? mem[59] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] : 
                        (N0)? mem[58] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] : 
                        (N0)? mem[57] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] : 
                        (N0)? mem[56] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] : 
                        (N0)? mem[55] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] : 
                        (N0)? mem[54] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] : 
                        (N0)? mem[53] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] : 
                        (N0)? mem[52] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] : 
                        (N0)? mem[51] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] : 
                        (N0)? mem[50] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] : 
                        (N0)? mem[49] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] : 
                        (N0)? mem[48] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] : 
                        (N0)? mem[47] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] : 
                        (N0)? mem[46] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] : 
                        (N0)? mem[45] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] : 
                        (N0)? mem[44] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] : 
                        (N0)? mem[43] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] : 
                        (N0)? mem[42] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] : 
                       (N0)? mem[41] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] : 
                       (N0)? mem[40] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] : 
                       (N0)? mem[39] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] : 
                       (N0)? mem[38] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[37] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[36] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[35] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[34] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[33] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[32] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_63_sv2v_reg <= w_data_i[31];
      mem_62_sv2v_reg <= w_data_i[30];
      mem_61_sv2v_reg <= w_data_i[29];
      mem_60_sv2v_reg <= w_data_i[28];
      mem_59_sv2v_reg <= w_data_i[27];
      mem_58_sv2v_reg <= w_data_i[26];
      mem_57_sv2v_reg <= w_data_i[25];
      mem_56_sv2v_reg <= w_data_i[24];
      mem_55_sv2v_reg <= w_data_i[23];
      mem_54_sv2v_reg <= w_data_i[22];
      mem_53_sv2v_reg <= w_data_i[21];
      mem_52_sv2v_reg <= w_data_i[20];
      mem_51_sv2v_reg <= w_data_i[19];
      mem_50_sv2v_reg <= w_data_i[18];
      mem_49_sv2v_reg <= w_data_i[17];
      mem_48_sv2v_reg <= w_data_i[16];
      mem_47_sv2v_reg <= w_data_i[15];
      mem_46_sv2v_reg <= w_data_i[14];
      mem_45_sv2v_reg <= w_data_i[13];
      mem_44_sv2v_reg <= w_data_i[12];
      mem_43_sv2v_reg <= w_data_i[11];
      mem_42_sv2v_reg <= w_data_i[10];
      mem_41_sv2v_reg <= w_data_i[9];
      mem_40_sv2v_reg <= w_data_i[8];
      mem_39_sv2v_reg <= w_data_i[7];
      mem_38_sv2v_reg <= w_data_i[6];
      mem_37_sv2v_reg <= w_data_i[5];
      mem_36_sv2v_reg <= w_data_i[4];
      mem_35_sv2v_reg <= w_data_i[3];
      mem_34_sv2v_reg <= w_data_i[2];
      mem_33_sv2v_reg <= w_data_i[1];
      mem_32_sv2v_reg <= w_data_i[0];
    end 
    if(N7) begin
      mem_31_sv2v_reg <= w_data_i[31];
      mem_30_sv2v_reg <= w_data_i[30];
      mem_29_sv2v_reg <= w_data_i[29];
      mem_28_sv2v_reg <= w_data_i[28];
      mem_27_sv2v_reg <= w_data_i[27];
      mem_26_sv2v_reg <= w_data_i[26];
      mem_25_sv2v_reg <= w_data_i[25];
      mem_24_sv2v_reg <= w_data_i[24];
      mem_23_sv2v_reg <= w_data_i[23];
      mem_22_sv2v_reg <= w_data_i[22];
      mem_21_sv2v_reg <= w_data_i[21];
      mem_20_sv2v_reg <= w_data_i[20];
      mem_19_sv2v_reg <= w_data_i[19];
      mem_18_sv2v_reg <= w_data_i[18];
      mem_17_sv2v_reg <= w_data_i[17];
      mem_16_sv2v_reg <= w_data_i[16];
      mem_15_sv2v_reg <= w_data_i[15];
      mem_14_sv2v_reg <= w_data_i[14];
      mem_13_sv2v_reg <= w_data_i[13];
      mem_12_sv2v_reg <= w_data_i[12];
      mem_11_sv2v_reg <= w_data_i[11];
      mem_10_sv2v_reg <= w_data_i[10];
      mem_9_sv2v_reg <= w_data_i[9];
      mem_8_sv2v_reg <= w_data_i[8];
      mem_7_sv2v_reg <= w_data_i[7];
      mem_6_sv2v_reg <= w_data_i[6];
      mem_5_sv2v_reg <= w_data_i[5];
      mem_4_sv2v_reg <= w_data_i[4];
      mem_3_sv2v_reg <= w_data_i[3];
      mem_2_sv2v_reg <= w_data_i[2];
      mem_1_sv2v_reg <= w_data_i[1];
      mem_0_sv2v_reg <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;

  bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p32
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,enq_i,tail_r,_0_net_,head_r,empty_r,full_r,N0,N1,N2,N3,N4,N5,N6,N7,
  N8,N9,N10,N11,N12,N13,N14;
  reg full_r_sv2v_reg,tail_r_sv2v_reg,head_r_sv2v_reg,empty_r_sv2v_reg;
  assign full_r = full_r_sv2v_reg;
  assign tail_r = tail_r_sv2v_reg;
  assign head_r = head_r_sv2v_reg;
  assign empty_r = empty_r_sv2v_reg;

  bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign _0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N5;
  assign N5 = ~full_r;
  assign N1 = enq_i;
  assign N0 = ~tail_r;
  assign N2 = ~head_r;
  assign N3 = N7 | N9;
  assign N7 = empty_r & N6;
  assign N6 = ~enq_i;
  assign N9 = N8 & N6;
  assign N8 = N5 & yumi_i;
  assign N4 = N13 | N14;
  assign N13 = N11 & N12;
  assign N11 = N10 & enq_i;
  assign N10 = ~empty_r;
  assign N12 = ~yumi_i;
  assign N14 = full_r & N12;

  always @(posedge clk_i) begin
    if(reset_i) begin
      full_r_sv2v_reg <= 1'b0;
      empty_r_sv2v_reg <= 1'b1;
    end else if(1'b1) begin
      full_r_sv2v_reg <= N4;
      empty_r_sv2v_reg <= N3;
    end 
    if(reset_i) begin
      tail_r_sv2v_reg <= 1'b0;
    end else if(N1) begin
      tail_r_sv2v_reg <= N0;
    end 
    if(reset_i) begin
      head_r_sv2v_reg <= 1'b0;
    end else if(yumi_i) begin
      head_r_sv2v_reg <= N2;
    end 
  end


endmodule



module bsg_assembler_in
(
  clk,
  reset,
  calibration_done_i,
  valid_i,
  data_i,
  yumi_o,
  in_top_channel_i,
  out_top_channel_i,
  valid_o,
  data_o,
  yumi_i
);

  input [9:0] valid_i;
  input [319:0] data_i;
  output [9:0] yumi_o;
  input [3:0] in_top_channel_i;
  input [2:0] out_top_channel_i;
  output [159:0] data_o;
  input clk;
  input reset;
  input calibration_done_i;
  input yumi_i;
  output valid_o;
  wire [9:0] yumi_o;
  wire [159:0] data_o,fifo_data_vec;
  wire valid_o,_0_net__9_,_0_net__8_,_0_net__7_,_0_net__6_,_0_net__5_,_0_net__4_,
  _0_net__3_,_0_net__2_,_0_net__1_,_0_net__0_,N0,N1,N2,N3;
  wire [4:0] fifo_enq_vec,fifo_not_full_vec,fifo_valid_vec;

  bsg_round_robin_fifo_to_fifo_width_p32_num_in_p10_num_out_p5_in_channel_count_mask_p512
  rr_fifo_to_fifo
  (
    .clk(clk),
    .reset(reset),
    .valid_i({ _0_net__9_, _0_net__8_, _0_net__7_, _0_net__6_, _0_net__5_, _0_net__4_, _0_net__3_, _0_net__2_, _0_net__1_, _0_net__0_ }),
    .data_i(data_i),
    .yumi_o(yumi_o),
    .in_top_channel_i(in_top_channel_i),
    .out_top_channel_i(out_top_channel_i),
    .valid_o(fifo_enq_vec),
    .data_o(fifo_data_vec),
    .ready_i(fifo_not_full_vec)
  );


  bsg_two_fifo_width_p32
  \fifos_0_.ring_packet_fifo 
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[0]),
    .data_i(fifo_data_vec[31:0]),
    .v_i(fifo_enq_vec[0]),
    .v_o(fifo_valid_vec[0]),
    .data_o(data_o[31:0]),
    .yumi_i(yumi_i)
  );


  bsg_two_fifo_width_p32
  \fifos_1_.ring_packet_fifo 
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[1]),
    .data_i(fifo_data_vec[63:32]),
    .v_i(fifo_enq_vec[1]),
    .v_o(fifo_valid_vec[1]),
    .data_o(data_o[63:32]),
    .yumi_i(yumi_i)
  );


  bsg_two_fifo_width_p32
  \fifos_2_.ring_packet_fifo 
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[2]),
    .data_i(fifo_data_vec[95:64]),
    .v_i(fifo_enq_vec[2]),
    .v_o(fifo_valid_vec[2]),
    .data_o(data_o[95:64]),
    .yumi_i(yumi_i)
  );


  bsg_two_fifo_width_p32
  \fifos_3_.ring_packet_fifo 
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[3]),
    .data_i(fifo_data_vec[127:96]),
    .v_i(fifo_enq_vec[3]),
    .v_o(fifo_valid_vec[3]),
    .data_o(data_o[127:96]),
    .yumi_i(yumi_i)
  );


  bsg_two_fifo_width_p32
  \fifos_4_.ring_packet_fifo 
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[4]),
    .data_i(fifo_data_vec[159:128]),
    .v_i(fifo_enq_vec[4]),
    .v_o(fifo_valid_vec[4]),
    .data_o(data_o[159:128]),
    .yumi_i(yumi_i)
  );

  assign _0_net__9_ = valid_i[9] & calibration_done_i;
  assign _0_net__8_ = valid_i[8] & calibration_done_i;
  assign _0_net__7_ = valid_i[7] & calibration_done_i;
  assign _0_net__6_ = valid_i[6] & calibration_done_i;
  assign _0_net__5_ = valid_i[5] & calibration_done_i;
  assign _0_net__4_ = valid_i[4] & calibration_done_i;
  assign _0_net__3_ = valid_i[3] & calibration_done_i;
  assign _0_net__2_ = valid_i[2] & calibration_done_i;
  assign _0_net__1_ = valid_i[1] & calibration_done_i;
  assign _0_net__0_ = valid_i[0] & calibration_done_i;
  assign valid_o = N3 & calibration_done_i;
  assign N3 = N2 & fifo_valid_vec[0];
  assign N2 = N1 & fifo_valid_vec[1];
  assign N1 = N0 & fifo_valid_vec[2];
  assign N0 = fifo_valid_vec[4] & fifo_valid_vec[3];

endmodule

