

module top
(
  clk,
  reset,
  calibration_done_i,
  valid_i,
  data_i,
  ready_o,
  in_top_channel_i,
  out_top_channel_i,
  valid_o,
  data_o,
  ready_i
);

  input [639:0] data_i;
  input [3:0] in_top_channel_i;
  input [3:0] out_top_channel_i;
  output [9:0] valid_o;
  output [639:0] data_o;
  input [9:0] ready_i;
  input clk;
  input reset;
  input calibration_done_i;
  input valid_i;
  output ready_o;

  bsg_assembler_out
  wrapper
  (
    .data_i(data_i),
    .in_top_channel_i(in_top_channel_i),
    .out_top_channel_i(out_top_channel_i),
    .valid_o(valid_o),
    .data_o(data_o),
    .ready_i(ready_i),
    .clk(clk),
    .reset(reset),
    .calibration_done_i(calibration_done_i),
    .valid_i(valid_i),
    .ready_o(ready_o)
  );


endmodule



module bsg_mem_1r1w_synth_width_p64_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [63:0] w_data_i;
  input [0:0] r_addr_i;
  output [63:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [63:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  reg [127:0] mem;
  assign r_data_o[63] = (N3)? mem[63] : 
                        (N0)? mem[127] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[62] = (N3)? mem[62] : 
                        (N0)? mem[126] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] : 
                        (N0)? mem[125] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] : 
                        (N0)? mem[124] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] : 
                        (N0)? mem[123] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] : 
                        (N0)? mem[122] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] : 
                        (N0)? mem[121] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] : 
                        (N0)? mem[120] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] : 
                        (N0)? mem[119] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] : 
                        (N0)? mem[118] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] : 
                        (N0)? mem[117] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] : 
                        (N0)? mem[116] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] : 
                        (N0)? mem[115] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] : 
                        (N0)? mem[114] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] : 
                        (N0)? mem[113] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] : 
                        (N0)? mem[112] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] : 
                        (N0)? mem[111] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] : 
                        (N0)? mem[110] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] : 
                        (N0)? mem[109] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] : 
                        (N0)? mem[108] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] : 
                        (N0)? mem[107] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] : 
                        (N0)? mem[106] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] : 
                        (N0)? mem[105] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] : 
                        (N0)? mem[104] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] : 
                        (N0)? mem[103] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] : 
                        (N0)? mem[102] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] : 
                        (N0)? mem[101] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] : 
                        (N0)? mem[100] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] : 
                        (N0)? mem[99] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] : 
                        (N0)? mem[98] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] : 
                        (N0)? mem[97] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] : 
                        (N0)? mem[96] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] : 
                        (N0)? mem[95] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] : 
                        (N0)? mem[94] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] : 
                        (N0)? mem[93] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] : 
                        (N0)? mem[92] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] : 
                        (N0)? mem[91] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] : 
                        (N0)? mem[90] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] : 
                        (N0)? mem[89] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] : 
                        (N0)? mem[88] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] : 
                        (N0)? mem[87] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] : 
                        (N0)? mem[86] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] : 
                        (N0)? mem[85] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] : 
                        (N0)? mem[84] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] : 
                        (N0)? mem[83] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] : 
                        (N0)? mem[82] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] : 
                        (N0)? mem[81] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] : 
                        (N0)? mem[80] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] : 
                        (N0)? mem[79] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] : 
                        (N0)? mem[78] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] : 
                        (N0)? mem[77] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] : 
                        (N0)? mem[76] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] : 
                        (N0)? mem[75] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] : 
                        (N0)? mem[74] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] : 
                       (N0)? mem[73] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] : 
                       (N0)? mem[72] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] : 
                       (N0)? mem[71] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] : 
                       (N0)? mem[70] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[69] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[68] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[67] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[66] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[65] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[64] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      { mem[127:64] } <= { w_data_i[63:0] };
    end 
    if(N7) begin
      { mem[63:0] } <= { w_data_i[63:0] };
    end 
  end


endmodule



module bsg_mem_1r1w_width_p64_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [63:0] w_data_i;
  input [0:0] r_addr_i;
  output [63:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [63:0] r_data_o;

  bsg_mem_1r1w_synth_width_p64_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p64_ready_THEN_valid_p1
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [63:0] data_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [63:0] data_o;
  wire ready_o,v_o,N0,N1,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,
  N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p64_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(v_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 : 
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 : 
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 : 
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 : 
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 : 
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 : 
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = v_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N16 | N19;
  assign N16 = empty_r & N15;
  assign N15 = ~v_i;
  assign N19 = N18 & N15;
  assign N18 = N17 & yumi_i;
  assign N17 = ~full_r;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & v_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end 
    if(N9) begin
      tail_r <= N10;
    end 
    if(N11) begin
      head_r <= N12;
    end 
  end


endmodule



module bsg_make_2D_array_width_p64_items_p10
(
  i,
  o
);

  input [639:0] i;
  output [639:0] o;
  wire [639:0] o;
  assign o[639] = i[639];
  assign o[638] = i[638];
  assign o[637] = i[637];
  assign o[636] = i[636];
  assign o[635] = i[635];
  assign o[634] = i[634];
  assign o[633] = i[633];
  assign o[632] = i[632];
  assign o[631] = i[631];
  assign o[630] = i[630];
  assign o[629] = i[629];
  assign o[628] = i[628];
  assign o[627] = i[627];
  assign o[626] = i[626];
  assign o[625] = i[625];
  assign o[624] = i[624];
  assign o[623] = i[623];
  assign o[622] = i[622];
  assign o[621] = i[621];
  assign o[620] = i[620];
  assign o[619] = i[619];
  assign o[618] = i[618];
  assign o[617] = i[617];
  assign o[616] = i[616];
  assign o[615] = i[615];
  assign o[614] = i[614];
  assign o[613] = i[613];
  assign o[612] = i[612];
  assign o[611] = i[611];
  assign o[610] = i[610];
  assign o[609] = i[609];
  assign o[608] = i[608];
  assign o[607] = i[607];
  assign o[606] = i[606];
  assign o[605] = i[605];
  assign o[604] = i[604];
  assign o[603] = i[603];
  assign o[602] = i[602];
  assign o[601] = i[601];
  assign o[600] = i[600];
  assign o[599] = i[599];
  assign o[598] = i[598];
  assign o[597] = i[597];
  assign o[596] = i[596];
  assign o[595] = i[595];
  assign o[594] = i[594];
  assign o[593] = i[593];
  assign o[592] = i[592];
  assign o[591] = i[591];
  assign o[590] = i[590];
  assign o[589] = i[589];
  assign o[588] = i[588];
  assign o[587] = i[587];
  assign o[586] = i[586];
  assign o[585] = i[585];
  assign o[584] = i[584];
  assign o[583] = i[583];
  assign o[582] = i[582];
  assign o[581] = i[581];
  assign o[580] = i[580];
  assign o[579] = i[579];
  assign o[578] = i[578];
  assign o[577] = i[577];
  assign o[576] = i[576];
  assign o[575] = i[575];
  assign o[574] = i[574];
  assign o[573] = i[573];
  assign o[572] = i[572];
  assign o[571] = i[571];
  assign o[570] = i[570];
  assign o[569] = i[569];
  assign o[568] = i[568];
  assign o[567] = i[567];
  assign o[566] = i[566];
  assign o[565] = i[565];
  assign o[564] = i[564];
  assign o[563] = i[563];
  assign o[562] = i[562];
  assign o[561] = i[561];
  assign o[560] = i[560];
  assign o[559] = i[559];
  assign o[558] = i[558];
  assign o[557] = i[557];
  assign o[556] = i[556];
  assign o[555] = i[555];
  assign o[554] = i[554];
  assign o[553] = i[553];
  assign o[552] = i[552];
  assign o[551] = i[551];
  assign o[550] = i[550];
  assign o[549] = i[549];
  assign o[548] = i[548];
  assign o[547] = i[547];
  assign o[546] = i[546];
  assign o[545] = i[545];
  assign o[544] = i[544];
  assign o[543] = i[543];
  assign o[542] = i[542];
  assign o[541] = i[541];
  assign o[540] = i[540];
  assign o[539] = i[539];
  assign o[538] = i[538];
  assign o[537] = i[537];
  assign o[536] = i[536];
  assign o[535] = i[535];
  assign o[534] = i[534];
  assign o[533] = i[533];
  assign o[532] = i[532];
  assign o[531] = i[531];
  assign o[530] = i[530];
  assign o[529] = i[529];
  assign o[528] = i[528];
  assign o[527] = i[527];
  assign o[526] = i[526];
  assign o[525] = i[525];
  assign o[524] = i[524];
  assign o[523] = i[523];
  assign o[522] = i[522];
  assign o[521] = i[521];
  assign o[520] = i[520];
  assign o[519] = i[519];
  assign o[518] = i[518];
  assign o[517] = i[517];
  assign o[516] = i[516];
  assign o[515] = i[515];
  assign o[514] = i[514];
  assign o[513] = i[513];
  assign o[512] = i[512];
  assign o[511] = i[511];
  assign o[510] = i[510];
  assign o[509] = i[509];
  assign o[508] = i[508];
  assign o[507] = i[507];
  assign o[506] = i[506];
  assign o[505] = i[505];
  assign o[504] = i[504];
  assign o[503] = i[503];
  assign o[502] = i[502];
  assign o[501] = i[501];
  assign o[500] = i[500];
  assign o[499] = i[499];
  assign o[498] = i[498];
  assign o[497] = i[497];
  assign o[496] = i[496];
  assign o[495] = i[495];
  assign o[494] = i[494];
  assign o[493] = i[493];
  assign o[492] = i[492];
  assign o[491] = i[491];
  assign o[490] = i[490];
  assign o[489] = i[489];
  assign o[488] = i[488];
  assign o[487] = i[487];
  assign o[486] = i[486];
  assign o[485] = i[485];
  assign o[484] = i[484];
  assign o[483] = i[483];
  assign o[482] = i[482];
  assign o[481] = i[481];
  assign o[480] = i[480];
  assign o[479] = i[479];
  assign o[478] = i[478];
  assign o[477] = i[477];
  assign o[476] = i[476];
  assign o[475] = i[475];
  assign o[474] = i[474];
  assign o[473] = i[473];
  assign o[472] = i[472];
  assign o[471] = i[471];
  assign o[470] = i[470];
  assign o[469] = i[469];
  assign o[468] = i[468];
  assign o[467] = i[467];
  assign o[466] = i[466];
  assign o[465] = i[465];
  assign o[464] = i[464];
  assign o[463] = i[463];
  assign o[462] = i[462];
  assign o[461] = i[461];
  assign o[460] = i[460];
  assign o[459] = i[459];
  assign o[458] = i[458];
  assign o[457] = i[457];
  assign o[456] = i[456];
  assign o[455] = i[455];
  assign o[454] = i[454];
  assign o[453] = i[453];
  assign o[452] = i[452];
  assign o[451] = i[451];
  assign o[450] = i[450];
  assign o[449] = i[449];
  assign o[448] = i[448];
  assign o[447] = i[447];
  assign o[446] = i[446];
  assign o[445] = i[445];
  assign o[444] = i[444];
  assign o[443] = i[443];
  assign o[442] = i[442];
  assign o[441] = i[441];
  assign o[440] = i[440];
  assign o[439] = i[439];
  assign o[438] = i[438];
  assign o[437] = i[437];
  assign o[436] = i[436];
  assign o[435] = i[435];
  assign o[434] = i[434];
  assign o[433] = i[433];
  assign o[432] = i[432];
  assign o[431] = i[431];
  assign o[430] = i[430];
  assign o[429] = i[429];
  assign o[428] = i[428];
  assign o[427] = i[427];
  assign o[426] = i[426];
  assign o[425] = i[425];
  assign o[424] = i[424];
  assign o[423] = i[423];
  assign o[422] = i[422];
  assign o[421] = i[421];
  assign o[420] = i[420];
  assign o[419] = i[419];
  assign o[418] = i[418];
  assign o[417] = i[417];
  assign o[416] = i[416];
  assign o[415] = i[415];
  assign o[414] = i[414];
  assign o[413] = i[413];
  assign o[412] = i[412];
  assign o[411] = i[411];
  assign o[410] = i[410];
  assign o[409] = i[409];
  assign o[408] = i[408];
  assign o[407] = i[407];
  assign o[406] = i[406];
  assign o[405] = i[405];
  assign o[404] = i[404];
  assign o[403] = i[403];
  assign o[402] = i[402];
  assign o[401] = i[401];
  assign o[400] = i[400];
  assign o[399] = i[399];
  assign o[398] = i[398];
  assign o[397] = i[397];
  assign o[396] = i[396];
  assign o[395] = i[395];
  assign o[394] = i[394];
  assign o[393] = i[393];
  assign o[392] = i[392];
  assign o[391] = i[391];
  assign o[390] = i[390];
  assign o[389] = i[389];
  assign o[388] = i[388];
  assign o[387] = i[387];
  assign o[386] = i[386];
  assign o[385] = i[385];
  assign o[384] = i[384];
  assign o[383] = i[383];
  assign o[382] = i[382];
  assign o[381] = i[381];
  assign o[380] = i[380];
  assign o[379] = i[379];
  assign o[378] = i[378];
  assign o[377] = i[377];
  assign o[376] = i[376];
  assign o[375] = i[375];
  assign o[374] = i[374];
  assign o[373] = i[373];
  assign o[372] = i[372];
  assign o[371] = i[371];
  assign o[370] = i[370];
  assign o[369] = i[369];
  assign o[368] = i[368];
  assign o[367] = i[367];
  assign o[366] = i[366];
  assign o[365] = i[365];
  assign o[364] = i[364];
  assign o[363] = i[363];
  assign o[362] = i[362];
  assign o[361] = i[361];
  assign o[360] = i[360];
  assign o[359] = i[359];
  assign o[358] = i[358];
  assign o[357] = i[357];
  assign o[356] = i[356];
  assign o[355] = i[355];
  assign o[354] = i[354];
  assign o[353] = i[353];
  assign o[352] = i[352];
  assign o[351] = i[351];
  assign o[350] = i[350];
  assign o[349] = i[349];
  assign o[348] = i[348];
  assign o[347] = i[347];
  assign o[346] = i[346];
  assign o[345] = i[345];
  assign o[344] = i[344];
  assign o[343] = i[343];
  assign o[342] = i[342];
  assign o[341] = i[341];
  assign o[340] = i[340];
  assign o[339] = i[339];
  assign o[338] = i[338];
  assign o[337] = i[337];
  assign o[336] = i[336];
  assign o[335] = i[335];
  assign o[334] = i[334];
  assign o[333] = i[333];
  assign o[332] = i[332];
  assign o[331] = i[331];
  assign o[330] = i[330];
  assign o[329] = i[329];
  assign o[328] = i[328];
  assign o[327] = i[327];
  assign o[326] = i[326];
  assign o[325] = i[325];
  assign o[324] = i[324];
  assign o[323] = i[323];
  assign o[322] = i[322];
  assign o[321] = i[321];
  assign o[320] = i[320];
  assign o[319] = i[319];
  assign o[318] = i[318];
  assign o[317] = i[317];
  assign o[316] = i[316];
  assign o[315] = i[315];
  assign o[314] = i[314];
  assign o[313] = i[313];
  assign o[312] = i[312];
  assign o[311] = i[311];
  assign o[310] = i[310];
  assign o[309] = i[309];
  assign o[308] = i[308];
  assign o[307] = i[307];
  assign o[306] = i[306];
  assign o[305] = i[305];
  assign o[304] = i[304];
  assign o[303] = i[303];
  assign o[302] = i[302];
  assign o[301] = i[301];
  assign o[300] = i[300];
  assign o[299] = i[299];
  assign o[298] = i[298];
  assign o[297] = i[297];
  assign o[296] = i[296];
  assign o[295] = i[295];
  assign o[294] = i[294];
  assign o[293] = i[293];
  assign o[292] = i[292];
  assign o[291] = i[291];
  assign o[290] = i[290];
  assign o[289] = i[289];
  assign o[288] = i[288];
  assign o[287] = i[287];
  assign o[286] = i[286];
  assign o[285] = i[285];
  assign o[284] = i[284];
  assign o[283] = i[283];
  assign o[282] = i[282];
  assign o[281] = i[281];
  assign o[280] = i[280];
  assign o[279] = i[279];
  assign o[278] = i[278];
  assign o[277] = i[277];
  assign o[276] = i[276];
  assign o[275] = i[275];
  assign o[274] = i[274];
  assign o[273] = i[273];
  assign o[272] = i[272];
  assign o[271] = i[271];
  assign o[270] = i[270];
  assign o[269] = i[269];
  assign o[268] = i[268];
  assign o[267] = i[267];
  assign o[266] = i[266];
  assign o[265] = i[265];
  assign o[264] = i[264];
  assign o[263] = i[263];
  assign o[262] = i[262];
  assign o[261] = i[261];
  assign o[260] = i[260];
  assign o[259] = i[259];
  assign o[258] = i[258];
  assign o[257] = i[257];
  assign o[256] = i[256];
  assign o[255] = i[255];
  assign o[254] = i[254];
  assign o[253] = i[253];
  assign o[252] = i[252];
  assign o[251] = i[251];
  assign o[250] = i[250];
  assign o[249] = i[249];
  assign o[248] = i[248];
  assign o[247] = i[247];
  assign o[246] = i[246];
  assign o[245] = i[245];
  assign o[244] = i[244];
  assign o[243] = i[243];
  assign o[242] = i[242];
  assign o[241] = i[241];
  assign o[240] = i[240];
  assign o[239] = i[239];
  assign o[238] = i[238];
  assign o[237] = i[237];
  assign o[236] = i[236];
  assign o[235] = i[235];
  assign o[234] = i[234];
  assign o[233] = i[233];
  assign o[232] = i[232];
  assign o[231] = i[231];
  assign o[230] = i[230];
  assign o[229] = i[229];
  assign o[228] = i[228];
  assign o[227] = i[227];
  assign o[226] = i[226];
  assign o[225] = i[225];
  assign o[224] = i[224];
  assign o[223] = i[223];
  assign o[222] = i[222];
  assign o[221] = i[221];
  assign o[220] = i[220];
  assign o[219] = i[219];
  assign o[218] = i[218];
  assign o[217] = i[217];
  assign o[216] = i[216];
  assign o[215] = i[215];
  assign o[214] = i[214];
  assign o[213] = i[213];
  assign o[212] = i[212];
  assign o[211] = i[211];
  assign o[210] = i[210];
  assign o[209] = i[209];
  assign o[208] = i[208];
  assign o[207] = i[207];
  assign o[206] = i[206];
  assign o[205] = i[205];
  assign o[204] = i[204];
  assign o[203] = i[203];
  assign o[202] = i[202];
  assign o[201] = i[201];
  assign o[200] = i[200];
  assign o[199] = i[199];
  assign o[198] = i[198];
  assign o[197] = i[197];
  assign o[196] = i[196];
  assign o[195] = i[195];
  assign o[194] = i[194];
  assign o[193] = i[193];
  assign o[192] = i[192];
  assign o[191] = i[191];
  assign o[190] = i[190];
  assign o[189] = i[189];
  assign o[188] = i[188];
  assign o[187] = i[187];
  assign o[186] = i[186];
  assign o[185] = i[185];
  assign o[184] = i[184];
  assign o[183] = i[183];
  assign o[182] = i[182];
  assign o[181] = i[181];
  assign o[180] = i[180];
  assign o[179] = i[179];
  assign o[178] = i[178];
  assign o[177] = i[177];
  assign o[176] = i[176];
  assign o[175] = i[175];
  assign o[174] = i[174];
  assign o[173] = i[173];
  assign o[172] = i[172];
  assign o[171] = i[171];
  assign o[170] = i[170];
  assign o[169] = i[169];
  assign o[168] = i[168];
  assign o[167] = i[167];
  assign o[166] = i[166];
  assign o[165] = i[165];
  assign o[164] = i[164];
  assign o[163] = i[163];
  assign o[162] = i[162];
  assign o[161] = i[161];
  assign o[160] = i[160];
  assign o[159] = i[159];
  assign o[158] = i[158];
  assign o[157] = i[157];
  assign o[156] = i[156];
  assign o[155] = i[155];
  assign o[154] = i[154];
  assign o[153] = i[153];
  assign o[152] = i[152];
  assign o[151] = i[151];
  assign o[150] = i[150];
  assign o[149] = i[149];
  assign o[148] = i[148];
  assign o[147] = i[147];
  assign o[146] = i[146];
  assign o[145] = i[145];
  assign o[144] = i[144];
  assign o[143] = i[143];
  assign o[142] = i[142];
  assign o[141] = i[141];
  assign o[140] = i[140];
  assign o[139] = i[139];
  assign o[138] = i[138];
  assign o[137] = i[137];
  assign o[136] = i[136];
  assign o[135] = i[135];
  assign o[134] = i[134];
  assign o[133] = i[133];
  assign o[132] = i[132];
  assign o[131] = i[131];
  assign o[130] = i[130];
  assign o[129] = i[129];
  assign o[128] = i[128];
  assign o[127] = i[127];
  assign o[126] = i[126];
  assign o[125] = i[125];
  assign o[124] = i[124];
  assign o[123] = i[123];
  assign o[122] = i[122];
  assign o[121] = i[121];
  assign o[120] = i[120];
  assign o[119] = i[119];
  assign o[118] = i[118];
  assign o[117] = i[117];
  assign o[116] = i[116];
  assign o[115] = i[115];
  assign o[114] = i[114];
  assign o[113] = i[113];
  assign o[112] = i[112];
  assign o[111] = i[111];
  assign o[110] = i[110];
  assign o[109] = i[109];
  assign o[108] = i[108];
  assign o[107] = i[107];
  assign o[106] = i[106];
  assign o[105] = i[105];
  assign o[104] = i[104];
  assign o[103] = i[103];
  assign o[102] = i[102];
  assign o[101] = i[101];
  assign o[100] = i[100];
  assign o[99] = i[99];
  assign o[98] = i[98];
  assign o[97] = i[97];
  assign o[96] = i[96];
  assign o[95] = i[95];
  assign o[94] = i[94];
  assign o[93] = i[93];
  assign o[92] = i[92];
  assign o[91] = i[91];
  assign o[90] = i[90];
  assign o[89] = i[89];
  assign o[88] = i[88];
  assign o[87] = i[87];
  assign o[86] = i[86];
  assign o[85] = i[85];
  assign o[84] = i[84];
  assign o[83] = i[83];
  assign o[82] = i[82];
  assign o[81] = i[81];
  assign o[80] = i[80];
  assign o[79] = i[79];
  assign o[78] = i[78];
  assign o[77] = i[77];
  assign o[76] = i[76];
  assign o[75] = i[75];
  assign o[74] = i[74];
  assign o[73] = i[73];
  assign o[72] = i[72];
  assign o[71] = i[71];
  assign o[70] = i[70];
  assign o[69] = i[69];
  assign o[68] = i[68];
  assign o[67] = i[67];
  assign o[66] = i[66];
  assign o[65] = i[65];
  assign o[64] = i[64];
  assign o[63] = i[63];
  assign o[62] = i[62];
  assign o[61] = i[61];
  assign o[60] = i[60];
  assign o[59] = i[59];
  assign o[58] = i[58];
  assign o[57] = i[57];
  assign o[56] = i[56];
  assign o[55] = i[55];
  assign o[54] = i[54];
  assign o[53] = i[53];
  assign o[52] = i[52];
  assign o[51] = i[51];
  assign o[50] = i[50];
  assign o[49] = i[49];
  assign o[48] = i[48];
  assign o[47] = i[47];
  assign o[46] = i[46];
  assign o[45] = i[45];
  assign o[44] = i[44];
  assign o[43] = i[43];
  assign o[42] = i[42];
  assign o[41] = i[41];
  assign o[40] = i[40];
  assign o[39] = i[39];
  assign o[38] = i[38];
  assign o[37] = i[37];
  assign o[36] = i[36];
  assign o[35] = i[35];
  assign o[34] = i[34];
  assign o[33] = i[33];
  assign o[32] = i[32];
  assign o[31] = i[31];
  assign o[30] = i[30];
  assign o[29] = i[29];
  assign o[28] = i[28];
  assign o[27] = i[27];
  assign o[26] = i[26];
  assign o[25] = i[25];
  assign o[24] = i[24];
  assign o[23] = i[23];
  assign o[22] = i[22];
  assign o[21] = i[21];
  assign o[20] = i[20];
  assign o[19] = i[19];
  assign o[18] = i[18];
  assign o[17] = i[17];
  assign o[16] = i[16];
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_rotate_right_width_p10
(
  data_i,
  rot_i,
  o
);

  input [9:0] data_i;
  input [3:0] rot_i;
  output [9:0] o;
  wire [9:0] o;
  wire SYNOPSYS_UNCONNECTED_1,SYNOPSYS_UNCONNECTED_2,SYNOPSYS_UNCONNECTED_3,
  SYNOPSYS_UNCONNECTED_4,SYNOPSYS_UNCONNECTED_5,SYNOPSYS_UNCONNECTED_6,
  SYNOPSYS_UNCONNECTED_7,SYNOPSYS_UNCONNECTED_8,SYNOPSYS_UNCONNECTED_9,SYNOPSYS_UNCONNECTED_10;
  assign { SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, o } = { data_i, data_i } >> rot_i;

endmodule



module bsg_circular_ptr_slots_p10_max_add_p10
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [3:0] add_i;
  output [3:0] o;
  output [3:0] n_o;
  input clk;
  input reset_i;
  wire [3:0] n_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;
  wire [4:0] ptr_wrap;
  reg [3:0] o;
  assign { N17, N16, N15, N14 } = o + add_i;
  assign { N13, N12, N11, N10, N9 } = o - { 1'b1, 1'b0, 1'b1, 1'b0 };
  assign ptr_wrap = { N13, N12, N11, N10, N9 } + add_i;
  assign { N8, N7, N6, N5 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N1)? n_o : 1'b0;
  assign N0 = reset_i;
  assign N1 = N4;
  assign n_o = (N2)? ptr_wrap[3:0] : 
               (N3)? { N17, N16, N15, N14 } : 1'b0;
  assign N2 = N18;
  assign N3 = ptr_wrap[4];
  assign N4 = ~reset_i;
  assign N18 = ~ptr_wrap[4];

  always @(posedge clk) begin
    if(1'b1) begin
      { o[3:0] } <= { N8, N7, N6, N5 };
    end 
  end


endmodule



module bsg_rr_f2f_input_width_p64_num_in_p10_middle_meet_p10
(
  clk,
  reset,
  valid_i,
  data_i,
  data_head_o,
  valid_head_o,
  go_channels_i,
  go_cnt_i,
  yumi_o
);

  input [9:0] valid_i;
  input [639:0] data_i;
  output [639:0] data_head_o;
  output [9:0] valid_head_o;
  input [9:0] go_channels_i;
  input [3:0] go_cnt_i;
  output [9:0] yumi_o;
  input clk;
  input reset;
  wire [639:0] data_head_o,data_head_o_flat_pretrunc;
  wire [9:0] valid_head_o,yumi_o;
  wire SYNOPSYS_UNCONNECTED_1,SYNOPSYS_UNCONNECTED_2,SYNOPSYS_UNCONNECTED_3,
  SYNOPSYS_UNCONNECTED_4,SYNOPSYS_UNCONNECTED_5,SYNOPSYS_UNCONNECTED_6,
  SYNOPSYS_UNCONNECTED_7,SYNOPSYS_UNCONNECTED_8,SYNOPSYS_UNCONNECTED_9,SYNOPSYS_UNCONNECTED_10,
  SYNOPSYS_UNCONNECTED_11,SYNOPSYS_UNCONNECTED_12,SYNOPSYS_UNCONNECTED_13,
  SYNOPSYS_UNCONNECTED_14,SYNOPSYS_UNCONNECTED_15,SYNOPSYS_UNCONNECTED_16,SYNOPSYS_UNCONNECTED_17,
  SYNOPSYS_UNCONNECTED_18,SYNOPSYS_UNCONNECTED_19,SYNOPSYS_UNCONNECTED_20,
  SYNOPSYS_UNCONNECTED_21,SYNOPSYS_UNCONNECTED_22,SYNOPSYS_UNCONNECTED_23,
  SYNOPSYS_UNCONNECTED_24,SYNOPSYS_UNCONNECTED_25,SYNOPSYS_UNCONNECTED_26,SYNOPSYS_UNCONNECTED_27,
  SYNOPSYS_UNCONNECTED_28,SYNOPSYS_UNCONNECTED_29,SYNOPSYS_UNCONNECTED_30,
  SYNOPSYS_UNCONNECTED_31,SYNOPSYS_UNCONNECTED_32,SYNOPSYS_UNCONNECTED_33,
  SYNOPSYS_UNCONNECTED_34,SYNOPSYS_UNCONNECTED_35,SYNOPSYS_UNCONNECTED_36,SYNOPSYS_UNCONNECTED_37,
  SYNOPSYS_UNCONNECTED_38,SYNOPSYS_UNCONNECTED_39,SYNOPSYS_UNCONNECTED_40,
  SYNOPSYS_UNCONNECTED_41,SYNOPSYS_UNCONNECTED_42,SYNOPSYS_UNCONNECTED_43,
  SYNOPSYS_UNCONNECTED_44,SYNOPSYS_UNCONNECTED_45,SYNOPSYS_UNCONNECTED_46,SYNOPSYS_UNCONNECTED_47,
  SYNOPSYS_UNCONNECTED_48,SYNOPSYS_UNCONNECTED_49,SYNOPSYS_UNCONNECTED_50,
  SYNOPSYS_UNCONNECTED_51,SYNOPSYS_UNCONNECTED_52,SYNOPSYS_UNCONNECTED_53,
  SYNOPSYS_UNCONNECTED_54,SYNOPSYS_UNCONNECTED_55,SYNOPSYS_UNCONNECTED_56,SYNOPSYS_UNCONNECTED_57,
  SYNOPSYS_UNCONNECTED_58,SYNOPSYS_UNCONNECTED_59,SYNOPSYS_UNCONNECTED_60,
  SYNOPSYS_UNCONNECTED_61,SYNOPSYS_UNCONNECTED_62,SYNOPSYS_UNCONNECTED_63,
  SYNOPSYS_UNCONNECTED_64,SYNOPSYS_UNCONNECTED_65,SYNOPSYS_UNCONNECTED_66,SYNOPSYS_UNCONNECTED_67,
  SYNOPSYS_UNCONNECTED_68,SYNOPSYS_UNCONNECTED_69,SYNOPSYS_UNCONNECTED_70,
  SYNOPSYS_UNCONNECTED_71,SYNOPSYS_UNCONNECTED_72,SYNOPSYS_UNCONNECTED_73,
  SYNOPSYS_UNCONNECTED_74,SYNOPSYS_UNCONNECTED_75,SYNOPSYS_UNCONNECTED_76,SYNOPSYS_UNCONNECTED_77,
  SYNOPSYS_UNCONNECTED_78,SYNOPSYS_UNCONNECTED_79,SYNOPSYS_UNCONNECTED_80,
  SYNOPSYS_UNCONNECTED_81,SYNOPSYS_UNCONNECTED_82,SYNOPSYS_UNCONNECTED_83,
  SYNOPSYS_UNCONNECTED_84,SYNOPSYS_UNCONNECTED_85,SYNOPSYS_UNCONNECTED_86,SYNOPSYS_UNCONNECTED_87,
  SYNOPSYS_UNCONNECTED_88,SYNOPSYS_UNCONNECTED_89,SYNOPSYS_UNCONNECTED_90,
  SYNOPSYS_UNCONNECTED_91,SYNOPSYS_UNCONNECTED_92,SYNOPSYS_UNCONNECTED_93,
  SYNOPSYS_UNCONNECTED_94,SYNOPSYS_UNCONNECTED_95,SYNOPSYS_UNCONNECTED_96,SYNOPSYS_UNCONNECTED_97,
  SYNOPSYS_UNCONNECTED_98,SYNOPSYS_UNCONNECTED_99,SYNOPSYS_UNCONNECTED_100,
  SYNOPSYS_UNCONNECTED_101,SYNOPSYS_UNCONNECTED_102,SYNOPSYS_UNCONNECTED_103,
  SYNOPSYS_UNCONNECTED_104,SYNOPSYS_UNCONNECTED_105,SYNOPSYS_UNCONNECTED_106,
  SYNOPSYS_UNCONNECTED_107,SYNOPSYS_UNCONNECTED_108,SYNOPSYS_UNCONNECTED_109,
  SYNOPSYS_UNCONNECTED_110,SYNOPSYS_UNCONNECTED_111,SYNOPSYS_UNCONNECTED_112,SYNOPSYS_UNCONNECTED_113,
  SYNOPSYS_UNCONNECTED_114,SYNOPSYS_UNCONNECTED_115,SYNOPSYS_UNCONNECTED_116,
  SYNOPSYS_UNCONNECTED_117,SYNOPSYS_UNCONNECTED_118,SYNOPSYS_UNCONNECTED_119,
  SYNOPSYS_UNCONNECTED_120,SYNOPSYS_UNCONNECTED_121,SYNOPSYS_UNCONNECTED_122,
  SYNOPSYS_UNCONNECTED_123,SYNOPSYS_UNCONNECTED_124,SYNOPSYS_UNCONNECTED_125,
  SYNOPSYS_UNCONNECTED_126,SYNOPSYS_UNCONNECTED_127,SYNOPSYS_UNCONNECTED_128,SYNOPSYS_UNCONNECTED_129,
  SYNOPSYS_UNCONNECTED_130,SYNOPSYS_UNCONNECTED_131,SYNOPSYS_UNCONNECTED_132,
  SYNOPSYS_UNCONNECTED_133,SYNOPSYS_UNCONNECTED_134,SYNOPSYS_UNCONNECTED_135,
  SYNOPSYS_UNCONNECTED_136,SYNOPSYS_UNCONNECTED_137,SYNOPSYS_UNCONNECTED_138,
  SYNOPSYS_UNCONNECTED_139,SYNOPSYS_UNCONNECTED_140,SYNOPSYS_UNCONNECTED_141,
  SYNOPSYS_UNCONNECTED_142,SYNOPSYS_UNCONNECTED_143,SYNOPSYS_UNCONNECTED_144,SYNOPSYS_UNCONNECTED_145,
  SYNOPSYS_UNCONNECTED_146,SYNOPSYS_UNCONNECTED_147,SYNOPSYS_UNCONNECTED_148,
  SYNOPSYS_UNCONNECTED_149,SYNOPSYS_UNCONNECTED_150,SYNOPSYS_UNCONNECTED_151,
  SYNOPSYS_UNCONNECTED_152,SYNOPSYS_UNCONNECTED_153,SYNOPSYS_UNCONNECTED_154,
  SYNOPSYS_UNCONNECTED_155,SYNOPSYS_UNCONNECTED_156,SYNOPSYS_UNCONNECTED_157,
  SYNOPSYS_UNCONNECTED_158,SYNOPSYS_UNCONNECTED_159,SYNOPSYS_UNCONNECTED_160,SYNOPSYS_UNCONNECTED_161,
  SYNOPSYS_UNCONNECTED_162,SYNOPSYS_UNCONNECTED_163,SYNOPSYS_UNCONNECTED_164,
  SYNOPSYS_UNCONNECTED_165,SYNOPSYS_UNCONNECTED_166,SYNOPSYS_UNCONNECTED_167,
  SYNOPSYS_UNCONNECTED_168,SYNOPSYS_UNCONNECTED_169,SYNOPSYS_UNCONNECTED_170,
  SYNOPSYS_UNCONNECTED_171,SYNOPSYS_UNCONNECTED_172,SYNOPSYS_UNCONNECTED_173,
  SYNOPSYS_UNCONNECTED_174,SYNOPSYS_UNCONNECTED_175,SYNOPSYS_UNCONNECTED_176,SYNOPSYS_UNCONNECTED_177,
  SYNOPSYS_UNCONNECTED_178,SYNOPSYS_UNCONNECTED_179,SYNOPSYS_UNCONNECTED_180,
  SYNOPSYS_UNCONNECTED_181,SYNOPSYS_UNCONNECTED_182,SYNOPSYS_UNCONNECTED_183,
  SYNOPSYS_UNCONNECTED_184,SYNOPSYS_UNCONNECTED_185,SYNOPSYS_UNCONNECTED_186,
  SYNOPSYS_UNCONNECTED_187,SYNOPSYS_UNCONNECTED_188,SYNOPSYS_UNCONNECTED_189,
  SYNOPSYS_UNCONNECTED_190,SYNOPSYS_UNCONNECTED_191,SYNOPSYS_UNCONNECTED_192,SYNOPSYS_UNCONNECTED_193,
  SYNOPSYS_UNCONNECTED_194,SYNOPSYS_UNCONNECTED_195,SYNOPSYS_UNCONNECTED_196,
  SYNOPSYS_UNCONNECTED_197,SYNOPSYS_UNCONNECTED_198,SYNOPSYS_UNCONNECTED_199,
  SYNOPSYS_UNCONNECTED_200,SYNOPSYS_UNCONNECTED_201,SYNOPSYS_UNCONNECTED_202,
  SYNOPSYS_UNCONNECTED_203,SYNOPSYS_UNCONNECTED_204,SYNOPSYS_UNCONNECTED_205,
  SYNOPSYS_UNCONNECTED_206,SYNOPSYS_UNCONNECTED_207,SYNOPSYS_UNCONNECTED_208,SYNOPSYS_UNCONNECTED_209,
  SYNOPSYS_UNCONNECTED_210,SYNOPSYS_UNCONNECTED_211,SYNOPSYS_UNCONNECTED_212,
  SYNOPSYS_UNCONNECTED_213,SYNOPSYS_UNCONNECTED_214,SYNOPSYS_UNCONNECTED_215,
  SYNOPSYS_UNCONNECTED_216,SYNOPSYS_UNCONNECTED_217,SYNOPSYS_UNCONNECTED_218,
  SYNOPSYS_UNCONNECTED_219,SYNOPSYS_UNCONNECTED_220,SYNOPSYS_UNCONNECTED_221,
  SYNOPSYS_UNCONNECTED_222,SYNOPSYS_UNCONNECTED_223,SYNOPSYS_UNCONNECTED_224,SYNOPSYS_UNCONNECTED_225,
  SYNOPSYS_UNCONNECTED_226,SYNOPSYS_UNCONNECTED_227,SYNOPSYS_UNCONNECTED_228,
  SYNOPSYS_UNCONNECTED_229,SYNOPSYS_UNCONNECTED_230,SYNOPSYS_UNCONNECTED_231,
  SYNOPSYS_UNCONNECTED_232,SYNOPSYS_UNCONNECTED_233,SYNOPSYS_UNCONNECTED_234,
  SYNOPSYS_UNCONNECTED_235,SYNOPSYS_UNCONNECTED_236,SYNOPSYS_UNCONNECTED_237,
  SYNOPSYS_UNCONNECTED_238,SYNOPSYS_UNCONNECTED_239,SYNOPSYS_UNCONNECTED_240,SYNOPSYS_UNCONNECTED_241,
  SYNOPSYS_UNCONNECTED_242,SYNOPSYS_UNCONNECTED_243,SYNOPSYS_UNCONNECTED_244,
  SYNOPSYS_UNCONNECTED_245,SYNOPSYS_UNCONNECTED_246,SYNOPSYS_UNCONNECTED_247,
  SYNOPSYS_UNCONNECTED_248,SYNOPSYS_UNCONNECTED_249,SYNOPSYS_UNCONNECTED_250,
  SYNOPSYS_UNCONNECTED_251,SYNOPSYS_UNCONNECTED_252,SYNOPSYS_UNCONNECTED_253,
  SYNOPSYS_UNCONNECTED_254,SYNOPSYS_UNCONNECTED_255,SYNOPSYS_UNCONNECTED_256,SYNOPSYS_UNCONNECTED_257,
  SYNOPSYS_UNCONNECTED_258,SYNOPSYS_UNCONNECTED_259,SYNOPSYS_UNCONNECTED_260,
  SYNOPSYS_UNCONNECTED_261,SYNOPSYS_UNCONNECTED_262,SYNOPSYS_UNCONNECTED_263,
  SYNOPSYS_UNCONNECTED_264,SYNOPSYS_UNCONNECTED_265,SYNOPSYS_UNCONNECTED_266,
  SYNOPSYS_UNCONNECTED_267,SYNOPSYS_UNCONNECTED_268,SYNOPSYS_UNCONNECTED_269,
  SYNOPSYS_UNCONNECTED_270,SYNOPSYS_UNCONNECTED_271,SYNOPSYS_UNCONNECTED_272,SYNOPSYS_UNCONNECTED_273,
  SYNOPSYS_UNCONNECTED_274,SYNOPSYS_UNCONNECTED_275,SYNOPSYS_UNCONNECTED_276,
  SYNOPSYS_UNCONNECTED_277,SYNOPSYS_UNCONNECTED_278,SYNOPSYS_UNCONNECTED_279,
  SYNOPSYS_UNCONNECTED_280,SYNOPSYS_UNCONNECTED_281,SYNOPSYS_UNCONNECTED_282,
  SYNOPSYS_UNCONNECTED_283,SYNOPSYS_UNCONNECTED_284,SYNOPSYS_UNCONNECTED_285,
  SYNOPSYS_UNCONNECTED_286,SYNOPSYS_UNCONNECTED_287,SYNOPSYS_UNCONNECTED_288,SYNOPSYS_UNCONNECTED_289,
  SYNOPSYS_UNCONNECTED_290,SYNOPSYS_UNCONNECTED_291,SYNOPSYS_UNCONNECTED_292,
  SYNOPSYS_UNCONNECTED_293,SYNOPSYS_UNCONNECTED_294,SYNOPSYS_UNCONNECTED_295,
  SYNOPSYS_UNCONNECTED_296,SYNOPSYS_UNCONNECTED_297,SYNOPSYS_UNCONNECTED_298,
  SYNOPSYS_UNCONNECTED_299,SYNOPSYS_UNCONNECTED_300,SYNOPSYS_UNCONNECTED_301,
  SYNOPSYS_UNCONNECTED_302,SYNOPSYS_UNCONNECTED_303,SYNOPSYS_UNCONNECTED_304,SYNOPSYS_UNCONNECTED_305,
  SYNOPSYS_UNCONNECTED_306,SYNOPSYS_UNCONNECTED_307,SYNOPSYS_UNCONNECTED_308,
  SYNOPSYS_UNCONNECTED_309,SYNOPSYS_UNCONNECTED_310,SYNOPSYS_UNCONNECTED_311,
  SYNOPSYS_UNCONNECTED_312,SYNOPSYS_UNCONNECTED_313,SYNOPSYS_UNCONNECTED_314,
  SYNOPSYS_UNCONNECTED_315,SYNOPSYS_UNCONNECTED_316,SYNOPSYS_UNCONNECTED_317,
  SYNOPSYS_UNCONNECTED_318,SYNOPSYS_UNCONNECTED_319,SYNOPSYS_UNCONNECTED_320,SYNOPSYS_UNCONNECTED_321,
  SYNOPSYS_UNCONNECTED_322,SYNOPSYS_UNCONNECTED_323,SYNOPSYS_UNCONNECTED_324,
  SYNOPSYS_UNCONNECTED_325,SYNOPSYS_UNCONNECTED_326,SYNOPSYS_UNCONNECTED_327,
  SYNOPSYS_UNCONNECTED_328,SYNOPSYS_UNCONNECTED_329,SYNOPSYS_UNCONNECTED_330,
  SYNOPSYS_UNCONNECTED_331,SYNOPSYS_UNCONNECTED_332,SYNOPSYS_UNCONNECTED_333,
  SYNOPSYS_UNCONNECTED_334,SYNOPSYS_UNCONNECTED_335,SYNOPSYS_UNCONNECTED_336,SYNOPSYS_UNCONNECTED_337,
  SYNOPSYS_UNCONNECTED_338,SYNOPSYS_UNCONNECTED_339,SYNOPSYS_UNCONNECTED_340,
  SYNOPSYS_UNCONNECTED_341,SYNOPSYS_UNCONNECTED_342,SYNOPSYS_UNCONNECTED_343,
  SYNOPSYS_UNCONNECTED_344,SYNOPSYS_UNCONNECTED_345,SYNOPSYS_UNCONNECTED_346,
  SYNOPSYS_UNCONNECTED_347,SYNOPSYS_UNCONNECTED_348,SYNOPSYS_UNCONNECTED_349,
  SYNOPSYS_UNCONNECTED_350,SYNOPSYS_UNCONNECTED_351,SYNOPSYS_UNCONNECTED_352,SYNOPSYS_UNCONNECTED_353,
  SYNOPSYS_UNCONNECTED_354,SYNOPSYS_UNCONNECTED_355,SYNOPSYS_UNCONNECTED_356,
  SYNOPSYS_UNCONNECTED_357,SYNOPSYS_UNCONNECTED_358,SYNOPSYS_UNCONNECTED_359,
  SYNOPSYS_UNCONNECTED_360,SYNOPSYS_UNCONNECTED_361,SYNOPSYS_UNCONNECTED_362,
  SYNOPSYS_UNCONNECTED_363,SYNOPSYS_UNCONNECTED_364,SYNOPSYS_UNCONNECTED_365,
  SYNOPSYS_UNCONNECTED_366,SYNOPSYS_UNCONNECTED_367,SYNOPSYS_UNCONNECTED_368,SYNOPSYS_UNCONNECTED_369,
  SYNOPSYS_UNCONNECTED_370,SYNOPSYS_UNCONNECTED_371,SYNOPSYS_UNCONNECTED_372,
  SYNOPSYS_UNCONNECTED_373,SYNOPSYS_UNCONNECTED_374,SYNOPSYS_UNCONNECTED_375,
  SYNOPSYS_UNCONNECTED_376,SYNOPSYS_UNCONNECTED_377,SYNOPSYS_UNCONNECTED_378,
  SYNOPSYS_UNCONNECTED_379,SYNOPSYS_UNCONNECTED_380,SYNOPSYS_UNCONNECTED_381,
  SYNOPSYS_UNCONNECTED_382,SYNOPSYS_UNCONNECTED_383,SYNOPSYS_UNCONNECTED_384,SYNOPSYS_UNCONNECTED_385,
  SYNOPSYS_UNCONNECTED_386,SYNOPSYS_UNCONNECTED_387,SYNOPSYS_UNCONNECTED_388,
  SYNOPSYS_UNCONNECTED_389,SYNOPSYS_UNCONNECTED_390,SYNOPSYS_UNCONNECTED_391,
  SYNOPSYS_UNCONNECTED_392,SYNOPSYS_UNCONNECTED_393,SYNOPSYS_UNCONNECTED_394,
  SYNOPSYS_UNCONNECTED_395,SYNOPSYS_UNCONNECTED_396,SYNOPSYS_UNCONNECTED_397,
  SYNOPSYS_UNCONNECTED_398,SYNOPSYS_UNCONNECTED_399,SYNOPSYS_UNCONNECTED_400,SYNOPSYS_UNCONNECTED_401,
  SYNOPSYS_UNCONNECTED_402,SYNOPSYS_UNCONNECTED_403,SYNOPSYS_UNCONNECTED_404,
  SYNOPSYS_UNCONNECTED_405,SYNOPSYS_UNCONNECTED_406,SYNOPSYS_UNCONNECTED_407,
  SYNOPSYS_UNCONNECTED_408,SYNOPSYS_UNCONNECTED_409,SYNOPSYS_UNCONNECTED_410,
  SYNOPSYS_UNCONNECTED_411,SYNOPSYS_UNCONNECTED_412,SYNOPSYS_UNCONNECTED_413,
  SYNOPSYS_UNCONNECTED_414,SYNOPSYS_UNCONNECTED_415,SYNOPSYS_UNCONNECTED_416,SYNOPSYS_UNCONNECTED_417,
  SYNOPSYS_UNCONNECTED_418,SYNOPSYS_UNCONNECTED_419,SYNOPSYS_UNCONNECTED_420,
  SYNOPSYS_UNCONNECTED_421,SYNOPSYS_UNCONNECTED_422,SYNOPSYS_UNCONNECTED_423,
  SYNOPSYS_UNCONNECTED_424,SYNOPSYS_UNCONNECTED_425,SYNOPSYS_UNCONNECTED_426,
  SYNOPSYS_UNCONNECTED_427,SYNOPSYS_UNCONNECTED_428,SYNOPSYS_UNCONNECTED_429,
  SYNOPSYS_UNCONNECTED_430,SYNOPSYS_UNCONNECTED_431,SYNOPSYS_UNCONNECTED_432,SYNOPSYS_UNCONNECTED_433,
  SYNOPSYS_UNCONNECTED_434,SYNOPSYS_UNCONNECTED_435,SYNOPSYS_UNCONNECTED_436,
  SYNOPSYS_UNCONNECTED_437,SYNOPSYS_UNCONNECTED_438,SYNOPSYS_UNCONNECTED_439,
  SYNOPSYS_UNCONNECTED_440,SYNOPSYS_UNCONNECTED_441,SYNOPSYS_UNCONNECTED_442,
  SYNOPSYS_UNCONNECTED_443,SYNOPSYS_UNCONNECTED_444,SYNOPSYS_UNCONNECTED_445,
  SYNOPSYS_UNCONNECTED_446,SYNOPSYS_UNCONNECTED_447,SYNOPSYS_UNCONNECTED_448,SYNOPSYS_UNCONNECTED_449,
  SYNOPSYS_UNCONNECTED_450,SYNOPSYS_UNCONNECTED_451,SYNOPSYS_UNCONNECTED_452,
  SYNOPSYS_UNCONNECTED_453,SYNOPSYS_UNCONNECTED_454,SYNOPSYS_UNCONNECTED_455,
  SYNOPSYS_UNCONNECTED_456,SYNOPSYS_UNCONNECTED_457,SYNOPSYS_UNCONNECTED_458,
  SYNOPSYS_UNCONNECTED_459,SYNOPSYS_UNCONNECTED_460,SYNOPSYS_UNCONNECTED_461,
  SYNOPSYS_UNCONNECTED_462,SYNOPSYS_UNCONNECTED_463,SYNOPSYS_UNCONNECTED_464,SYNOPSYS_UNCONNECTED_465,
  SYNOPSYS_UNCONNECTED_466,SYNOPSYS_UNCONNECTED_467,SYNOPSYS_UNCONNECTED_468,
  SYNOPSYS_UNCONNECTED_469,SYNOPSYS_UNCONNECTED_470,SYNOPSYS_UNCONNECTED_471,
  SYNOPSYS_UNCONNECTED_472,SYNOPSYS_UNCONNECTED_473,SYNOPSYS_UNCONNECTED_474,
  SYNOPSYS_UNCONNECTED_475,SYNOPSYS_UNCONNECTED_476,SYNOPSYS_UNCONNECTED_477,
  SYNOPSYS_UNCONNECTED_478,SYNOPSYS_UNCONNECTED_479,SYNOPSYS_UNCONNECTED_480,SYNOPSYS_UNCONNECTED_481,
  SYNOPSYS_UNCONNECTED_482,SYNOPSYS_UNCONNECTED_483,SYNOPSYS_UNCONNECTED_484,
  SYNOPSYS_UNCONNECTED_485,SYNOPSYS_UNCONNECTED_486,SYNOPSYS_UNCONNECTED_487,
  SYNOPSYS_UNCONNECTED_488,SYNOPSYS_UNCONNECTED_489,SYNOPSYS_UNCONNECTED_490,
  SYNOPSYS_UNCONNECTED_491,SYNOPSYS_UNCONNECTED_492,SYNOPSYS_UNCONNECTED_493,
  SYNOPSYS_UNCONNECTED_494,SYNOPSYS_UNCONNECTED_495,SYNOPSYS_UNCONNECTED_496,SYNOPSYS_UNCONNECTED_497,
  SYNOPSYS_UNCONNECTED_498,SYNOPSYS_UNCONNECTED_499,SYNOPSYS_UNCONNECTED_500,
  SYNOPSYS_UNCONNECTED_501,SYNOPSYS_UNCONNECTED_502,SYNOPSYS_UNCONNECTED_503,
  SYNOPSYS_UNCONNECTED_504,SYNOPSYS_UNCONNECTED_505,SYNOPSYS_UNCONNECTED_506,
  SYNOPSYS_UNCONNECTED_507,SYNOPSYS_UNCONNECTED_508,SYNOPSYS_UNCONNECTED_509,
  SYNOPSYS_UNCONNECTED_510,SYNOPSYS_UNCONNECTED_511,SYNOPSYS_UNCONNECTED_512,SYNOPSYS_UNCONNECTED_513,
  SYNOPSYS_UNCONNECTED_514,SYNOPSYS_UNCONNECTED_515,SYNOPSYS_UNCONNECTED_516,
  SYNOPSYS_UNCONNECTED_517,SYNOPSYS_UNCONNECTED_518,SYNOPSYS_UNCONNECTED_519,
  SYNOPSYS_UNCONNECTED_520,SYNOPSYS_UNCONNECTED_521,SYNOPSYS_UNCONNECTED_522,
  SYNOPSYS_UNCONNECTED_523,SYNOPSYS_UNCONNECTED_524,SYNOPSYS_UNCONNECTED_525,
  SYNOPSYS_UNCONNECTED_526,SYNOPSYS_UNCONNECTED_527,SYNOPSYS_UNCONNECTED_528,SYNOPSYS_UNCONNECTED_529,
  SYNOPSYS_UNCONNECTED_530,SYNOPSYS_UNCONNECTED_531,SYNOPSYS_UNCONNECTED_532,
  SYNOPSYS_UNCONNECTED_533,SYNOPSYS_UNCONNECTED_534,SYNOPSYS_UNCONNECTED_535,
  SYNOPSYS_UNCONNECTED_536,SYNOPSYS_UNCONNECTED_537,SYNOPSYS_UNCONNECTED_538,
  SYNOPSYS_UNCONNECTED_539,SYNOPSYS_UNCONNECTED_540,SYNOPSYS_UNCONNECTED_541,
  SYNOPSYS_UNCONNECTED_542,SYNOPSYS_UNCONNECTED_543,SYNOPSYS_UNCONNECTED_544,SYNOPSYS_UNCONNECTED_545,
  SYNOPSYS_UNCONNECTED_546,SYNOPSYS_UNCONNECTED_547,SYNOPSYS_UNCONNECTED_548,
  SYNOPSYS_UNCONNECTED_549,SYNOPSYS_UNCONNECTED_550,SYNOPSYS_UNCONNECTED_551,
  SYNOPSYS_UNCONNECTED_552,SYNOPSYS_UNCONNECTED_553,SYNOPSYS_UNCONNECTED_554,
  SYNOPSYS_UNCONNECTED_555,SYNOPSYS_UNCONNECTED_556,SYNOPSYS_UNCONNECTED_557,
  SYNOPSYS_UNCONNECTED_558,SYNOPSYS_UNCONNECTED_559,SYNOPSYS_UNCONNECTED_560,SYNOPSYS_UNCONNECTED_561,
  SYNOPSYS_UNCONNECTED_562,SYNOPSYS_UNCONNECTED_563,SYNOPSYS_UNCONNECTED_564,
  SYNOPSYS_UNCONNECTED_565,SYNOPSYS_UNCONNECTED_566,SYNOPSYS_UNCONNECTED_567,
  SYNOPSYS_UNCONNECTED_568,SYNOPSYS_UNCONNECTED_569,SYNOPSYS_UNCONNECTED_570,
  SYNOPSYS_UNCONNECTED_571,SYNOPSYS_UNCONNECTED_572,SYNOPSYS_UNCONNECTED_573,
  SYNOPSYS_UNCONNECTED_574,SYNOPSYS_UNCONNECTED_575,SYNOPSYS_UNCONNECTED_576,SYNOPSYS_UNCONNECTED_577,
  SYNOPSYS_UNCONNECTED_578,SYNOPSYS_UNCONNECTED_579,SYNOPSYS_UNCONNECTED_580,
  SYNOPSYS_UNCONNECTED_581,SYNOPSYS_UNCONNECTED_582,SYNOPSYS_UNCONNECTED_583,
  SYNOPSYS_UNCONNECTED_584,SYNOPSYS_UNCONNECTED_585,SYNOPSYS_UNCONNECTED_586,
  SYNOPSYS_UNCONNECTED_587,SYNOPSYS_UNCONNECTED_588,SYNOPSYS_UNCONNECTED_589,
  SYNOPSYS_UNCONNECTED_590,SYNOPSYS_UNCONNECTED_591,SYNOPSYS_UNCONNECTED_592,SYNOPSYS_UNCONNECTED_593,
  SYNOPSYS_UNCONNECTED_594,SYNOPSYS_UNCONNECTED_595,SYNOPSYS_UNCONNECTED_596,
  SYNOPSYS_UNCONNECTED_597,SYNOPSYS_UNCONNECTED_598,SYNOPSYS_UNCONNECTED_599,
  SYNOPSYS_UNCONNECTED_600,SYNOPSYS_UNCONNECTED_601,SYNOPSYS_UNCONNECTED_602,
  SYNOPSYS_UNCONNECTED_603,SYNOPSYS_UNCONNECTED_604,SYNOPSYS_UNCONNECTED_605,
  SYNOPSYS_UNCONNECTED_606,SYNOPSYS_UNCONNECTED_607,SYNOPSYS_UNCONNECTED_608,SYNOPSYS_UNCONNECTED_609,
  SYNOPSYS_UNCONNECTED_610,SYNOPSYS_UNCONNECTED_611,SYNOPSYS_UNCONNECTED_612,
  SYNOPSYS_UNCONNECTED_613,SYNOPSYS_UNCONNECTED_614,SYNOPSYS_UNCONNECTED_615,
  SYNOPSYS_UNCONNECTED_616,SYNOPSYS_UNCONNECTED_617,SYNOPSYS_UNCONNECTED_618,
  SYNOPSYS_UNCONNECTED_619,SYNOPSYS_UNCONNECTED_620,SYNOPSYS_UNCONNECTED_621,
  SYNOPSYS_UNCONNECTED_622,SYNOPSYS_UNCONNECTED_623,SYNOPSYS_UNCONNECTED_624,SYNOPSYS_UNCONNECTED_625,
  SYNOPSYS_UNCONNECTED_626,SYNOPSYS_UNCONNECTED_627,SYNOPSYS_UNCONNECTED_628,
  SYNOPSYS_UNCONNECTED_629,SYNOPSYS_UNCONNECTED_630,SYNOPSYS_UNCONNECTED_631,
  SYNOPSYS_UNCONNECTED_632,SYNOPSYS_UNCONNECTED_633,SYNOPSYS_UNCONNECTED_634,
  SYNOPSYS_UNCONNECTED_635,SYNOPSYS_UNCONNECTED_636,SYNOPSYS_UNCONNECTED_637,
  SYNOPSYS_UNCONNECTED_638,SYNOPSYS_UNCONNECTED_639,SYNOPSYS_UNCONNECTED_640,SYNOPSYS_UNCONNECTED_641,
  SYNOPSYS_UNCONNECTED_642,SYNOPSYS_UNCONNECTED_643,SYNOPSYS_UNCONNECTED_644,
  SYNOPSYS_UNCONNECTED_645,SYNOPSYS_UNCONNECTED_646,SYNOPSYS_UNCONNECTED_647,
  SYNOPSYS_UNCONNECTED_648,SYNOPSYS_UNCONNECTED_649,SYNOPSYS_UNCONNECTED_650,
  SYNOPSYS_UNCONNECTED_651,SYNOPSYS_UNCONNECTED_652,SYNOPSYS_UNCONNECTED_653,
  SYNOPSYS_UNCONNECTED_654,SYNOPSYS_UNCONNECTED_655,SYNOPSYS_UNCONNECTED_656,SYNOPSYS_UNCONNECTED_657,
  SYNOPSYS_UNCONNECTED_658;
  wire [3:0] iptr_r,iptr_r_data;

  bsg_make_2D_array_width_p64_items_p10
  bm2Da
  (
    .i(data_head_o_flat_pretrunc),
    .o(data_head_o)
  );


  bsg_rotate_right_width_p10
  valid_rr
  (
    .data_i(valid_i),
    .rot_i(iptr_r),
    .o(valid_head_o)
  );

  assign { SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306, SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340, SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342, SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366, SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368, SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370, SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372, SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374, SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413, SYNOPSYS_UNCONNECTED_414, SYNOPSYS_UNCONNECTED_415, SYNOPSYS_UNCONNECTED_416, SYNOPSYS_UNCONNECTED_417, SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_419, SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_421, SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_423, SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_425, SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_427, SYNOPSYS_UNCONNECTED_428, SYNOPSYS_UNCONNECTED_429, SYNOPSYS_UNCONNECTED_430, SYNOPSYS_UNCONNECTED_431, SYNOPSYS_UNCONNECTED_432, SYNOPSYS_UNCONNECTED_433, SYNOPSYS_UNCONNECTED_434, SYNOPSYS_UNCONNECTED_435, SYNOPSYS_UNCONNECTED_436, SYNOPSYS_UNCONNECTED_437, SYNOPSYS_UNCONNECTED_438, SYNOPSYS_UNCONNECTED_439, SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_441, SYNOPSYS_UNCONNECTED_442, SYNOPSYS_UNCONNECTED_443, SYNOPSYS_UNCONNECTED_444, SYNOPSYS_UNCONNECTED_445, SYNOPSYS_UNCONNECTED_446, SYNOPSYS_UNCONNECTED_447, SYNOPSYS_UNCONNECTED_448, SYNOPSYS_UNCONNECTED_449, SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_451, SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_453, SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_455, SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_457, SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_459, SYNOPSYS_UNCONNECTED_460, SYNOPSYS_UNCONNECTED_461, SYNOPSYS_UNCONNECTED_462, SYNOPSYS_UNCONNECTED_463, SYNOPSYS_UNCONNECTED_464, SYNOPSYS_UNCONNECTED_465, SYNOPSYS_UNCONNECTED_466, SYNOPSYS_UNCONNECTED_467, SYNOPSYS_UNCONNECTED_468, SYNOPSYS_UNCONNECTED_469, SYNOPSYS_UNCONNECTED_470, SYNOPSYS_UNCONNECTED_471, SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_473, SYNOPSYS_UNCONNECTED_474, SYNOPSYS_UNCONNECTED_475, SYNOPSYS_UNCONNECTED_476, SYNOPSYS_UNCONNECTED_477, SYNOPSYS_UNCONNECTED_478, SYNOPSYS_UNCONNECTED_479, SYNOPSYS_UNCONNECTED_480, SYNOPSYS_UNCONNECTED_481, SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_483, SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_485, SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_487, SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_489, SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_491, SYNOPSYS_UNCONNECTED_492, SYNOPSYS_UNCONNECTED_493, SYNOPSYS_UNCONNECTED_494, SYNOPSYS_UNCONNECTED_495, SYNOPSYS_UNCONNECTED_496, SYNOPSYS_UNCONNECTED_497, SYNOPSYS_UNCONNECTED_498, SYNOPSYS_UNCONNECTED_499, SYNOPSYS_UNCONNECTED_500, SYNOPSYS_UNCONNECTED_501, SYNOPSYS_UNCONNECTED_502, SYNOPSYS_UNCONNECTED_503, SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_505, SYNOPSYS_UNCONNECTED_506, SYNOPSYS_UNCONNECTED_507, SYNOPSYS_UNCONNECTED_508, SYNOPSYS_UNCONNECTED_509, SYNOPSYS_UNCONNECTED_510, SYNOPSYS_UNCONNECTED_511, SYNOPSYS_UNCONNECTED_512, SYNOPSYS_UNCONNECTED_513, SYNOPSYS_UNCONNECTED_514, SYNOPSYS_UNCONNECTED_515, SYNOPSYS_UNCONNECTED_516, SYNOPSYS_UNCONNECTED_517, SYNOPSYS_UNCONNECTED_518, SYNOPSYS_UNCONNECTED_519, SYNOPSYS_UNCONNECTED_520, SYNOPSYS_UNCONNECTED_521, SYNOPSYS_UNCONNECTED_522, SYNOPSYS_UNCONNECTED_523, SYNOPSYS_UNCONNECTED_524, SYNOPSYS_UNCONNECTED_525, SYNOPSYS_UNCONNECTED_526, SYNOPSYS_UNCONNECTED_527, SYNOPSYS_UNCONNECTED_528, SYNOPSYS_UNCONNECTED_529, SYNOPSYS_UNCONNECTED_530, SYNOPSYS_UNCONNECTED_531, SYNOPSYS_UNCONNECTED_532, SYNOPSYS_UNCONNECTED_533, SYNOPSYS_UNCONNECTED_534, SYNOPSYS_UNCONNECTED_535, SYNOPSYS_UNCONNECTED_536, SYNOPSYS_UNCONNECTED_537, SYNOPSYS_UNCONNECTED_538, SYNOPSYS_UNCONNECTED_539, SYNOPSYS_UNCONNECTED_540, SYNOPSYS_UNCONNECTED_541, SYNOPSYS_UNCONNECTED_542, SYNOPSYS_UNCONNECTED_543, SYNOPSYS_UNCONNECTED_544, SYNOPSYS_UNCONNECTED_545, SYNOPSYS_UNCONNECTED_546, SYNOPSYS_UNCONNECTED_547, SYNOPSYS_UNCONNECTED_548, SYNOPSYS_UNCONNECTED_549, SYNOPSYS_UNCONNECTED_550, SYNOPSYS_UNCONNECTED_551, SYNOPSYS_UNCONNECTED_552, SYNOPSYS_UNCONNECTED_553, SYNOPSYS_UNCONNECTED_554, SYNOPSYS_UNCONNECTED_555, SYNOPSYS_UNCONNECTED_556, SYNOPSYS_UNCONNECTED_557, SYNOPSYS_UNCONNECTED_558, SYNOPSYS_UNCONNECTED_559, SYNOPSYS_UNCONNECTED_560, SYNOPSYS_UNCONNECTED_561, SYNOPSYS_UNCONNECTED_562, SYNOPSYS_UNCONNECTED_563, SYNOPSYS_UNCONNECTED_564, SYNOPSYS_UNCONNECTED_565, SYNOPSYS_UNCONNECTED_566, SYNOPSYS_UNCONNECTED_567, SYNOPSYS_UNCONNECTED_568, SYNOPSYS_UNCONNECTED_569, SYNOPSYS_UNCONNECTED_570, SYNOPSYS_UNCONNECTED_571, SYNOPSYS_UNCONNECTED_572, SYNOPSYS_UNCONNECTED_573, SYNOPSYS_UNCONNECTED_574, SYNOPSYS_UNCONNECTED_575, SYNOPSYS_UNCONNECTED_576, SYNOPSYS_UNCONNECTED_577, SYNOPSYS_UNCONNECTED_578, SYNOPSYS_UNCONNECTED_579, SYNOPSYS_UNCONNECTED_580, SYNOPSYS_UNCONNECTED_581, SYNOPSYS_UNCONNECTED_582, SYNOPSYS_UNCONNECTED_583, SYNOPSYS_UNCONNECTED_584, SYNOPSYS_UNCONNECTED_585, SYNOPSYS_UNCONNECTED_586, SYNOPSYS_UNCONNECTED_587, SYNOPSYS_UNCONNECTED_588, SYNOPSYS_UNCONNECTED_589, SYNOPSYS_UNCONNECTED_590, SYNOPSYS_UNCONNECTED_591, SYNOPSYS_UNCONNECTED_592, SYNOPSYS_UNCONNECTED_593, SYNOPSYS_UNCONNECTED_594, SYNOPSYS_UNCONNECTED_595, SYNOPSYS_UNCONNECTED_596, SYNOPSYS_UNCONNECTED_597, SYNOPSYS_UNCONNECTED_598, SYNOPSYS_UNCONNECTED_599, SYNOPSYS_UNCONNECTED_600, SYNOPSYS_UNCONNECTED_601, SYNOPSYS_UNCONNECTED_602, SYNOPSYS_UNCONNECTED_603, SYNOPSYS_UNCONNECTED_604, SYNOPSYS_UNCONNECTED_605, SYNOPSYS_UNCONNECTED_606, SYNOPSYS_UNCONNECTED_607, SYNOPSYS_UNCONNECTED_608, SYNOPSYS_UNCONNECTED_609, SYNOPSYS_UNCONNECTED_610, SYNOPSYS_UNCONNECTED_611, SYNOPSYS_UNCONNECTED_612, SYNOPSYS_UNCONNECTED_613, SYNOPSYS_UNCONNECTED_614, SYNOPSYS_UNCONNECTED_615, SYNOPSYS_UNCONNECTED_616, SYNOPSYS_UNCONNECTED_617, SYNOPSYS_UNCONNECTED_618, SYNOPSYS_UNCONNECTED_619, SYNOPSYS_UNCONNECTED_620, SYNOPSYS_UNCONNECTED_621, SYNOPSYS_UNCONNECTED_622, SYNOPSYS_UNCONNECTED_623, SYNOPSYS_UNCONNECTED_624, SYNOPSYS_UNCONNECTED_625, SYNOPSYS_UNCONNECTED_626, SYNOPSYS_UNCONNECTED_627, SYNOPSYS_UNCONNECTED_628, SYNOPSYS_UNCONNECTED_629, SYNOPSYS_UNCONNECTED_630, SYNOPSYS_UNCONNECTED_631, SYNOPSYS_UNCONNECTED_632, SYNOPSYS_UNCONNECTED_633, SYNOPSYS_UNCONNECTED_634, SYNOPSYS_UNCONNECTED_635, SYNOPSYS_UNCONNECTED_636, SYNOPSYS_UNCONNECTED_637, SYNOPSYS_UNCONNECTED_638, SYNOPSYS_UNCONNECTED_639, SYNOPSYS_UNCONNECTED_640, data_head_o_flat_pretrunc } = { data_i, data_i } >> { iptr_r_data, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign { yumi_o, SYNOPSYS_UNCONNECTED_641, SYNOPSYS_UNCONNECTED_642, SYNOPSYS_UNCONNECTED_643, SYNOPSYS_UNCONNECTED_644, SYNOPSYS_UNCONNECTED_645, SYNOPSYS_UNCONNECTED_646, SYNOPSYS_UNCONNECTED_647, SYNOPSYS_UNCONNECTED_648, SYNOPSYS_UNCONNECTED_649, SYNOPSYS_UNCONNECTED_650 } = { go_channels_i, go_channels_i } << iptr_r;

  bsg_circular_ptr_slots_p10_max_add_p10
  c_ptr
  (
    .clk(clk),
    .reset_i(reset),
    .add_i(go_cnt_i),
    .o(iptr_r),
    .n_o({ SYNOPSYS_UNCONNECTED_651, SYNOPSYS_UNCONNECTED_652, SYNOPSYS_UNCONNECTED_653, SYNOPSYS_UNCONNECTED_654 })
  );


  bsg_circular_ptr_slots_p10_max_add_p10
  c_ptr_data
  (
    .clk(clk),
    .reset_i(reset),
    .add_i(go_cnt_i),
    .o(iptr_r_data),
    .n_o({ SYNOPSYS_UNCONNECTED_655, SYNOPSYS_UNCONNECTED_656, SYNOPSYS_UNCONNECTED_657, SYNOPSYS_UNCONNECTED_658 })
  );


endmodule



module bsg_scan_width_p10_and_p1_lo_to_hi_p1
(
  i,
  o
);

  input [9:0] i;
  output [9:0] o;
  wire [9:0] o;
  wire t_3__9_,t_3__8_,t_3__7_,t_3__6_,t_3__5_,t_3__4_,t_3__3_,t_3__2_,t_3__1_,t_3__0_,
  t_2__9_,t_2__8_,t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,
  t_1__9_,t_1__8_,t_1__7_,t_1__6_,t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__9_ = i[0] & 1'b1;
  assign t_1__8_ = i[1] & i[0];
  assign t_1__7_ = i[2] & i[1];
  assign t_1__6_ = i[3] & i[2];
  assign t_1__5_ = i[4] & i[3];
  assign t_1__4_ = i[5] & i[4];
  assign t_1__3_ = i[6] & i[5];
  assign t_1__2_ = i[7] & i[6];
  assign t_1__1_ = i[8] & i[7];
  assign t_1__0_ = i[9] & i[8];
  assign t_2__9_ = t_1__9_ & 1'b1;
  assign t_2__8_ = t_1__8_ & 1'b1;
  assign t_2__7_ = t_1__7_ & t_1__9_;
  assign t_2__6_ = t_1__6_ & t_1__8_;
  assign t_2__5_ = t_1__5_ & t_1__7_;
  assign t_2__4_ = t_1__4_ & t_1__6_;
  assign t_2__3_ = t_1__3_ & t_1__5_;
  assign t_2__2_ = t_1__2_ & t_1__4_;
  assign t_2__1_ = t_1__1_ & t_1__3_;
  assign t_2__0_ = t_1__0_ & t_1__2_;
  assign t_3__9_ = t_2__9_ & 1'b1;
  assign t_3__8_ = t_2__8_ & 1'b1;
  assign t_3__7_ = t_2__7_ & 1'b1;
  assign t_3__6_ = t_2__6_ & 1'b1;
  assign t_3__5_ = t_2__5_ & t_2__9_;
  assign t_3__4_ = t_2__4_ & t_2__8_;
  assign t_3__3_ = t_2__3_ & t_2__7_;
  assign t_3__2_ = t_2__2_ & t_2__6_;
  assign t_3__1_ = t_2__1_ & t_2__5_;
  assign t_3__0_ = t_2__0_ & t_2__4_;
  assign o[0] = t_3__9_ & 1'b1;
  assign o[1] = t_3__8_ & 1'b1;
  assign o[2] = t_3__7_ & 1'b1;
  assign o[3] = t_3__6_ & 1'b1;
  assign o[4] = t_3__5_ & 1'b1;
  assign o[5] = t_3__4_ & 1'b1;
  assign o[6] = t_3__3_ & 1'b1;
  assign o[7] = t_3__2_ & 1'b1;
  assign o[8] = t_3__1_ & t_3__9_;
  assign o[9] = t_3__0_ & t_3__8_;

endmodule



module bsg_encode_one_hot_width_p1
(
  i,
  addr_o,
  v_o
);

  input [0:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  assign v_o = i[0];
  assign addr_o[0] = 1'b0;

endmodule



module bsg_encode_one_hot_width_p2
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o,aligned_vs;
  wire v_o;
  wire [1:0] aligned_addrs;

  bsg_encode_one_hot_width_p1
  aligned_left
  (
    .i(i[0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p1
  aligned_right
  (
    .i(i[1]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[0])
  );

  assign v_o = addr_o[0] | aligned_vs[0];

endmodule



module bsg_encode_one_hot_width_p4
(
  i,
  addr_o,
  v_o
);

  input [3:0] i;
  output [1:0] addr_o;
  output v_o;
  wire [1:0] addr_o,aligned_addrs;
  wire v_o;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p2
  aligned_left
  (
    .i(i[1:0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p2
  aligned_right
  (
    .i(i[3:2]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[1])
  );

  assign v_o = addr_o[1] | aligned_vs[0];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[1];

endmodule



module bsg_encode_one_hot_width_p8
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [3:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p4
  aligned_left
  (
    .i(i[3:0]),
    .addr_o(aligned_addrs[1:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p4
  aligned_right
  (
    .i(i[7:4]),
    .addr_o(aligned_addrs[3:2]),
    .v_o(addr_o[2])
  );

  assign v_o = addr_o[2] | aligned_vs[0];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[3];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[2];

endmodule



module bsg_encode_one_hot_width_p16
(
  i,
  addr_o,
  v_o
);

  input [15:0] i;
  output [3:0] addr_o;
  output v_o;
  wire [3:0] addr_o;
  wire v_o;
  wire [5:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p8
  aligned_left
  (
    .i(i[7:0]),
    .addr_o(aligned_addrs[2:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p8
  aligned_right
  (
    .i(i[15:8]),
    .addr_o(aligned_addrs[5:3]),
    .v_o(addr_o[3])
  );

  assign v_o = addr_o[3] | aligned_vs[0];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[5];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[4];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[3];

endmodule



module bsg_encode_one_hot_width_p11
(
  i,
  addr_o,
  v_o
);

  input [10:0] i;
  output [3:0] addr_o;
  output v_o;
  wire [3:0] addr_o;
  wire v_o;

  bsg_encode_one_hot_width_p16
  unaligned_align
  (
    .i({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, i }),
    .addr_o(addr_o),
    .v_o(v_o)
  );


endmodule



module bsg_thermometer_count_width_p10
(
  i,
  o
);

  input [9:0] i;
  output [3:0] o;
  wire [3:0] o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8;
  wire [9:0] big_one_hot;

  bsg_encode_one_hot_width_p11
  big_encode_one_hot
  (
    .i({ i[9:9], big_one_hot }),
    .addr_o(o)
  );

  assign big_one_hot[9] = N0 & i[8];
  assign N0 = ~i[9];
  assign big_one_hot[8] = N1 & i[7];
  assign N1 = ~i[8];
  assign big_one_hot[7] = N2 & i[6];
  assign N2 = ~i[7];
  assign big_one_hot[6] = N3 & i[5];
  assign N3 = ~i[6];
  assign big_one_hot[5] = N4 & i[4];
  assign N4 = ~i[5];
  assign big_one_hot[4] = N5 & i[3];
  assign N5 = ~i[4];
  assign big_one_hot[3] = N6 & i[2];
  assign N6 = ~i[3];
  assign big_one_hot[2] = N7 & i[1];
  assign N7 = ~i[2];
  assign big_one_hot[1] = N8 & i[0];
  assign N8 = ~i[1];
  assign big_one_hot[0] = ~i[0];

endmodule



module bsg_rr_f2f_middle_width_p64_middle_meet_p10
(
  valid_head_i,
  ready_head_i,
  go_channels_o,
  go_cnt_o
);

  input [9:0] valid_head_i;
  input [9:0] ready_head_i;
  output [9:0] go_channels_o;
  output [3:0] go_cnt_o;
  wire [9:0] go_channels_o,happy_channels;
  wire [3:0] go_cnt_o;

  bsg_scan_width_p10_and_p1_lo_to_hi_p1
  and_scan
  (
    .i(happy_channels),
    .o(go_channels_o)
  );


  bsg_thermometer_count_width_p10
  genblk1_genblk1_thermo
  (
    .i(go_channels_o),
    .o(go_cnt_o)
  );

  assign happy_channels[9] = valid_head_i[9] & ready_head_i[9];
  assign happy_channels[8] = valid_head_i[8] & ready_head_i[8];
  assign happy_channels[7] = valid_head_i[7] & ready_head_i[7];
  assign happy_channels[6] = valid_head_i[6] & ready_head_i[6];
  assign happy_channels[5] = valid_head_i[5] & ready_head_i[5];
  assign happy_channels[4] = valid_head_i[4] & ready_head_i[4];
  assign happy_channels[3] = valid_head_i[3] & ready_head_i[3];
  assign happy_channels[2] = valid_head_i[2] & ready_head_i[2];
  assign happy_channels[1] = valid_head_i[1] & ready_head_i[1];
  assign happy_channels[0] = valid_head_i[0] & ready_head_i[0];

endmodule



module bsg_rr_f2f_output_width_p64_num_out_p10_middle_meet_p10
(
  clk,
  reset,
  ready_i,
  ready_head_o,
  go_channels_i,
  go_cnt_i,
  data_head_i,
  valid_o,
  data_o
);

  input [9:0] ready_i;
  output [9:0] ready_head_o;
  input [9:0] go_channels_i;
  input [3:0] go_cnt_i;
  input [639:0] data_head_i;
  output [9:0] valid_o;
  output [639:0] data_o;
  input clk;
  input reset;
  wire [9:0] ready_head_o,valid_o;
  wire [639:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,SYNOPSYS_UNCONNECTED_1,
  SYNOPSYS_UNCONNECTED_2,SYNOPSYS_UNCONNECTED_3,SYNOPSYS_UNCONNECTED_4,
  SYNOPSYS_UNCONNECTED_5,SYNOPSYS_UNCONNECTED_6,SYNOPSYS_UNCONNECTED_7,SYNOPSYS_UNCONNECTED_8,
  SYNOPSYS_UNCONNECTED_9,SYNOPSYS_UNCONNECTED_10,SYNOPSYS_UNCONNECTED_11,
  SYNOPSYS_UNCONNECTED_12,SYNOPSYS_UNCONNECTED_13,SYNOPSYS_UNCONNECTED_14,
  SYNOPSYS_UNCONNECTED_15,SYNOPSYS_UNCONNECTED_16,SYNOPSYS_UNCONNECTED_17,SYNOPSYS_UNCONNECTED_18;
  wire [3:0] optr_r,optr_r_data;

  bsg_rotate_right_width_p10
  ready_rr
  (
    .data_i(ready_i),
    .rot_i(optr_r),
    .o(ready_head_o)
  );

  assign { valid_o, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10 } = { go_channels_i, go_channels_i } << optr_r;

  bsg_circular_ptr_slots_p10_max_add_p10
  c_ptr
  (
    .clk(clk),
    .reset_i(reset),
    .add_i(go_cnt_i),
    .o(optr_r),
    .n_o({ SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14 })
  );


  bsg_circular_ptr_slots_p10_max_add_p10
  c_ptr_data
  (
    .clk(clk),
    .reset_i(reset),
    .add_i(go_cnt_i),
    .o(optr_r_data),
    .n_o({ SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18 })
  );

  assign N370 = N0 & optr_r_data[3];
  assign N0 = ~optr_r_data[2];
  assign N371 = optr_r_data[2] & N1;
  assign N1 = ~optr_r_data[3];
  assign N372 = N2 & N3;
  assign N2 = ~optr_r_data[2];
  assign N3 = ~optr_r_data[3];
  assign N373 = optr_r_data[0] & optr_r_data[1];
  assign N374 = N4 & optr_r_data[1];
  assign N4 = ~optr_r_data[0];
  assign N375 = optr_r_data[0] & N5;
  assign N5 = ~optr_r_data[1];
  assign N376 = N6 & N7;
  assign N6 = ~optr_r_data[0];
  assign N7 = ~optr_r_data[1];
  assign N235 = N370 & N374;
  assign N234 = N370 & N375;
  assign N233 = N370 & N376;
  assign N232 = N371 & N373;
  assign N231 = N371 & N374;
  assign N230 = N371 & N375;
  assign N229 = N371 & N376;
  assign N228 = N372 & N373;
  assign N227 = N372 & N374;
  assign N226 = N372 & N375;
  assign N225 = N372 & N376;
  assign N377 = N8 & optr_r_data[3];
  assign N8 = ~optr_r_data[2];
  assign N378 = optr_r_data[2] & N9;
  assign N9 = ~optr_r_data[3];
  assign N379 = N10 & N11;
  assign N10 = ~optr_r_data[2];
  assign N11 = ~optr_r_data[3];
  assign N380 = optr_r_data[0] & optr_r_data[1];
  assign N381 = N12 & optr_r_data[1];
  assign N12 = ~optr_r_data[0];
  assign N382 = optr_r_data[0] & N13;
  assign N13 = ~optr_r_data[1];
  assign N383 = N14 & N15;
  assign N14 = ~optr_r_data[0];
  assign N15 = ~optr_r_data[1];
  assign N247 = N377 & N380;
  assign N246 = N377 & N381;
  assign N245 = N377 & N382;
  assign N244 = N377 & N383;
  assign N243 = N378 & N380;
  assign N242 = N378 & N381;
  assign N241 = N378 & N382;
  assign N240 = N378 & N383;
  assign N239 = N379 & N380;
  assign N238 = N379 & N381;
  assign N237 = N379 & N382;
  assign N236 = N379 & N383;
  assign N384 = optr_r_data[2] & optr_r_data[3];
  assign N385 = N16 & optr_r_data[3];
  assign N16 = ~optr_r_data[2];
  assign N386 = optr_r_data[2] & N17;
  assign N17 = ~optr_r_data[3];
  assign N387 = N18 & N19;
  assign N18 = ~optr_r_data[2];
  assign N19 = ~optr_r_data[3];
  assign N388 = optr_r_data[0] & optr_r_data[1];
  assign N389 = N20 & optr_r_data[1];
  assign N20 = ~optr_r_data[0];
  assign N390 = optr_r_data[0] & N21;
  assign N21 = ~optr_r_data[1];
  assign N391 = N22 & N23;
  assign N22 = ~optr_r_data[0];
  assign N23 = ~optr_r_data[1];
  assign N260 = N384 & N391;
  assign N259 = N385 & N388;
  assign N258 = N385 & N389;
  assign N257 = N385 & N390;
  assign N256 = N385 & N391;
  assign N255 = N386 & N388;
  assign N254 = N386 & N389;
  assign N253 = N386 & N390;
  assign N252 = N386 & N391;
  assign N251 = N387 & N388;
  assign N250 = N387 & N389;
  assign N249 = N387 & N390;
  assign N248 = N387 & N391;
  assign N392 = optr_r_data[2] & optr_r_data[3];
  assign N393 = N24 & optr_r_data[3];
  assign N24 = ~optr_r_data[2];
  assign N394 = optr_r_data[2] & N25;
  assign N25 = ~optr_r_data[3];
  assign N395 = N26 & N27;
  assign N26 = ~optr_r_data[2];
  assign N27 = ~optr_r_data[3];
  assign N396 = optr_r_data[0] & optr_r_data[1];
  assign N397 = N28 & optr_r_data[1];
  assign N28 = ~optr_r_data[0];
  assign N398 = optr_r_data[0] & N29;
  assign N29 = ~optr_r_data[1];
  assign N399 = N30 & N31;
  assign N30 = ~optr_r_data[0];
  assign N31 = ~optr_r_data[1];
  assign N274 = N392 & N398;
  assign N273 = N392 & N399;
  assign N272 = N393 & N396;
  assign N271 = N393 & N397;
  assign N270 = N393 & N398;
  assign N269 = N393 & N399;
  assign N268 = N394 & N396;
  assign N267 = N394 & N397;
  assign N266 = N394 & N398;
  assign N265 = N394 & N399;
  assign N264 = N395 & N396;
  assign N263 = N395 & N397;
  assign N262 = N395 & N398;
  assign N261 = N395 & N399;
  assign N400 = optr_r_data[2] & optr_r_data[3];
  assign N401 = N32 & optr_r_data[3];
  assign N32 = ~optr_r_data[2];
  assign N402 = optr_r_data[2] & N33;
  assign N33 = ~optr_r_data[3];
  assign N403 = N34 & N35;
  assign N34 = ~optr_r_data[2];
  assign N35 = ~optr_r_data[3];
  assign N404 = optr_r_data[0] & optr_r_data[1];
  assign N405 = N36 & optr_r_data[1];
  assign N36 = ~optr_r_data[0];
  assign N406 = optr_r_data[0] & N37;
  assign N37 = ~optr_r_data[1];
  assign N407 = N38 & N39;
  assign N38 = ~optr_r_data[0];
  assign N39 = ~optr_r_data[1];
  assign N289 = N400 & N405;
  assign N288 = N400 & N406;
  assign N287 = N400 & N407;
  assign N286 = N401 & N404;
  assign N285 = N401 & N405;
  assign N284 = N401 & N406;
  assign N283 = N401 & N407;
  assign N282 = N402 & N404;
  assign N281 = N402 & N405;
  assign N280 = N402 & N406;
  assign N279 = N402 & N407;
  assign N278 = N403 & N404;
  assign N277 = N403 & N405;
  assign N276 = N403 & N406;
  assign N275 = N403 & N407;
  assign N408 = optr_r_data[2] & optr_r_data[3];
  assign N409 = N40 & optr_r_data[3];
  assign N40 = ~optr_r_data[2];
  assign N410 = optr_r_data[2] & N41;
  assign N41 = ~optr_r_data[3];
  assign N411 = N42 & N43;
  assign N42 = ~optr_r_data[2];
  assign N43 = ~optr_r_data[3];
  assign N412 = optr_r_data[0] & optr_r_data[1];
  assign N413 = N44 & optr_r_data[1];
  assign N44 = ~optr_r_data[0];
  assign N414 = optr_r_data[0] & N45;
  assign N45 = ~optr_r_data[1];
  assign N415 = N46 & N47;
  assign N46 = ~optr_r_data[0];
  assign N47 = ~optr_r_data[1];
  assign N305 = N408 & N412;
  assign N304 = N408 & N413;
  assign N303 = N408 & N414;
  assign N302 = N408 & N415;
  assign N301 = N409 & N412;
  assign N300 = N409 & N413;
  assign N299 = N409 & N414;
  assign N298 = N409 & N415;
  assign N297 = N410 & N412;
  assign N296 = N410 & N413;
  assign N295 = N410 & N414;
  assign N294 = N410 & N415;
  assign N293 = N411 & N412;
  assign N292 = N411 & N413;
  assign N291 = N411 & N414;
  assign N290 = N411 & N415;
  assign N416 = optr_r_data[2] & optr_r_data[3];
  assign N417 = N48 & optr_r_data[3];
  assign N48 = ~optr_r_data[2];
  assign N418 = optr_r_data[2] & N49;
  assign N49 = ~optr_r_data[3];
  assign N419 = N50 & N51;
  assign N50 = ~optr_r_data[2];
  assign N51 = ~optr_r_data[3];
  assign N420 = optr_r_data[0] & optr_r_data[1];
  assign N421 = N52 & optr_r_data[1];
  assign N52 = ~optr_r_data[0];
  assign N422 = optr_r_data[0] & N53;
  assign N53 = ~optr_r_data[1];
  assign N423 = N54 & N55;
  assign N54 = ~optr_r_data[0];
  assign N55 = ~optr_r_data[1];
  assign N321 = N416 & N420;
  assign N320 = N416 & N421;
  assign N319 = N416 & N422;
  assign N318 = N416 & N423;
  assign N317 = N417 & N420;
  assign N316 = N417 & N421;
  assign N315 = N417 & N422;
  assign N314 = N417 & N423;
  assign N313 = N418 & N420;
  assign N312 = N418 & N421;
  assign N311 = N418 & N422;
  assign N310 = N418 & N423;
  assign N309 = N419 & N420;
  assign N308 = N419 & N421;
  assign N307 = N419 & N422;
  assign N306 = N419 & N423;
  assign N424 = optr_r_data[2] & optr_r_data[3];
  assign N425 = N56 & optr_r_data[3];
  assign N56 = ~optr_r_data[2];
  assign N426 = optr_r_data[2] & N57;
  assign N57 = ~optr_r_data[3];
  assign N427 = N58 & N59;
  assign N58 = ~optr_r_data[2];
  assign N59 = ~optr_r_data[3];
  assign N428 = optr_r_data[0] & optr_r_data[1];
  assign N429 = N60 & optr_r_data[1];
  assign N60 = ~optr_r_data[0];
  assign N430 = optr_r_data[0] & N61;
  assign N61 = ~optr_r_data[1];
  assign N431 = N62 & N63;
  assign N62 = ~optr_r_data[0];
  assign N63 = ~optr_r_data[1];
  assign N337 = N424 & N428;
  assign N336 = N424 & N429;
  assign N335 = N424 & N430;
  assign N334 = N424 & N431;
  assign N333 = N425 & N428;
  assign N332 = N425 & N429;
  assign N331 = N425 & N430;
  assign N330 = N425 & N431;
  assign N329 = N426 & N428;
  assign N328 = N426 & N429;
  assign N327 = N426 & N430;
  assign N326 = N426 & N431;
  assign N325 = N427 & N428;
  assign N324 = N427 & N429;
  assign N323 = N427 & N430;
  assign N322 = N427 & N431;
  assign N432 = optr_r_data[2] & optr_r_data[3];
  assign N433 = N64 & optr_r_data[3];
  assign N64 = ~optr_r_data[2];
  assign N434 = optr_r_data[2] & N65;
  assign N65 = ~optr_r_data[3];
  assign N435 = N66 & N67;
  assign N66 = ~optr_r_data[2];
  assign N67 = ~optr_r_data[3];
  assign N436 = optr_r_data[0] & optr_r_data[1];
  assign N437 = N68 & optr_r_data[1];
  assign N68 = ~optr_r_data[0];
  assign N438 = optr_r_data[0] & N69;
  assign N69 = ~optr_r_data[1];
  assign N439 = N70 & N71;
  assign N70 = ~optr_r_data[0];
  assign N71 = ~optr_r_data[1];
  assign N353 = N432 & N436;
  assign N352 = N432 & N437;
  assign N351 = N432 & N438;
  assign N350 = N432 & N439;
  assign N349 = N433 & N436;
  assign N348 = N433 & N437;
  assign N347 = N433 & N438;
  assign N346 = N433 & N439;
  assign N345 = N434 & N436;
  assign N344 = N434 & N437;
  assign N343 = N434 & N438;
  assign N342 = N434 & N439;
  assign N341 = N435 & N436;
  assign N340 = N435 & N437;
  assign N339 = N435 & N438;
  assign N338 = N435 & N439;
  assign N440 = optr_r_data[2] & optr_r_data[3];
  assign N441 = N72 & optr_r_data[3];
  assign N72 = ~optr_r_data[2];
  assign N442 = optr_r_data[2] & N73;
  assign N73 = ~optr_r_data[3];
  assign N443 = N74 & N75;
  assign N74 = ~optr_r_data[2];
  assign N75 = ~optr_r_data[3];
  assign N444 = optr_r_data[0] & optr_r_data[1];
  assign N445 = N76 & optr_r_data[1];
  assign N76 = ~optr_r_data[0];
  assign N446 = optr_r_data[0] & N77;
  assign N77 = ~optr_r_data[1];
  assign N447 = N78 & N79;
  assign N78 = ~optr_r_data[0];
  assign N79 = ~optr_r_data[1];
  assign N369 = N440 & N444;
  assign N368 = N440 & N445;
  assign N367 = N440 & N446;
  assign N366 = N440 & N447;
  assign N365 = N441 & N444;
  assign N364 = N441 & N445;
  assign N363 = N441 & N446;
  assign N362 = N441 & N447;
  assign N361 = N442 & N444;
  assign N360 = N442 & N445;
  assign N359 = N442 & N446;
  assign N358 = N442 & N447;
  assign N357 = N443 & N444;
  assign N356 = N443 & N445;
  assign N355 = N443 & N446;
  assign N354 = N443 & N447;
  assign data_o[63:0] = (N80)? data_head_i[63:0] : 
                        (N81)? data_head_i[127:64] : 
                        (N82)? data_head_i[191:128] : 
                        (N83)? data_head_i[255:192] : 
                        (N84)? data_head_i[319:256] : 
                        (N85)? data_head_i[383:320] : 
                        (N86)? data_head_i[447:384] : 
                        (N87)? data_head_i[511:448] : 
                        (N88)? data_head_i[575:512] : 
                        (N89)? data_head_i[639:576] : 
                        (N90)? data_head_i[63:0] : 1'b0;
  assign N80 = N235;
  assign N81 = N234;
  assign N82 = N233;
  assign N83 = N232;
  assign N84 = N231;
  assign N85 = N230;
  assign N86 = N229;
  assign N87 = N228;
  assign N88 = N227;
  assign N89 = N226;
  assign N90 = N225;
  assign data_o[127:64] = (N91)? data_head_i[63:0] : 
                          (N92)? data_head_i[127:64] : 
                          (N93)? data_head_i[191:128] : 
                          (N94)? data_head_i[255:192] : 
                          (N95)? data_head_i[319:256] : 
                          (N96)? data_head_i[383:320] : 
                          (N97)? data_head_i[447:384] : 
                          (N98)? data_head_i[511:448] : 
                          (N99)? data_head_i[575:512] : 
                          (N100)? data_head_i[639:576] : 
                          (N101)? data_head_i[63:0] : 
                          (N102)? data_head_i[127:64] : 1'b0;
  assign N91 = N247;
  assign N92 = N246;
  assign N93 = N245;
  assign N94 = N244;
  assign N95 = N243;
  assign N96 = N242;
  assign N97 = N241;
  assign N98 = N240;
  assign N99 = N239;
  assign N100 = N238;
  assign N101 = N237;
  assign N102 = N236;
  assign data_o[191:128] = (N103)? data_head_i[63:0] : 
                           (N104)? data_head_i[127:64] : 
                           (N105)? data_head_i[191:128] : 
                           (N106)? data_head_i[255:192] : 
                           (N107)? data_head_i[319:256] : 
                           (N108)? data_head_i[383:320] : 
                           (N109)? data_head_i[447:384] : 
                           (N110)? data_head_i[511:448] : 
                           (N111)? data_head_i[575:512] : 
                           (N112)? data_head_i[639:576] : 
                           (N113)? data_head_i[63:0] : 
                           (N114)? data_head_i[127:64] : 
                           (N115)? data_head_i[191:128] : 1'b0;
  assign N103 = N260;
  assign N104 = N259;
  assign N105 = N258;
  assign N106 = N257;
  assign N107 = N256;
  assign N108 = N255;
  assign N109 = N254;
  assign N110 = N253;
  assign N111 = N252;
  assign N112 = N251;
  assign N113 = N250;
  assign N114 = N249;
  assign N115 = N248;
  assign data_o[255:192] = (N116)? data_head_i[63:0] : 
                           (N117)? data_head_i[127:64] : 
                           (N118)? data_head_i[191:128] : 
                           (N119)? data_head_i[255:192] : 
                           (N120)? data_head_i[319:256] : 
                           (N121)? data_head_i[383:320] : 
                           (N122)? data_head_i[447:384] : 
                           (N123)? data_head_i[511:448] : 
                           (N124)? data_head_i[575:512] : 
                           (N125)? data_head_i[639:576] : 
                           (N126)? data_head_i[63:0] : 
                           (N127)? data_head_i[127:64] : 
                           (N128)? data_head_i[191:128] : 
                           (N129)? data_head_i[255:192] : 1'b0;
  assign N116 = N274;
  assign N117 = N273;
  assign N118 = N272;
  assign N119 = N271;
  assign N120 = N270;
  assign N121 = N269;
  assign N122 = N268;
  assign N123 = N267;
  assign N124 = N266;
  assign N125 = N265;
  assign N126 = N264;
  assign N127 = N263;
  assign N128 = N262;
  assign N129 = N261;
  assign data_o[319:256] = (N130)? data_head_i[63:0] : 
                           (N131)? data_head_i[127:64] : 
                           (N132)? data_head_i[191:128] : 
                           (N133)? data_head_i[255:192] : 
                           (N134)? data_head_i[319:256] : 
                           (N135)? data_head_i[383:320] : 
                           (N136)? data_head_i[447:384] : 
                           (N137)? data_head_i[511:448] : 
                           (N138)? data_head_i[575:512] : 
                           (N139)? data_head_i[639:576] : 
                           (N140)? data_head_i[63:0] : 
                           (N141)? data_head_i[127:64] : 
                           (N142)? data_head_i[191:128] : 
                           (N143)? data_head_i[255:192] : 
                           (N144)? data_head_i[319:256] : 1'b0;
  assign N130 = N289;
  assign N131 = N288;
  assign N132 = N287;
  assign N133 = N286;
  assign N134 = N285;
  assign N135 = N284;
  assign N136 = N283;
  assign N137 = N282;
  assign N138 = N281;
  assign N139 = N280;
  assign N140 = N279;
  assign N141 = N278;
  assign N142 = N277;
  assign N143 = N276;
  assign N144 = N275;
  assign data_o[383:320] = (N145)? data_head_i[63:0] : 
                           (N146)? data_head_i[127:64] : 
                           (N147)? data_head_i[191:128] : 
                           (N148)? data_head_i[255:192] : 
                           (N149)? data_head_i[319:256] : 
                           (N150)? data_head_i[383:320] : 
                           (N151)? data_head_i[447:384] : 
                           (N152)? data_head_i[511:448] : 
                           (N153)? data_head_i[575:512] : 
                           (N154)? data_head_i[639:576] : 
                           (N155)? data_head_i[63:0] : 
                           (N156)? data_head_i[127:64] : 
                           (N157)? data_head_i[191:128] : 
                           (N158)? data_head_i[255:192] : 
                           (N159)? data_head_i[319:256] : 
                           (N160)? data_head_i[383:320] : 1'b0;
  assign N145 = N305;
  assign N146 = N304;
  assign N147 = N303;
  assign N148 = N302;
  assign N149 = N301;
  assign N150 = N300;
  assign N151 = N299;
  assign N152 = N298;
  assign N153 = N297;
  assign N154 = N296;
  assign N155 = N295;
  assign N156 = N294;
  assign N157 = N293;
  assign N158 = N292;
  assign N159 = N291;
  assign N160 = N290;
  assign data_o[447:384] = (N161)? data_head_i[127:64] : 
                           (N162)? data_head_i[191:128] : 
                           (N163)? data_head_i[255:192] : 
                           (N164)? data_head_i[319:256] : 
                           (N165)? data_head_i[383:320] : 
                           (N166)? data_head_i[447:384] : 
                           (N167)? data_head_i[511:448] : 
                           (N168)? data_head_i[575:512] : 
                           (N169)? data_head_i[639:576] : 
                           (N170)? data_head_i[63:0] : 
                           (N171)? data_head_i[127:64] : 
                           (N172)? data_head_i[191:128] : 
                           (N173)? data_head_i[255:192] : 
                           (N174)? data_head_i[319:256] : 
                           (N175)? data_head_i[383:320] : 
                           (N176)? data_head_i[447:384] : 1'b0;
  assign N161 = N321;
  assign N162 = N320;
  assign N163 = N319;
  assign N164 = N318;
  assign N165 = N317;
  assign N166 = N316;
  assign N167 = N315;
  assign N168 = N314;
  assign N169 = N313;
  assign N170 = N312;
  assign N171 = N311;
  assign N172 = N310;
  assign N173 = N309;
  assign N174 = N308;
  assign N175 = N307;
  assign N176 = N306;
  assign data_o[511:448] = (N177)? data_head_i[191:128] : 
                           (N178)? data_head_i[255:192] : 
                           (N179)? data_head_i[319:256] : 
                           (N180)? data_head_i[383:320] : 
                           (N181)? data_head_i[447:384] : 
                           (N182)? data_head_i[511:448] : 
                           (N183)? data_head_i[575:512] : 
                           (N184)? data_head_i[639:576] : 
                           (N185)? data_head_i[63:0] : 
                           (N186)? data_head_i[127:64] : 
                           (N187)? data_head_i[191:128] : 
                           (N188)? data_head_i[255:192] : 
                           (N189)? data_head_i[319:256] : 
                           (N190)? data_head_i[383:320] : 
                           (N191)? data_head_i[447:384] : 
                           (N192)? data_head_i[511:448] : 1'b0;
  assign N177 = N337;
  assign N178 = N336;
  assign N179 = N335;
  assign N180 = N334;
  assign N181 = N333;
  assign N182 = N332;
  assign N183 = N331;
  assign N184 = N330;
  assign N185 = N329;
  assign N186 = N328;
  assign N187 = N327;
  assign N188 = N326;
  assign N189 = N325;
  assign N190 = N324;
  assign N191 = N323;
  assign N192 = N322;
  assign data_o[575:512] = (N193)? data_head_i[255:192] : 
                           (N194)? data_head_i[319:256] : 
                           (N195)? data_head_i[383:320] : 
                           (N196)? data_head_i[447:384] : 
                           (N197)? data_head_i[511:448] : 
                           (N198)? data_head_i[575:512] : 
                           (N199)? data_head_i[639:576] : 
                           (N200)? data_head_i[63:0] : 
                           (N201)? data_head_i[127:64] : 
                           (N202)? data_head_i[191:128] : 
                           (N203)? data_head_i[255:192] : 
                           (N204)? data_head_i[319:256] : 
                           (N205)? data_head_i[383:320] : 
                           (N206)? data_head_i[447:384] : 
                           (N207)? data_head_i[511:448] : 
                           (N208)? data_head_i[575:512] : 1'b0;
  assign N193 = N353;
  assign N194 = N352;
  assign N195 = N351;
  assign N196 = N350;
  assign N197 = N349;
  assign N198 = N348;
  assign N199 = N347;
  assign N200 = N346;
  assign N201 = N345;
  assign N202 = N344;
  assign N203 = N343;
  assign N204 = N342;
  assign N205 = N341;
  assign N206 = N340;
  assign N207 = N339;
  assign N208 = N338;
  assign data_o[639:576] = (N209)? data_head_i[319:256] : 
                           (N210)? data_head_i[383:320] : 
                           (N211)? data_head_i[447:384] : 
                           (N212)? data_head_i[511:448] : 
                           (N213)? data_head_i[575:512] : 
                           (N214)? data_head_i[639:576] : 
                           (N215)? data_head_i[63:0] : 
                           (N216)? data_head_i[127:64] : 
                           (N217)? data_head_i[191:128] : 
                           (N218)? data_head_i[255:192] : 
                           (N219)? data_head_i[319:256] : 
                           (N220)? data_head_i[383:320] : 
                           (N221)? data_head_i[447:384] : 
                           (N222)? data_head_i[511:448] : 
                           (N223)? data_head_i[575:512] : 
                           (N224)? data_head_i[639:576] : 1'b0;
  assign N209 = N369;
  assign N210 = N368;
  assign N211 = N367;
  assign N212 = N366;
  assign N213 = N365;
  assign N214 = N364;
  assign N215 = N363;
  assign N216 = N362;
  assign N217 = N361;
  assign N218 = N360;
  assign N219 = N359;
  assign N220 = N358;
  assign N221 = N357;
  assign N222 = N356;
  assign N223 = N355;
  assign N224 = N354;

endmodule



module bsg_round_robin_fifo_to_fifo_width_p64_num_in_p10_num_out_p10_out_channel_count_mask_p512
(
  clk,
  reset,
  valid_i,
  data_i,
  yumi_o,
  in_top_channel_i,
  out_top_channel_i,
  valid_o,
  data_o,
  ready_i
);

  input [9:0] valid_i;
  input [639:0] data_i;
  output [9:0] yumi_o;
  input [3:0] in_top_channel_i;
  input [3:0] out_top_channel_i;
  output [9:0] valid_o;
  output [639:0] data_o;
  input [9:0] ready_i;
  input clk;
  input reset;
  wire [9:0] yumi_o,valid_o,go_channels;
  wire [639:0] data_o,data_o_flat,oc_9__out_chan_data_head_array;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,yumi_int_o_9__9_,yumi_int_o_9__8_,
  yumi_int_o_9__7_,yumi_int_o_9__6_,yumi_int_o_9__5_,yumi_int_o_9__4_,yumi_int_o_9__3_,
  yumi_int_o_9__2_,yumi_int_o_9__1_,yumi_int_o_9__0_,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,valid_int_o_9__9_,valid_int_o_9__8_,valid_int_o_9__7_,
  valid_int_o_9__6_,valid_int_o_9__5_,valid_int_o_9__4_,valid_int_o_9__3_,valid_int_o_9__2_,
  valid_int_o_9__1_,valid_int_o_9__0_,N135,N136,N137,N138,N139,N140,N141,N142,N143,
  N144,data_int_o_9__639_,data_int_o_9__638_,data_int_o_9__637_,
  data_int_o_9__636_,data_int_o_9__635_,data_int_o_9__634_,data_int_o_9__633_,data_int_o_9__632_,
  data_int_o_9__631_,data_int_o_9__630_,data_int_o_9__629_,data_int_o_9__628_,
  data_int_o_9__627_,data_int_o_9__626_,data_int_o_9__625_,data_int_o_9__624_,
  data_int_o_9__623_,data_int_o_9__622_,data_int_o_9__621_,data_int_o_9__620_,
  data_int_o_9__619_,data_int_o_9__618_,data_int_o_9__617_,data_int_o_9__616_,data_int_o_9__615_,
  data_int_o_9__614_,data_int_o_9__613_,data_int_o_9__612_,data_int_o_9__611_,
  data_int_o_9__610_,data_int_o_9__609_,data_int_o_9__608_,data_int_o_9__607_,
  data_int_o_9__606_,data_int_o_9__605_,data_int_o_9__604_,data_int_o_9__603_,
  data_int_o_9__602_,data_int_o_9__601_,data_int_o_9__600_,data_int_o_9__599_,
  data_int_o_9__598_,data_int_o_9__597_,data_int_o_9__596_,data_int_o_9__595_,data_int_o_9__594_,
  data_int_o_9__593_,data_int_o_9__592_,data_int_o_9__591_,data_int_o_9__590_,
  data_int_o_9__589_,data_int_o_9__588_,data_int_o_9__587_,data_int_o_9__586_,
  data_int_o_9__585_,data_int_o_9__584_,data_int_o_9__583_,data_int_o_9__582_,
  data_int_o_9__581_,data_int_o_9__580_,data_int_o_9__579_,data_int_o_9__578_,
  data_int_o_9__577_,data_int_o_9__576_,data_int_o_9__575_,data_int_o_9__574_,data_int_o_9__573_,
  data_int_o_9__572_,data_int_o_9__571_,data_int_o_9__570_,data_int_o_9__569_,
  data_int_o_9__568_,data_int_o_9__567_,data_int_o_9__566_,data_int_o_9__565_,
  data_int_o_9__564_,data_int_o_9__563_,data_int_o_9__562_,data_int_o_9__561_,
  data_int_o_9__560_,data_int_o_9__559_,data_int_o_9__558_,data_int_o_9__557_,
  data_int_o_9__556_,data_int_o_9__555_,data_int_o_9__554_,data_int_o_9__553_,data_int_o_9__552_,
  data_int_o_9__551_,data_int_o_9__550_,data_int_o_9__549_,data_int_o_9__548_,
  data_int_o_9__547_,data_int_o_9__546_,data_int_o_9__545_,data_int_o_9__544_,
  data_int_o_9__543_,data_int_o_9__542_,data_int_o_9__541_,data_int_o_9__540_,
  data_int_o_9__539_,data_int_o_9__538_,data_int_o_9__537_,data_int_o_9__536_,data_int_o_9__535_,
  data_int_o_9__534_,data_int_o_9__533_,data_int_o_9__532_,data_int_o_9__531_,
  data_int_o_9__530_,data_int_o_9__529_,data_int_o_9__528_,data_int_o_9__527_,
  data_int_o_9__526_,data_int_o_9__525_,data_int_o_9__524_,data_int_o_9__523_,
  data_int_o_9__522_,data_int_o_9__521_,data_int_o_9__520_,data_int_o_9__519_,
  data_int_o_9__518_,data_int_o_9__517_,data_int_o_9__516_,data_int_o_9__515_,data_int_o_9__514_,
  data_int_o_9__513_,data_int_o_9__512_,data_int_o_9__511_,data_int_o_9__510_,
  data_int_o_9__509_,data_int_o_9__508_,data_int_o_9__507_,data_int_o_9__506_,
  data_int_o_9__505_,data_int_o_9__504_,data_int_o_9__503_,data_int_o_9__502_,
  data_int_o_9__501_,data_int_o_9__500_,data_int_o_9__499_,data_int_o_9__498_,
  data_int_o_9__497_,data_int_o_9__496_,data_int_o_9__495_,data_int_o_9__494_,data_int_o_9__493_,
  data_int_o_9__492_,data_int_o_9__491_,data_int_o_9__490_,data_int_o_9__489_,
  data_int_o_9__488_,data_int_o_9__487_,data_int_o_9__486_,data_int_o_9__485_,
  data_int_o_9__484_,data_int_o_9__483_,data_int_o_9__482_,data_int_o_9__481_,
  data_int_o_9__480_,data_int_o_9__479_,data_int_o_9__478_,data_int_o_9__477_,
  data_int_o_9__476_,data_int_o_9__475_,data_int_o_9__474_,data_int_o_9__473_,data_int_o_9__472_,
  data_int_o_9__471_,data_int_o_9__470_,data_int_o_9__469_,data_int_o_9__468_,
  data_int_o_9__467_,data_int_o_9__466_,data_int_o_9__465_,data_int_o_9__464_,
  data_int_o_9__463_,data_int_o_9__462_,data_int_o_9__461_,data_int_o_9__460_,
  data_int_o_9__459_,data_int_o_9__458_,data_int_o_9__457_,data_int_o_9__456_,data_int_o_9__455_,
  data_int_o_9__454_,data_int_o_9__453_,data_int_o_9__452_,data_int_o_9__451_,
  data_int_o_9__450_,data_int_o_9__449_,data_int_o_9__448_,data_int_o_9__447_,
  data_int_o_9__446_,data_int_o_9__445_,data_int_o_9__444_,data_int_o_9__443_,
  data_int_o_9__442_,data_int_o_9__441_,data_int_o_9__440_,data_int_o_9__439_,
  data_int_o_9__438_,data_int_o_9__437_,data_int_o_9__436_,data_int_o_9__435_,data_int_o_9__434_,
  data_int_o_9__433_,data_int_o_9__432_,data_int_o_9__431_,data_int_o_9__430_,
  data_int_o_9__429_,data_int_o_9__428_,data_int_o_9__427_,data_int_o_9__426_,
  data_int_o_9__425_,data_int_o_9__424_,data_int_o_9__423_,data_int_o_9__422_,
  data_int_o_9__421_,data_int_o_9__420_,data_int_o_9__419_,data_int_o_9__418_,
  data_int_o_9__417_,data_int_o_9__416_,data_int_o_9__415_,data_int_o_9__414_,data_int_o_9__413_,
  data_int_o_9__412_,data_int_o_9__411_,data_int_o_9__410_,data_int_o_9__409_,
  data_int_o_9__408_,data_int_o_9__407_,data_int_o_9__406_,data_int_o_9__405_,
  data_int_o_9__404_,data_int_o_9__403_,data_int_o_9__402_,data_int_o_9__401_,
  data_int_o_9__400_,data_int_o_9__399_,data_int_o_9__398_,data_int_o_9__397_,
  data_int_o_9__396_,data_int_o_9__395_,data_int_o_9__394_,data_int_o_9__393_,data_int_o_9__392_,
  data_int_o_9__391_,data_int_o_9__390_,data_int_o_9__389_,data_int_o_9__388_,
  data_int_o_9__387_,data_int_o_9__386_,data_int_o_9__385_,data_int_o_9__384_,
  data_int_o_9__383_,data_int_o_9__382_,data_int_o_9__381_,data_int_o_9__380_,
  data_int_o_9__379_,data_int_o_9__378_,data_int_o_9__377_,data_int_o_9__376_,data_int_o_9__375_,
  data_int_o_9__374_,data_int_o_9__373_,data_int_o_9__372_,data_int_o_9__371_,
  data_int_o_9__370_,data_int_o_9__369_,data_int_o_9__368_,data_int_o_9__367_,
  data_int_o_9__366_,data_int_o_9__365_,data_int_o_9__364_,data_int_o_9__363_,
  data_int_o_9__362_,data_int_o_9__361_,data_int_o_9__360_,data_int_o_9__359_,
  data_int_o_9__358_,data_int_o_9__357_,data_int_o_9__356_,data_int_o_9__355_,data_int_o_9__354_,
  data_int_o_9__353_,data_int_o_9__352_,data_int_o_9__351_,data_int_o_9__350_,
  data_int_o_9__349_,data_int_o_9__348_,data_int_o_9__347_,data_int_o_9__346_,
  data_int_o_9__345_,data_int_o_9__344_,data_int_o_9__343_,data_int_o_9__342_,
  data_int_o_9__341_,data_int_o_9__340_,data_int_o_9__339_,data_int_o_9__338_,
  data_int_o_9__337_,data_int_o_9__336_,data_int_o_9__335_,data_int_o_9__334_,data_int_o_9__333_,
  data_int_o_9__332_,data_int_o_9__331_,data_int_o_9__330_,data_int_o_9__329_,
  data_int_o_9__328_,data_int_o_9__327_,data_int_o_9__326_,data_int_o_9__325_,
  data_int_o_9__324_,data_int_o_9__323_,data_int_o_9__322_,data_int_o_9__321_,
  data_int_o_9__320_,data_int_o_9__319_,data_int_o_9__318_,data_int_o_9__317_,
  data_int_o_9__316_,data_int_o_9__315_,data_int_o_9__314_,data_int_o_9__313_,data_int_o_9__312_,
  data_int_o_9__311_,data_int_o_9__310_,data_int_o_9__309_,data_int_o_9__308_,
  data_int_o_9__307_,data_int_o_9__306_,data_int_o_9__305_,data_int_o_9__304_,
  data_int_o_9__303_,data_int_o_9__302_,data_int_o_9__301_,data_int_o_9__300_,
  data_int_o_9__299_,data_int_o_9__298_,data_int_o_9__297_,data_int_o_9__296_,data_int_o_9__295_,
  data_int_o_9__294_,data_int_o_9__293_,data_int_o_9__292_,data_int_o_9__291_,
  data_int_o_9__290_,data_int_o_9__289_,data_int_o_9__288_,data_int_o_9__287_,
  data_int_o_9__286_,data_int_o_9__285_,data_int_o_9__284_,data_int_o_9__283_,
  data_int_o_9__282_,data_int_o_9__281_,data_int_o_9__280_,data_int_o_9__279_,
  data_int_o_9__278_,data_int_o_9__277_,data_int_o_9__276_,data_int_o_9__275_,data_int_o_9__274_,
  data_int_o_9__273_,data_int_o_9__272_,data_int_o_9__271_,data_int_o_9__270_,
  data_int_o_9__269_,data_int_o_9__268_,data_int_o_9__267_,data_int_o_9__266_,
  data_int_o_9__265_,data_int_o_9__264_,data_int_o_9__263_,data_int_o_9__262_,
  data_int_o_9__261_,data_int_o_9__260_,data_int_o_9__259_,data_int_o_9__258_,
  data_int_o_9__257_,data_int_o_9__256_,data_int_o_9__255_,data_int_o_9__254_,data_int_o_9__253_,
  data_int_o_9__252_,data_int_o_9__251_,data_int_o_9__250_,data_int_o_9__249_,
  data_int_o_9__248_,data_int_o_9__247_,data_int_o_9__246_,data_int_o_9__245_,
  data_int_o_9__244_,data_int_o_9__243_,data_int_o_9__242_,data_int_o_9__241_,
  data_int_o_9__240_,data_int_o_9__239_,data_int_o_9__238_,data_int_o_9__237_,
  data_int_o_9__236_,data_int_o_9__235_,data_int_o_9__234_,data_int_o_9__233_,data_int_o_9__232_,
  data_int_o_9__231_,data_int_o_9__230_,data_int_o_9__229_,data_int_o_9__228_,
  data_int_o_9__227_,data_int_o_9__226_,data_int_o_9__225_,data_int_o_9__224_,
  data_int_o_9__223_,data_int_o_9__222_,data_int_o_9__221_,data_int_o_9__220_,
  data_int_o_9__219_,data_int_o_9__218_,data_int_o_9__217_,data_int_o_9__216_,data_int_o_9__215_,
  data_int_o_9__214_,data_int_o_9__213_,data_int_o_9__212_,data_int_o_9__211_,
  data_int_o_9__210_,data_int_o_9__209_,data_int_o_9__208_,data_int_o_9__207_,
  data_int_o_9__206_,data_int_o_9__205_,data_int_o_9__204_,data_int_o_9__203_,
  data_int_o_9__202_,data_int_o_9__201_,data_int_o_9__200_,data_int_o_9__199_,
  data_int_o_9__198_,data_int_o_9__197_,data_int_o_9__196_,data_int_o_9__195_,data_int_o_9__194_,
  data_int_o_9__193_,data_int_o_9__192_,data_int_o_9__191_,data_int_o_9__190_,
  data_int_o_9__189_,data_int_o_9__188_,data_int_o_9__187_,data_int_o_9__186_,
  data_int_o_9__185_,data_int_o_9__184_,data_int_o_9__183_,data_int_o_9__182_,
  data_int_o_9__181_,data_int_o_9__180_,data_int_o_9__179_,data_int_o_9__178_,
  data_int_o_9__177_,data_int_o_9__176_,data_int_o_9__175_,data_int_o_9__174_,data_int_o_9__173_,
  data_int_o_9__172_,data_int_o_9__171_,data_int_o_9__170_,data_int_o_9__169_,
  data_int_o_9__168_,data_int_o_9__167_,data_int_o_9__166_,data_int_o_9__165_,
  data_int_o_9__164_,data_int_o_9__163_,data_int_o_9__162_,data_int_o_9__161_,
  data_int_o_9__160_,data_int_o_9__159_,data_int_o_9__158_,data_int_o_9__157_,
  data_int_o_9__156_,data_int_o_9__155_,data_int_o_9__154_,data_int_o_9__153_,data_int_o_9__152_,
  data_int_o_9__151_,data_int_o_9__150_,data_int_o_9__149_,data_int_o_9__148_,
  data_int_o_9__147_,data_int_o_9__146_,data_int_o_9__145_,data_int_o_9__144_,
  data_int_o_9__143_,data_int_o_9__142_,data_int_o_9__141_,data_int_o_9__140_,
  data_int_o_9__139_,data_int_o_9__138_,data_int_o_9__137_,data_int_o_9__136_,data_int_o_9__135_,
  data_int_o_9__134_,data_int_o_9__133_,data_int_o_9__132_,data_int_o_9__131_,
  data_int_o_9__130_,data_int_o_9__129_,data_int_o_9__128_,data_int_o_9__127_,
  data_int_o_9__126_,data_int_o_9__125_,data_int_o_9__124_,data_int_o_9__123_,
  data_int_o_9__122_,data_int_o_9__121_,data_int_o_9__120_,data_int_o_9__119_,
  data_int_o_9__118_,data_int_o_9__117_,data_int_o_9__116_,data_int_o_9__115_,data_int_o_9__114_,
  data_int_o_9__113_,data_int_o_9__112_,data_int_o_9__111_,data_int_o_9__110_,
  data_int_o_9__109_,data_int_o_9__108_,data_int_o_9__107_,data_int_o_9__106_,
  data_int_o_9__105_,data_int_o_9__104_,data_int_o_9__103_,data_int_o_9__102_,
  data_int_o_9__101_,data_int_o_9__100_,data_int_o_9__99_,data_int_o_9__98_,data_int_o_9__97_,
  data_int_o_9__96_,data_int_o_9__95_,data_int_o_9__94_,data_int_o_9__93_,
  data_int_o_9__92_,data_int_o_9__91_,data_int_o_9__90_,data_int_o_9__89_,
  data_int_o_9__88_,data_int_o_9__87_,data_int_o_9__86_,data_int_o_9__85_,data_int_o_9__84_,
  data_int_o_9__83_,data_int_o_9__82_,data_int_o_9__81_,data_int_o_9__80_,
  data_int_o_9__79_,data_int_o_9__78_,data_int_o_9__77_,data_int_o_9__76_,data_int_o_9__75_,
  data_int_o_9__74_,data_int_o_9__73_,data_int_o_9__72_,data_int_o_9__71_,
  data_int_o_9__70_,data_int_o_9__69_,data_int_o_9__68_,data_int_o_9__67_,data_int_o_9__66_,
  data_int_o_9__65_,data_int_o_9__64_,data_int_o_9__63_,data_int_o_9__62_,
  data_int_o_9__61_,data_int_o_9__60_,data_int_o_9__59_,data_int_o_9__58_,data_int_o_9__57_,
  data_int_o_9__56_,data_int_o_9__55_,data_int_o_9__54_,data_int_o_9__53_,
  data_int_o_9__52_,data_int_o_9__51_,data_int_o_9__50_,data_int_o_9__49_,
  data_int_o_9__48_,data_int_o_9__47_,data_int_o_9__46_,data_int_o_9__45_,data_int_o_9__44_,
  data_int_o_9__43_,data_int_o_9__42_,data_int_o_9__41_,data_int_o_9__40_,
  data_int_o_9__39_,data_int_o_9__38_,data_int_o_9__37_,data_int_o_9__36_,data_int_o_9__35_,
  data_int_o_9__34_,data_int_o_9__33_,data_int_o_9__32_,data_int_o_9__31_,
  data_int_o_9__30_,data_int_o_9__29_,data_int_o_9__28_,data_int_o_9__27_,data_int_o_9__26_,
  data_int_o_9__25_,data_int_o_9__24_,data_int_o_9__23_,data_int_o_9__22_,
  data_int_o_9__21_,data_int_o_9__20_,data_int_o_9__19_,data_int_o_9__18_,data_int_o_9__17_,
  data_int_o_9__16_,data_int_o_9__15_,data_int_o_9__14_,data_int_o_9__13_,
  data_int_o_9__12_,data_int_o_9__11_,data_int_o_9__10_,data_int_o_9__9_,data_int_o_9__8_,
  data_int_o_9__7_,data_int_o_9__6_,data_int_o_9__5_,data_int_o_9__4_,
  data_int_o_9__3_,data_int_o_9__2_,data_int_o_9__1_,data_int_o_9__0_,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,data_head_9__639_,data_head_9__638_,data_head_9__637_,
  data_head_9__636_,data_head_9__635_,data_head_9__634_,data_head_9__633_,
  data_head_9__632_,data_head_9__631_,data_head_9__630_,data_head_9__629_,
  data_head_9__628_,data_head_9__627_,data_head_9__626_,data_head_9__625_,data_head_9__624_,
  data_head_9__623_,data_head_9__622_,data_head_9__621_,data_head_9__620_,
  data_head_9__619_,data_head_9__618_,data_head_9__617_,data_head_9__616_,data_head_9__615_,
  data_head_9__614_,data_head_9__613_,data_head_9__612_,data_head_9__611_,
  data_head_9__610_,data_head_9__609_,data_head_9__608_,data_head_9__607_,data_head_9__606_,
  data_head_9__605_,data_head_9__604_,data_head_9__603_,data_head_9__602_,
  data_head_9__601_,data_head_9__600_,data_head_9__599_,data_head_9__598_,data_head_9__597_,
  data_head_9__596_,data_head_9__595_,data_head_9__594_,data_head_9__593_,
  data_head_9__592_,data_head_9__591_,data_head_9__590_,data_head_9__589_,
  data_head_9__588_,data_head_9__587_,data_head_9__586_,data_head_9__585_,data_head_9__584_,
  data_head_9__583_,data_head_9__582_,data_head_9__581_,data_head_9__580_,
  data_head_9__579_,data_head_9__578_,data_head_9__577_,data_head_9__576_,data_head_9__575_,
  data_head_9__574_,data_head_9__573_,data_head_9__572_,data_head_9__571_,
  data_head_9__570_,data_head_9__569_,data_head_9__568_,data_head_9__567_,data_head_9__566_,
  data_head_9__565_,data_head_9__564_,data_head_9__563_,data_head_9__562_,
  data_head_9__561_,data_head_9__560_,data_head_9__559_,data_head_9__558_,data_head_9__557_,
  data_head_9__556_,data_head_9__555_,data_head_9__554_,data_head_9__553_,
  data_head_9__552_,data_head_9__551_,data_head_9__550_,data_head_9__549_,
  data_head_9__548_,data_head_9__547_,data_head_9__546_,data_head_9__545_,data_head_9__544_,
  data_head_9__543_,data_head_9__542_,data_head_9__541_,data_head_9__540_,
  data_head_9__539_,data_head_9__538_,data_head_9__537_,data_head_9__536_,data_head_9__535_,
  data_head_9__534_,data_head_9__533_,data_head_9__532_,data_head_9__531_,
  data_head_9__530_,data_head_9__529_,data_head_9__528_,data_head_9__527_,data_head_9__526_,
  data_head_9__525_,data_head_9__524_,data_head_9__523_,data_head_9__522_,
  data_head_9__521_,data_head_9__520_,data_head_9__519_,data_head_9__518_,data_head_9__517_,
  data_head_9__516_,data_head_9__515_,data_head_9__514_,data_head_9__513_,
  data_head_9__512_,data_head_9__511_,data_head_9__510_,data_head_9__509_,
  data_head_9__508_,data_head_9__507_,data_head_9__506_,data_head_9__505_,data_head_9__504_,
  data_head_9__503_,data_head_9__502_,data_head_9__501_,data_head_9__500_,
  data_head_9__499_,data_head_9__498_,data_head_9__497_,data_head_9__496_,data_head_9__495_,
  data_head_9__494_,data_head_9__493_,data_head_9__492_,data_head_9__491_,
  data_head_9__490_,data_head_9__489_,data_head_9__488_,data_head_9__487_,data_head_9__486_,
  data_head_9__485_,data_head_9__484_,data_head_9__483_,data_head_9__482_,
  data_head_9__481_,data_head_9__480_,data_head_9__479_,data_head_9__478_,data_head_9__477_,
  data_head_9__476_,data_head_9__475_,data_head_9__474_,data_head_9__473_,
  data_head_9__472_,data_head_9__471_,data_head_9__470_,data_head_9__469_,
  data_head_9__468_,data_head_9__467_,data_head_9__466_,data_head_9__465_,data_head_9__464_,
  data_head_9__463_,data_head_9__462_,data_head_9__461_,data_head_9__460_,
  data_head_9__459_,data_head_9__458_,data_head_9__457_,data_head_9__456_,data_head_9__455_,
  data_head_9__454_,data_head_9__453_,data_head_9__452_,data_head_9__451_,
  data_head_9__450_,data_head_9__449_,data_head_9__448_,data_head_9__447_,data_head_9__446_,
  data_head_9__445_,data_head_9__444_,data_head_9__443_,data_head_9__442_,
  data_head_9__441_,data_head_9__440_,data_head_9__439_,data_head_9__438_,data_head_9__437_,
  data_head_9__436_,data_head_9__435_,data_head_9__434_,data_head_9__433_,
  data_head_9__432_,data_head_9__431_,data_head_9__430_,data_head_9__429_,
  data_head_9__428_,data_head_9__427_,data_head_9__426_,data_head_9__425_,data_head_9__424_,
  data_head_9__423_,data_head_9__422_,data_head_9__421_,data_head_9__420_,
  data_head_9__419_,data_head_9__418_,data_head_9__417_,data_head_9__416_,data_head_9__415_,
  data_head_9__414_,data_head_9__413_,data_head_9__412_,data_head_9__411_,
  data_head_9__410_,data_head_9__409_,data_head_9__408_,data_head_9__407_,data_head_9__406_,
  data_head_9__405_,data_head_9__404_,data_head_9__403_,data_head_9__402_,
  data_head_9__401_,data_head_9__400_,data_head_9__399_,data_head_9__398_,data_head_9__397_,
  data_head_9__396_,data_head_9__395_,data_head_9__394_,data_head_9__393_,
  data_head_9__392_,data_head_9__391_,data_head_9__390_,data_head_9__389_,
  data_head_9__388_,data_head_9__387_,data_head_9__386_,data_head_9__385_,data_head_9__384_,
  data_head_9__383_,data_head_9__382_,data_head_9__381_,data_head_9__380_,
  data_head_9__379_,data_head_9__378_,data_head_9__377_,data_head_9__376_,data_head_9__375_,
  data_head_9__374_,data_head_9__373_,data_head_9__372_,data_head_9__371_,
  data_head_9__370_,data_head_9__369_,data_head_9__368_,data_head_9__367_,data_head_9__366_,
  data_head_9__365_,data_head_9__364_,data_head_9__363_,data_head_9__362_,
  data_head_9__361_,data_head_9__360_,data_head_9__359_,data_head_9__358_,data_head_9__357_,
  data_head_9__356_,data_head_9__355_,data_head_9__354_,data_head_9__353_,
  data_head_9__352_,data_head_9__351_,data_head_9__350_,data_head_9__349_,
  data_head_9__348_,data_head_9__347_,data_head_9__346_,data_head_9__345_,data_head_9__344_,
  data_head_9__343_,data_head_9__342_,data_head_9__341_,data_head_9__340_,
  data_head_9__339_,data_head_9__338_,data_head_9__337_,data_head_9__336_,data_head_9__335_,
  data_head_9__334_,data_head_9__333_,data_head_9__332_,data_head_9__331_,
  data_head_9__330_,data_head_9__329_,data_head_9__328_,data_head_9__327_,data_head_9__326_,
  data_head_9__325_,data_head_9__324_,data_head_9__323_,data_head_9__322_,
  data_head_9__321_,data_head_9__320_,data_head_9__319_,data_head_9__318_,data_head_9__317_,
  data_head_9__316_,data_head_9__315_,data_head_9__314_,data_head_9__313_,
  data_head_9__312_,data_head_9__311_,data_head_9__310_,data_head_9__309_,
  data_head_9__308_,data_head_9__307_,data_head_9__306_,data_head_9__305_,data_head_9__304_,
  data_head_9__303_,data_head_9__302_,data_head_9__301_,data_head_9__300_,
  data_head_9__299_,data_head_9__298_,data_head_9__297_,data_head_9__296_,data_head_9__295_,
  data_head_9__294_,data_head_9__293_,data_head_9__292_,data_head_9__291_,
  data_head_9__290_,data_head_9__289_,data_head_9__288_,data_head_9__287_,data_head_9__286_,
  data_head_9__285_,data_head_9__284_,data_head_9__283_,data_head_9__282_,
  data_head_9__281_,data_head_9__280_,data_head_9__279_,data_head_9__278_,data_head_9__277_,
  data_head_9__276_,data_head_9__275_,data_head_9__274_,data_head_9__273_,
  data_head_9__272_,data_head_9__271_,data_head_9__270_,data_head_9__269_,
  data_head_9__268_,data_head_9__267_,data_head_9__266_,data_head_9__265_,data_head_9__264_,
  data_head_9__263_,data_head_9__262_,data_head_9__261_,data_head_9__260_,
  data_head_9__259_,data_head_9__258_,data_head_9__257_,data_head_9__256_,data_head_9__255_,
  data_head_9__254_,data_head_9__253_,data_head_9__252_,data_head_9__251_,
  data_head_9__250_,data_head_9__249_,data_head_9__248_,data_head_9__247_,data_head_9__246_,
  data_head_9__245_,data_head_9__244_,data_head_9__243_,data_head_9__242_,
  data_head_9__241_,data_head_9__240_,data_head_9__239_,data_head_9__238_,data_head_9__237_,
  data_head_9__236_,data_head_9__235_,data_head_9__234_,data_head_9__233_,
  data_head_9__232_,data_head_9__231_,data_head_9__230_,data_head_9__229_,
  data_head_9__228_,data_head_9__227_,data_head_9__226_,data_head_9__225_,data_head_9__224_,
  data_head_9__223_,data_head_9__222_,data_head_9__221_,data_head_9__220_,
  data_head_9__219_,data_head_9__218_,data_head_9__217_,data_head_9__216_,data_head_9__215_,
  data_head_9__214_,data_head_9__213_,data_head_9__212_,data_head_9__211_,
  data_head_9__210_,data_head_9__209_,data_head_9__208_,data_head_9__207_,data_head_9__206_,
  data_head_9__205_,data_head_9__204_,data_head_9__203_,data_head_9__202_,
  data_head_9__201_,data_head_9__200_,data_head_9__199_,data_head_9__198_,data_head_9__197_,
  data_head_9__196_,data_head_9__195_,data_head_9__194_,data_head_9__193_,
  data_head_9__192_,data_head_9__191_,data_head_9__190_,data_head_9__189_,
  data_head_9__188_,data_head_9__187_,data_head_9__186_,data_head_9__185_,data_head_9__184_,
  data_head_9__183_,data_head_9__182_,data_head_9__181_,data_head_9__180_,
  data_head_9__179_,data_head_9__178_,data_head_9__177_,data_head_9__176_,data_head_9__175_,
  data_head_9__174_,data_head_9__173_,data_head_9__172_,data_head_9__171_,
  data_head_9__170_,data_head_9__169_,data_head_9__168_,data_head_9__167_,data_head_9__166_,
  data_head_9__165_,data_head_9__164_,data_head_9__163_,data_head_9__162_,
  data_head_9__161_,data_head_9__160_,data_head_9__159_,data_head_9__158_,data_head_9__157_,
  data_head_9__156_,data_head_9__155_,data_head_9__154_,data_head_9__153_,
  data_head_9__152_,data_head_9__151_,data_head_9__150_,data_head_9__149_,
  data_head_9__148_,data_head_9__147_,data_head_9__146_,data_head_9__145_,data_head_9__144_,
  data_head_9__143_,data_head_9__142_,data_head_9__141_,data_head_9__140_,
  data_head_9__139_,data_head_9__138_,data_head_9__137_,data_head_9__136_,data_head_9__135_,
  data_head_9__134_,data_head_9__133_,data_head_9__132_,data_head_9__131_,
  data_head_9__130_,data_head_9__129_,data_head_9__128_,data_head_9__127_,data_head_9__126_,
  data_head_9__125_,data_head_9__124_,data_head_9__123_,data_head_9__122_,
  data_head_9__121_,data_head_9__120_,data_head_9__119_,data_head_9__118_,data_head_9__117_,
  data_head_9__116_,data_head_9__115_,data_head_9__114_,data_head_9__113_,
  data_head_9__112_,data_head_9__111_,data_head_9__110_,data_head_9__109_,
  data_head_9__108_,data_head_9__107_,data_head_9__106_,data_head_9__105_,data_head_9__104_,
  data_head_9__103_,data_head_9__102_,data_head_9__101_,data_head_9__100_,
  data_head_9__99_,data_head_9__98_,data_head_9__97_,data_head_9__96_,data_head_9__95_,
  data_head_9__94_,data_head_9__93_,data_head_9__92_,data_head_9__91_,data_head_9__90_,
  data_head_9__89_,data_head_9__88_,data_head_9__87_,data_head_9__86_,data_head_9__85_,
  data_head_9__84_,data_head_9__83_,data_head_9__82_,data_head_9__81_,
  data_head_9__80_,data_head_9__79_,data_head_9__78_,data_head_9__77_,data_head_9__76_,
  data_head_9__75_,data_head_9__74_,data_head_9__73_,data_head_9__72_,data_head_9__71_,
  data_head_9__70_,data_head_9__69_,data_head_9__68_,data_head_9__67_,
  data_head_9__66_,data_head_9__65_,data_head_9__64_,data_head_9__63_,data_head_9__62_,
  data_head_9__61_,data_head_9__60_,data_head_9__59_,data_head_9__58_,data_head_9__57_,
  data_head_9__56_,data_head_9__55_,data_head_9__54_,data_head_9__53_,
  data_head_9__52_,data_head_9__51_,data_head_9__50_,data_head_9__49_,data_head_9__48_,
  data_head_9__47_,data_head_9__46_,data_head_9__45_,data_head_9__44_,data_head_9__43_,
  data_head_9__42_,data_head_9__41_,data_head_9__40_,data_head_9__39_,data_head_9__38_,
  data_head_9__37_,data_head_9__36_,data_head_9__35_,data_head_9__34_,
  data_head_9__33_,data_head_9__32_,data_head_9__31_,data_head_9__30_,data_head_9__29_,
  data_head_9__28_,data_head_9__27_,data_head_9__26_,data_head_9__25_,data_head_9__24_,
  data_head_9__23_,data_head_9__22_,data_head_9__21_,data_head_9__20_,
  data_head_9__19_,data_head_9__18_,data_head_9__17_,data_head_9__16_,data_head_9__15_,
  data_head_9__14_,data_head_9__13_,data_head_9__12_,data_head_9__11_,data_head_9__10_,
  data_head_9__9_,data_head_9__8_,data_head_9__7_,data_head_9__6_,data_head_9__5_,
  data_head_9__4_,data_head_9__3_,data_head_9__2_,data_head_9__1_,data_head_9__0_,
  n_0_net_,valid_head_9__9_,valid_head_9__8_,valid_head_9__7_,valid_head_9__6_,
  valid_head_9__5_,valid_head_9__4_,valid_head_9__3_,valid_head_9__2_,valid_head_9__1_,
  valid_head_9__0_,n_2_net__9_,n_2_net__8_,n_2_net__7_,n_2_net__6_,n_2_net__5_,
  n_2_net__4_,n_2_net__3_,n_2_net__2_,n_2_net__1_,n_2_net__0_,n_3_net__9_,n_3_net__8_,
  n_3_net__7_,n_3_net__6_,n_3_net__5_,n_3_net__4_,n_3_net__3_,n_3_net__2_,
  n_3_net__1_,n_3_net__0_,ready_head_9__9_,ready_head_9__8_,ready_head_9__7_,
  ready_head_9__6_,ready_head_9__5_,ready_head_9__4_,ready_head_9__3_,ready_head_9__2_,
  ready_head_9__1_,ready_head_9__0_,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,
  n_4_net__639_,n_4_net__638_,n_4_net__637_,n_4_net__636_,n_4_net__635_,n_4_net__634_,
  n_4_net__633_,n_4_net__632_,n_4_net__631_,n_4_net__630_,n_4_net__629_,
  n_4_net__628_,n_4_net__627_,n_4_net__626_,n_4_net__625_,n_4_net__624_,n_4_net__623_,
  n_4_net__622_,n_4_net__621_,n_4_net__620_,n_4_net__619_,n_4_net__618_,n_4_net__617_,
  n_4_net__616_,n_4_net__615_,n_4_net__614_,n_4_net__613_,n_4_net__612_,n_4_net__611_,
  n_4_net__610_,n_4_net__609_,n_4_net__608_,n_4_net__607_,n_4_net__606_,
  n_4_net__605_,n_4_net__604_,n_4_net__603_,n_4_net__602_,n_4_net__601_,n_4_net__600_,
  n_4_net__599_,n_4_net__598_,n_4_net__597_,n_4_net__596_,n_4_net__595_,n_4_net__594_,
  n_4_net__593_,n_4_net__592_,n_4_net__591_,n_4_net__590_,n_4_net__589_,
  n_4_net__588_,n_4_net__587_,n_4_net__586_,n_4_net__585_,n_4_net__584_,n_4_net__583_,
  n_4_net__582_,n_4_net__581_,n_4_net__580_,n_4_net__579_,n_4_net__578_,n_4_net__577_,
  n_4_net__576_,n_4_net__575_,n_4_net__574_,n_4_net__573_,n_4_net__572_,n_4_net__571_,
  n_4_net__570_,n_4_net__569_,n_4_net__568_,n_4_net__567_,n_4_net__566_,
  n_4_net__565_,n_4_net__564_,n_4_net__563_,n_4_net__562_,n_4_net__561_,n_4_net__560_,
  n_4_net__559_,n_4_net__558_,n_4_net__557_,n_4_net__556_,n_4_net__555_,n_4_net__554_,
  n_4_net__553_,n_4_net__552_,n_4_net__551_,n_4_net__550_,n_4_net__549_,
  n_4_net__548_,n_4_net__547_,n_4_net__546_,n_4_net__545_,n_4_net__544_,n_4_net__543_,
  n_4_net__542_,n_4_net__541_,n_4_net__540_,n_4_net__539_,n_4_net__538_,n_4_net__537_,
  n_4_net__536_,n_4_net__535_,n_4_net__534_,n_4_net__533_,n_4_net__532_,n_4_net__531_,
  n_4_net__530_,n_4_net__529_,n_4_net__528_,n_4_net__527_,n_4_net__526_,
  n_4_net__525_,n_4_net__524_,n_4_net__523_,n_4_net__522_,n_4_net__521_,n_4_net__520_,
  n_4_net__519_,n_4_net__518_,n_4_net__517_,n_4_net__516_,n_4_net__515_,n_4_net__514_,
  n_4_net__513_,n_4_net__512_,n_4_net__511_,n_4_net__510_,n_4_net__509_,
  n_4_net__508_,n_4_net__507_,n_4_net__506_,n_4_net__505_,n_4_net__504_,n_4_net__503_,
  n_4_net__502_,n_4_net__501_,n_4_net__500_,n_4_net__499_,n_4_net__498_,n_4_net__497_,
  n_4_net__496_,n_4_net__495_,n_4_net__494_,n_4_net__493_,n_4_net__492_,n_4_net__491_,
  n_4_net__490_,n_4_net__489_,n_4_net__488_,n_4_net__487_,n_4_net__486_,
  n_4_net__485_,n_4_net__484_,n_4_net__483_,n_4_net__482_,n_4_net__481_,n_4_net__480_,
  n_4_net__479_,n_4_net__478_,n_4_net__477_,n_4_net__476_,n_4_net__475_,n_4_net__474_,
  n_4_net__473_,n_4_net__472_,n_4_net__471_,n_4_net__470_,n_4_net__469_,
  n_4_net__468_,n_4_net__467_,n_4_net__466_,n_4_net__465_,n_4_net__464_,n_4_net__463_,
  n_4_net__462_,n_4_net__461_,n_4_net__460_,n_4_net__459_,n_4_net__458_,n_4_net__457_,
  n_4_net__456_,n_4_net__455_,n_4_net__454_,n_4_net__453_,n_4_net__452_,n_4_net__451_,
  n_4_net__450_,n_4_net__449_,n_4_net__448_,n_4_net__447_,n_4_net__446_,
  n_4_net__445_,n_4_net__444_,n_4_net__443_,n_4_net__442_,n_4_net__441_,n_4_net__440_,
  n_4_net__439_,n_4_net__438_,n_4_net__437_,n_4_net__436_,n_4_net__435_,n_4_net__434_,
  n_4_net__433_,n_4_net__432_,n_4_net__431_,n_4_net__430_,n_4_net__429_,
  n_4_net__428_,n_4_net__427_,n_4_net__426_,n_4_net__425_,n_4_net__424_,n_4_net__423_,
  n_4_net__422_,n_4_net__421_,n_4_net__420_,n_4_net__419_,n_4_net__418_,n_4_net__417_,
  n_4_net__416_,n_4_net__415_,n_4_net__414_,n_4_net__413_,n_4_net__412_,n_4_net__411_,
  n_4_net__410_,n_4_net__409_,n_4_net__408_,n_4_net__407_,n_4_net__406_,
  n_4_net__405_,n_4_net__404_,n_4_net__403_,n_4_net__402_,n_4_net__401_,n_4_net__400_,
  n_4_net__399_,n_4_net__398_,n_4_net__397_,n_4_net__396_,n_4_net__395_,n_4_net__394_,
  n_4_net__393_,n_4_net__392_,n_4_net__391_,n_4_net__390_,n_4_net__389_,
  n_4_net__388_,n_4_net__387_,n_4_net__386_,n_4_net__385_,n_4_net__384_,n_4_net__383_,
  n_4_net__382_,n_4_net__381_,n_4_net__380_,n_4_net__379_,n_4_net__378_,n_4_net__377_,
  n_4_net__376_,n_4_net__375_,n_4_net__374_,n_4_net__373_,n_4_net__372_,n_4_net__371_,
  n_4_net__370_,n_4_net__369_,n_4_net__368_,n_4_net__367_,n_4_net__366_,
  n_4_net__365_,n_4_net__364_,n_4_net__363_,n_4_net__362_,n_4_net__361_,n_4_net__360_,
  n_4_net__359_,n_4_net__358_,n_4_net__357_,n_4_net__356_,n_4_net__355_,n_4_net__354_,
  n_4_net__353_,n_4_net__352_,n_4_net__351_,n_4_net__350_,n_4_net__349_,
  n_4_net__348_,n_4_net__347_,n_4_net__346_,n_4_net__345_,n_4_net__344_,n_4_net__343_,
  n_4_net__342_,n_4_net__341_,n_4_net__340_,n_4_net__339_,n_4_net__338_,n_4_net__337_,
  n_4_net__336_,n_4_net__335_,n_4_net__334_,n_4_net__333_,n_4_net__332_,n_4_net__331_,
  n_4_net__330_,n_4_net__329_,n_4_net__328_,n_4_net__327_,n_4_net__326_,
  n_4_net__325_,n_4_net__324_,n_4_net__323_,n_4_net__322_,n_4_net__321_,n_4_net__320_,
  n_4_net__319_,n_4_net__318_,n_4_net__317_,n_4_net__316_,n_4_net__315_,n_4_net__314_,
  n_4_net__313_,n_4_net__312_,n_4_net__311_,n_4_net__310_,n_4_net__309_,
  n_4_net__308_,n_4_net__307_,n_4_net__306_,n_4_net__305_,n_4_net__304_,n_4_net__303_,
  n_4_net__302_,n_4_net__301_,n_4_net__300_,n_4_net__299_,n_4_net__298_,n_4_net__297_,
  n_4_net__296_,n_4_net__295_,n_4_net__294_,n_4_net__293_,n_4_net__292_,n_4_net__291_,
  n_4_net__290_,n_4_net__289_,n_4_net__288_,n_4_net__287_,n_4_net__286_,
  n_4_net__285_,n_4_net__284_,n_4_net__283_,n_4_net__282_,n_4_net__281_,n_4_net__280_,
  n_4_net__279_,n_4_net__278_,n_4_net__277_,n_4_net__276_,n_4_net__275_,n_4_net__274_,
  n_4_net__273_,n_4_net__272_,n_4_net__271_,n_4_net__270_,n_4_net__269_,
  n_4_net__268_,n_4_net__267_,n_4_net__266_,n_4_net__265_,n_4_net__264_,n_4_net__263_,
  n_4_net__262_,n_4_net__261_,n_4_net__260_,n_4_net__259_,n_4_net__258_,n_4_net__257_,
  n_4_net__256_,n_4_net__255_,n_4_net__254_,n_4_net__253_,n_4_net__252_,n_4_net__251_,
  n_4_net__250_,n_4_net__249_,n_4_net__248_,n_4_net__247_,n_4_net__246_,
  n_4_net__245_,n_4_net__244_,n_4_net__243_,n_4_net__242_,n_4_net__241_,n_4_net__240_,
  n_4_net__239_,n_4_net__238_,n_4_net__237_,n_4_net__236_,n_4_net__235_,n_4_net__234_,
  n_4_net__233_,n_4_net__232_,n_4_net__231_,n_4_net__230_,n_4_net__229_,
  n_4_net__228_,n_4_net__227_,n_4_net__226_,n_4_net__225_,n_4_net__224_,n_4_net__223_,
  n_4_net__222_,n_4_net__221_,n_4_net__220_,n_4_net__219_,n_4_net__218_,n_4_net__217_,
  n_4_net__216_,n_4_net__215_,n_4_net__214_,n_4_net__213_,n_4_net__212_,n_4_net__211_,
  n_4_net__210_,n_4_net__209_,n_4_net__208_,n_4_net__207_,n_4_net__206_,
  n_4_net__205_,n_4_net__204_,n_4_net__203_,n_4_net__202_,n_4_net__201_,n_4_net__200_,
  n_4_net__199_,n_4_net__198_,n_4_net__197_,n_4_net__196_,n_4_net__195_,n_4_net__194_,
  n_4_net__193_,n_4_net__192_,n_4_net__191_,n_4_net__190_,n_4_net__189_,
  n_4_net__188_,n_4_net__187_,n_4_net__186_,n_4_net__185_,n_4_net__184_,n_4_net__183_,
  n_4_net__182_,n_4_net__181_,n_4_net__180_,n_4_net__179_,n_4_net__178_,n_4_net__177_,
  n_4_net__176_,n_4_net__175_,n_4_net__174_,n_4_net__173_,n_4_net__172_,n_4_net__171_,
  n_4_net__170_,n_4_net__169_,n_4_net__168_,n_4_net__167_,n_4_net__166_,
  n_4_net__165_,n_4_net__164_,n_4_net__163_,n_4_net__162_,n_4_net__161_,n_4_net__160_,
  n_4_net__159_,n_4_net__158_,n_4_net__157_,n_4_net__156_,n_4_net__155_,n_4_net__154_,
  n_4_net__153_,n_4_net__152_,n_4_net__151_,n_4_net__150_,n_4_net__149_,
  n_4_net__148_,n_4_net__147_,n_4_net__146_,n_4_net__145_,n_4_net__144_,n_4_net__143_,
  n_4_net__142_,n_4_net__141_,n_4_net__140_,n_4_net__139_,n_4_net__138_,n_4_net__137_,
  n_4_net__136_,n_4_net__135_,n_4_net__134_,n_4_net__133_,n_4_net__132_,n_4_net__131_,
  n_4_net__130_,n_4_net__129_,n_4_net__128_,n_4_net__127_,n_4_net__126_,
  n_4_net__125_,n_4_net__124_,n_4_net__123_,n_4_net__122_,n_4_net__121_,n_4_net__120_,
  n_4_net__119_,n_4_net__118_,n_4_net__117_,n_4_net__116_,n_4_net__115_,n_4_net__114_,
  n_4_net__113_,n_4_net__112_,n_4_net__111_,n_4_net__110_,n_4_net__109_,
  n_4_net__108_,n_4_net__107_,n_4_net__106_,n_4_net__105_,n_4_net__104_,n_4_net__103_,
  n_4_net__102_,n_4_net__101_,n_4_net__100_,n_4_net__99_,n_4_net__98_,n_4_net__97_,
  n_4_net__96_,n_4_net__95_,n_4_net__94_,n_4_net__93_,n_4_net__92_,n_4_net__91_,
  n_4_net__90_,n_4_net__89_,n_4_net__88_,n_4_net__87_,n_4_net__86_,n_4_net__85_,
  n_4_net__84_,n_4_net__83_,n_4_net__82_,n_4_net__81_,n_4_net__80_,n_4_net__79_,n_4_net__78_,
  n_4_net__77_,n_4_net__76_,n_4_net__75_,n_4_net__74_,n_4_net__73_,n_4_net__72_,
  n_4_net__71_,n_4_net__70_,n_4_net__69_,n_4_net__68_,n_4_net__67_,n_4_net__66_,
  n_4_net__65_,n_4_net__64_,n_4_net__63_,n_4_net__62_,n_4_net__61_,n_4_net__60_,
  n_4_net__59_,n_4_net__58_,n_4_net__57_,n_4_net__56_,n_4_net__55_,n_4_net__54_,
  n_4_net__53_,n_4_net__52_,n_4_net__51_,n_4_net__50_,n_4_net__49_,n_4_net__48_,
  n_4_net__47_,n_4_net__46_,n_4_net__45_,n_4_net__44_,n_4_net__43_,n_4_net__42_,
  n_4_net__41_,n_4_net__40_,n_4_net__39_,n_4_net__38_,n_4_net__37_,n_4_net__36_,n_4_net__35_,
  n_4_net__34_,n_4_net__33_,n_4_net__32_,n_4_net__31_,n_4_net__30_,n_4_net__29_,
  n_4_net__28_,n_4_net__27_,n_4_net__26_,n_4_net__25_,n_4_net__24_,n_4_net__23_,
  n_4_net__22_,n_4_net__21_,n_4_net__20_,n_4_net__19_,n_4_net__18_,n_4_net__17_,
  n_4_net__16_,n_4_net__15_,n_4_net__14_,n_4_net__13_,n_4_net__12_,n_4_net__11_,
  n_4_net__10_,n_4_net__9_,n_4_net__8_,n_4_net__7_,n_4_net__6_,n_4_net__5_,n_4_net__4_,
  n_4_net__3_,n_4_net__2_,n_4_net__1_,n_4_net__0_,N165,N166,N167,N168,N169,N170,N171,
  N172,N173,N174,n_5_net_,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184;
  wire [3:0] go_cnt;

  bsg_make_2D_array_width_p64_items_p10
  bm2Da
  (
    .i(data_o_flat),
    .o(data_o)
  );


  bsg_rr_f2f_input_width_p64_num_in_p10_middle_meet_p10
  ic_9__in_chan_bsg_rr_ff_in
  (
    .clk(clk),
    .reset(n_0_net_),
    .valid_i(valid_i),
    .data_i(data_i),
    .data_head_o({ data_head_9__639_, data_head_9__638_, data_head_9__637_, data_head_9__636_, data_head_9__635_, data_head_9__634_, data_head_9__633_, data_head_9__632_, data_head_9__631_, data_head_9__630_, data_head_9__629_, data_head_9__628_, data_head_9__627_, data_head_9__626_, data_head_9__625_, data_head_9__624_, data_head_9__623_, data_head_9__622_, data_head_9__621_, data_head_9__620_, data_head_9__619_, data_head_9__618_, data_head_9__617_, data_head_9__616_, data_head_9__615_, data_head_9__614_, data_head_9__613_, data_head_9__612_, data_head_9__611_, data_head_9__610_, data_head_9__609_, data_head_9__608_, data_head_9__607_, data_head_9__606_, data_head_9__605_, data_head_9__604_, data_head_9__603_, data_head_9__602_, data_head_9__601_, data_head_9__600_, data_head_9__599_, data_head_9__598_, data_head_9__597_, data_head_9__596_, data_head_9__595_, data_head_9__594_, data_head_9__593_, data_head_9__592_, data_head_9__591_, data_head_9__590_, data_head_9__589_, data_head_9__588_, data_head_9__587_, data_head_9__586_, data_head_9__585_, data_head_9__584_, data_head_9__583_, data_head_9__582_, data_head_9__581_, data_head_9__580_, data_head_9__579_, data_head_9__578_, data_head_9__577_, data_head_9__576_, data_head_9__575_, data_head_9__574_, data_head_9__573_, data_head_9__572_, data_head_9__571_, data_head_9__570_, data_head_9__569_, data_head_9__568_, data_head_9__567_, data_head_9__566_, data_head_9__565_, data_head_9__564_, data_head_9__563_, data_head_9__562_, data_head_9__561_, data_head_9__560_, data_head_9__559_, data_head_9__558_, data_head_9__557_, data_head_9__556_, data_head_9__555_, data_head_9__554_, data_head_9__553_, data_head_9__552_, data_head_9__551_, data_head_9__550_, data_head_9__549_, data_head_9__548_, data_head_9__547_, data_head_9__546_, data_head_9__545_, data_head_9__544_, data_head_9__543_, data_head_9__542_, data_head_9__541_, data_head_9__540_, data_head_9__539_, data_head_9__538_, data_head_9__537_, data_head_9__536_, data_head_9__535_, data_head_9__534_, data_head_9__533_, data_head_9__532_, data_head_9__531_, data_head_9__530_, data_head_9__529_, data_head_9__528_, data_head_9__527_, data_head_9__526_, data_head_9__525_, data_head_9__524_, data_head_9__523_, data_head_9__522_, data_head_9__521_, data_head_9__520_, data_head_9__519_, data_head_9__518_, data_head_9__517_, data_head_9__516_, data_head_9__515_, data_head_9__514_, data_head_9__513_, data_head_9__512_, data_head_9__511_, data_head_9__510_, data_head_9__509_, data_head_9__508_, data_head_9__507_, data_head_9__506_, data_head_9__505_, data_head_9__504_, data_head_9__503_, data_head_9__502_, data_head_9__501_, data_head_9__500_, data_head_9__499_, data_head_9__498_, data_head_9__497_, data_head_9__496_, data_head_9__495_, data_head_9__494_, data_head_9__493_, data_head_9__492_, data_head_9__491_, data_head_9__490_, data_head_9__489_, data_head_9__488_, data_head_9__487_, data_head_9__486_, data_head_9__485_, data_head_9__484_, data_head_9__483_, data_head_9__482_, data_head_9__481_, data_head_9__480_, data_head_9__479_, data_head_9__478_, data_head_9__477_, data_head_9__476_, data_head_9__475_, data_head_9__474_, data_head_9__473_, data_head_9__472_, data_head_9__471_, data_head_9__470_, data_head_9__469_, data_head_9__468_, data_head_9__467_, data_head_9__466_, data_head_9__465_, data_head_9__464_, data_head_9__463_, data_head_9__462_, data_head_9__461_, data_head_9__460_, data_head_9__459_, data_head_9__458_, data_head_9__457_, data_head_9__456_, data_head_9__455_, data_head_9__454_, data_head_9__453_, data_head_9__452_, data_head_9__451_, data_head_9__450_, data_head_9__449_, data_head_9__448_, data_head_9__447_, data_head_9__446_, data_head_9__445_, data_head_9__444_, data_head_9__443_, data_head_9__442_, data_head_9__441_, data_head_9__440_, data_head_9__439_, data_head_9__438_, data_head_9__437_, data_head_9__436_, data_head_9__435_, data_head_9__434_, data_head_9__433_, data_head_9__432_, data_head_9__431_, data_head_9__430_, data_head_9__429_, data_head_9__428_, data_head_9__427_, data_head_9__426_, data_head_9__425_, data_head_9__424_, data_head_9__423_, data_head_9__422_, data_head_9__421_, data_head_9__420_, data_head_9__419_, data_head_9__418_, data_head_9__417_, data_head_9__416_, data_head_9__415_, data_head_9__414_, data_head_9__413_, data_head_9__412_, data_head_9__411_, data_head_9__410_, data_head_9__409_, data_head_9__408_, data_head_9__407_, data_head_9__406_, data_head_9__405_, data_head_9__404_, data_head_9__403_, data_head_9__402_, data_head_9__401_, data_head_9__400_, data_head_9__399_, data_head_9__398_, data_head_9__397_, data_head_9__396_, data_head_9__395_, data_head_9__394_, data_head_9__393_, data_head_9__392_, data_head_9__391_, data_head_9__390_, data_head_9__389_, data_head_9__388_, data_head_9__387_, data_head_9__386_, data_head_9__385_, data_head_9__384_, data_head_9__383_, data_head_9__382_, data_head_9__381_, data_head_9__380_, data_head_9__379_, data_head_9__378_, data_head_9__377_, data_head_9__376_, data_head_9__375_, data_head_9__374_, data_head_9__373_, data_head_9__372_, data_head_9__371_, data_head_9__370_, data_head_9__369_, data_head_9__368_, data_head_9__367_, data_head_9__366_, data_head_9__365_, data_head_9__364_, data_head_9__363_, data_head_9__362_, data_head_9__361_, data_head_9__360_, data_head_9__359_, data_head_9__358_, data_head_9__357_, data_head_9__356_, data_head_9__355_, data_head_9__354_, data_head_9__353_, data_head_9__352_, data_head_9__351_, data_head_9__350_, data_head_9__349_, data_head_9__348_, data_head_9__347_, data_head_9__346_, data_head_9__345_, data_head_9__344_, data_head_9__343_, data_head_9__342_, data_head_9__341_, data_head_9__340_, data_head_9__339_, data_head_9__338_, data_head_9__337_, data_head_9__336_, data_head_9__335_, data_head_9__334_, data_head_9__333_, data_head_9__332_, data_head_9__331_, data_head_9__330_, data_head_9__329_, data_head_9__328_, data_head_9__327_, data_head_9__326_, data_head_9__325_, data_head_9__324_, data_head_9__323_, data_head_9__322_, data_head_9__321_, data_head_9__320_, data_head_9__319_, data_head_9__318_, data_head_9__317_, data_head_9__316_, data_head_9__315_, data_head_9__314_, data_head_9__313_, data_head_9__312_, data_head_9__311_, data_head_9__310_, data_head_9__309_, data_head_9__308_, data_head_9__307_, data_head_9__306_, data_head_9__305_, data_head_9__304_, data_head_9__303_, data_head_9__302_, data_head_9__301_, data_head_9__300_, data_head_9__299_, data_head_9__298_, data_head_9__297_, data_head_9__296_, data_head_9__295_, data_head_9__294_, data_head_9__293_, data_head_9__292_, data_head_9__291_, data_head_9__290_, data_head_9__289_, data_head_9__288_, data_head_9__287_, data_head_9__286_, data_head_9__285_, data_head_9__284_, data_head_9__283_, data_head_9__282_, data_head_9__281_, data_head_9__280_, data_head_9__279_, data_head_9__278_, data_head_9__277_, data_head_9__276_, data_head_9__275_, data_head_9__274_, data_head_9__273_, data_head_9__272_, data_head_9__271_, data_head_9__270_, data_head_9__269_, data_head_9__268_, data_head_9__267_, data_head_9__266_, data_head_9__265_, data_head_9__264_, data_head_9__263_, data_head_9__262_, data_head_9__261_, data_head_9__260_, data_head_9__259_, data_head_9__258_, data_head_9__257_, data_head_9__256_, data_head_9__255_, data_head_9__254_, data_head_9__253_, data_head_9__252_, data_head_9__251_, data_head_9__250_, data_head_9__249_, data_head_9__248_, data_head_9__247_, data_head_9__246_, data_head_9__245_, data_head_9__244_, data_head_9__243_, data_head_9__242_, data_head_9__241_, data_head_9__240_, data_head_9__239_, data_head_9__238_, data_head_9__237_, data_head_9__236_, data_head_9__235_, data_head_9__234_, data_head_9__233_, data_head_9__232_, data_head_9__231_, data_head_9__230_, data_head_9__229_, data_head_9__228_, data_head_9__227_, data_head_9__226_, data_head_9__225_, data_head_9__224_, data_head_9__223_, data_head_9__222_, data_head_9__221_, data_head_9__220_, data_head_9__219_, data_head_9__218_, data_head_9__217_, data_head_9__216_, data_head_9__215_, data_head_9__214_, data_head_9__213_, data_head_9__212_, data_head_9__211_, data_head_9__210_, data_head_9__209_, data_head_9__208_, data_head_9__207_, data_head_9__206_, data_head_9__205_, data_head_9__204_, data_head_9__203_, data_head_9__202_, data_head_9__201_, data_head_9__200_, data_head_9__199_, data_head_9__198_, data_head_9__197_, data_head_9__196_, data_head_9__195_, data_head_9__194_, data_head_9__193_, data_head_9__192_, data_head_9__191_, data_head_9__190_, data_head_9__189_, data_head_9__188_, data_head_9__187_, data_head_9__186_, data_head_9__185_, data_head_9__184_, data_head_9__183_, data_head_9__182_, data_head_9__181_, data_head_9__180_, data_head_9__179_, data_head_9__178_, data_head_9__177_, data_head_9__176_, data_head_9__175_, data_head_9__174_, data_head_9__173_, data_head_9__172_, data_head_9__171_, data_head_9__170_, data_head_9__169_, data_head_9__168_, data_head_9__167_, data_head_9__166_, data_head_9__165_, data_head_9__164_, data_head_9__163_, data_head_9__162_, data_head_9__161_, data_head_9__160_, data_head_9__159_, data_head_9__158_, data_head_9__157_, data_head_9__156_, data_head_9__155_, data_head_9__154_, data_head_9__153_, data_head_9__152_, data_head_9__151_, data_head_9__150_, data_head_9__149_, data_head_9__148_, data_head_9__147_, data_head_9__146_, data_head_9__145_, data_head_9__144_, data_head_9__143_, data_head_9__142_, data_head_9__141_, data_head_9__140_, data_head_9__139_, data_head_9__138_, data_head_9__137_, data_head_9__136_, data_head_9__135_, data_head_9__134_, data_head_9__133_, data_head_9__132_, data_head_9__131_, data_head_9__130_, data_head_9__129_, data_head_9__128_, data_head_9__127_, data_head_9__126_, data_head_9__125_, data_head_9__124_, data_head_9__123_, data_head_9__122_, data_head_9__121_, data_head_9__120_, data_head_9__119_, data_head_9__118_, data_head_9__117_, data_head_9__116_, data_head_9__115_, data_head_9__114_, data_head_9__113_, data_head_9__112_, data_head_9__111_, data_head_9__110_, data_head_9__109_, data_head_9__108_, data_head_9__107_, data_head_9__106_, data_head_9__105_, data_head_9__104_, data_head_9__103_, data_head_9__102_, data_head_9__101_, data_head_9__100_, data_head_9__99_, data_head_9__98_, data_head_9__97_, data_head_9__96_, data_head_9__95_, data_head_9__94_, data_head_9__93_, data_head_9__92_, data_head_9__91_, data_head_9__90_, data_head_9__89_, data_head_9__88_, data_head_9__87_, data_head_9__86_, data_head_9__85_, data_head_9__84_, data_head_9__83_, data_head_9__82_, data_head_9__81_, data_head_9__80_, data_head_9__79_, data_head_9__78_, data_head_9__77_, data_head_9__76_, data_head_9__75_, data_head_9__74_, data_head_9__73_, data_head_9__72_, data_head_9__71_, data_head_9__70_, data_head_9__69_, data_head_9__68_, data_head_9__67_, data_head_9__66_, data_head_9__65_, data_head_9__64_, data_head_9__63_, data_head_9__62_, data_head_9__61_, data_head_9__60_, data_head_9__59_, data_head_9__58_, data_head_9__57_, data_head_9__56_, data_head_9__55_, data_head_9__54_, data_head_9__53_, data_head_9__52_, data_head_9__51_, data_head_9__50_, data_head_9__49_, data_head_9__48_, data_head_9__47_, data_head_9__46_, data_head_9__45_, data_head_9__44_, data_head_9__43_, data_head_9__42_, data_head_9__41_, data_head_9__40_, data_head_9__39_, data_head_9__38_, data_head_9__37_, data_head_9__36_, data_head_9__35_, data_head_9__34_, data_head_9__33_, data_head_9__32_, data_head_9__31_, data_head_9__30_, data_head_9__29_, data_head_9__28_, data_head_9__27_, data_head_9__26_, data_head_9__25_, data_head_9__24_, data_head_9__23_, data_head_9__22_, data_head_9__21_, data_head_9__20_, data_head_9__19_, data_head_9__18_, data_head_9__17_, data_head_9__16_, data_head_9__15_, data_head_9__14_, data_head_9__13_, data_head_9__12_, data_head_9__11_, data_head_9__10_, data_head_9__9_, data_head_9__8_, data_head_9__7_, data_head_9__6_, data_head_9__5_, data_head_9__4_, data_head_9__3_, data_head_9__2_, data_head_9__1_, data_head_9__0_ }),
    .valid_head_o({ valid_head_9__9_, valid_head_9__8_, valid_head_9__7_, valid_head_9__6_, valid_head_9__5_, valid_head_9__4_, valid_head_9__3_, valid_head_9__2_, valid_head_9__1_, valid_head_9__0_ }),
    .go_channels_i(go_channels),
    .go_cnt_i(go_cnt),
    .yumi_o({ yumi_int_o_9__9_, yumi_int_o_9__8_, yumi_int_o_9__7_, yumi_int_o_9__6_, yumi_int_o_9__5_, yumi_int_o_9__4_, yumi_int_o_9__3_, yumi_int_o_9__2_, yumi_int_o_9__1_, yumi_int_o_9__0_ })
  );


  bsg_rr_f2f_middle_width_p64_middle_meet_p10
  brrf2fm
  (
    .valid_head_i({ n_2_net__9_, n_2_net__8_, n_2_net__7_, n_2_net__6_, n_2_net__5_, n_2_net__4_, n_2_net__3_, n_2_net__2_, n_2_net__1_, n_2_net__0_ }),
    .ready_head_i({ n_3_net__9_, n_3_net__8_, n_3_net__7_, n_3_net__6_, n_3_net__5_, n_3_net__4_, n_3_net__3_, n_3_net__2_, n_3_net__1_, n_3_net__0_ }),
    .go_channels_o(go_channels),
    .go_cnt_o(go_cnt)
  );


  bsg_make_2D_array_width_p64_items_p10
  oc_9__out_chan_bm2Da
  (
    .i({ n_4_net__639_, n_4_net__638_, n_4_net__637_, n_4_net__636_, n_4_net__635_, n_4_net__634_, n_4_net__633_, n_4_net__632_, n_4_net__631_, n_4_net__630_, n_4_net__629_, n_4_net__628_, n_4_net__627_, n_4_net__626_, n_4_net__625_, n_4_net__624_, n_4_net__623_, n_4_net__622_, n_4_net__621_, n_4_net__620_, n_4_net__619_, n_4_net__618_, n_4_net__617_, n_4_net__616_, n_4_net__615_, n_4_net__614_, n_4_net__613_, n_4_net__612_, n_4_net__611_, n_4_net__610_, n_4_net__609_, n_4_net__608_, n_4_net__607_, n_4_net__606_, n_4_net__605_, n_4_net__604_, n_4_net__603_, n_4_net__602_, n_4_net__601_, n_4_net__600_, n_4_net__599_, n_4_net__598_, n_4_net__597_, n_4_net__596_, n_4_net__595_, n_4_net__594_, n_4_net__593_, n_4_net__592_, n_4_net__591_, n_4_net__590_, n_4_net__589_, n_4_net__588_, n_4_net__587_, n_4_net__586_, n_4_net__585_, n_4_net__584_, n_4_net__583_, n_4_net__582_, n_4_net__581_, n_4_net__580_, n_4_net__579_, n_4_net__578_, n_4_net__577_, n_4_net__576_, n_4_net__575_, n_4_net__574_, n_4_net__573_, n_4_net__572_, n_4_net__571_, n_4_net__570_, n_4_net__569_, n_4_net__568_, n_4_net__567_, n_4_net__566_, n_4_net__565_, n_4_net__564_, n_4_net__563_, n_4_net__562_, n_4_net__561_, n_4_net__560_, n_4_net__559_, n_4_net__558_, n_4_net__557_, n_4_net__556_, n_4_net__555_, n_4_net__554_, n_4_net__553_, n_4_net__552_, n_4_net__551_, n_4_net__550_, n_4_net__549_, n_4_net__548_, n_4_net__547_, n_4_net__546_, n_4_net__545_, n_4_net__544_, n_4_net__543_, n_4_net__542_, n_4_net__541_, n_4_net__540_, n_4_net__539_, n_4_net__538_, n_4_net__537_, n_4_net__536_, n_4_net__535_, n_4_net__534_, n_4_net__533_, n_4_net__532_, n_4_net__531_, n_4_net__530_, n_4_net__529_, n_4_net__528_, n_4_net__527_, n_4_net__526_, n_4_net__525_, n_4_net__524_, n_4_net__523_, n_4_net__522_, n_4_net__521_, n_4_net__520_, n_4_net__519_, n_4_net__518_, n_4_net__517_, n_4_net__516_, n_4_net__515_, n_4_net__514_, n_4_net__513_, n_4_net__512_, n_4_net__511_, n_4_net__510_, n_4_net__509_, n_4_net__508_, n_4_net__507_, n_4_net__506_, n_4_net__505_, n_4_net__504_, n_4_net__503_, n_4_net__502_, n_4_net__501_, n_4_net__500_, n_4_net__499_, n_4_net__498_, n_4_net__497_, n_4_net__496_, n_4_net__495_, n_4_net__494_, n_4_net__493_, n_4_net__492_, n_4_net__491_, n_4_net__490_, n_4_net__489_, n_4_net__488_, n_4_net__487_, n_4_net__486_, n_4_net__485_, n_4_net__484_, n_4_net__483_, n_4_net__482_, n_4_net__481_, n_4_net__480_, n_4_net__479_, n_4_net__478_, n_4_net__477_, n_4_net__476_, n_4_net__475_, n_4_net__474_, n_4_net__473_, n_4_net__472_, n_4_net__471_, n_4_net__470_, n_4_net__469_, n_4_net__468_, n_4_net__467_, n_4_net__466_, n_4_net__465_, n_4_net__464_, n_4_net__463_, n_4_net__462_, n_4_net__461_, n_4_net__460_, n_4_net__459_, n_4_net__458_, n_4_net__457_, n_4_net__456_, n_4_net__455_, n_4_net__454_, n_4_net__453_, n_4_net__452_, n_4_net__451_, n_4_net__450_, n_4_net__449_, n_4_net__448_, n_4_net__447_, n_4_net__446_, n_4_net__445_, n_4_net__444_, n_4_net__443_, n_4_net__442_, n_4_net__441_, n_4_net__440_, n_4_net__439_, n_4_net__438_, n_4_net__437_, n_4_net__436_, n_4_net__435_, n_4_net__434_, n_4_net__433_, n_4_net__432_, n_4_net__431_, n_4_net__430_, n_4_net__429_, n_4_net__428_, n_4_net__427_, n_4_net__426_, n_4_net__425_, n_4_net__424_, n_4_net__423_, n_4_net__422_, n_4_net__421_, n_4_net__420_, n_4_net__419_, n_4_net__418_, n_4_net__417_, n_4_net__416_, n_4_net__415_, n_4_net__414_, n_4_net__413_, n_4_net__412_, n_4_net__411_, n_4_net__410_, n_4_net__409_, n_4_net__408_, n_4_net__407_, n_4_net__406_, n_4_net__405_, n_4_net__404_, n_4_net__403_, n_4_net__402_, n_4_net__401_, n_4_net__400_, n_4_net__399_, n_4_net__398_, n_4_net__397_, n_4_net__396_, n_4_net__395_, n_4_net__394_, n_4_net__393_, n_4_net__392_, n_4_net__391_, n_4_net__390_, n_4_net__389_, n_4_net__388_, n_4_net__387_, n_4_net__386_, n_4_net__385_, n_4_net__384_, n_4_net__383_, n_4_net__382_, n_4_net__381_, n_4_net__380_, n_4_net__379_, n_4_net__378_, n_4_net__377_, n_4_net__376_, n_4_net__375_, n_4_net__374_, n_4_net__373_, n_4_net__372_, n_4_net__371_, n_4_net__370_, n_4_net__369_, n_4_net__368_, n_4_net__367_, n_4_net__366_, n_4_net__365_, n_4_net__364_, n_4_net__363_, n_4_net__362_, n_4_net__361_, n_4_net__360_, n_4_net__359_, n_4_net__358_, n_4_net__357_, n_4_net__356_, n_4_net__355_, n_4_net__354_, n_4_net__353_, n_4_net__352_, n_4_net__351_, n_4_net__350_, n_4_net__349_, n_4_net__348_, n_4_net__347_, n_4_net__346_, n_4_net__345_, n_4_net__344_, n_4_net__343_, n_4_net__342_, n_4_net__341_, n_4_net__340_, n_4_net__339_, n_4_net__338_, n_4_net__337_, n_4_net__336_, n_4_net__335_, n_4_net__334_, n_4_net__333_, n_4_net__332_, n_4_net__331_, n_4_net__330_, n_4_net__329_, n_4_net__328_, n_4_net__327_, n_4_net__326_, n_4_net__325_, n_4_net__324_, n_4_net__323_, n_4_net__322_, n_4_net__321_, n_4_net__320_, n_4_net__319_, n_4_net__318_, n_4_net__317_, n_4_net__316_, n_4_net__315_, n_4_net__314_, n_4_net__313_, n_4_net__312_, n_4_net__311_, n_4_net__310_, n_4_net__309_, n_4_net__308_, n_4_net__307_, n_4_net__306_, n_4_net__305_, n_4_net__304_, n_4_net__303_, n_4_net__302_, n_4_net__301_, n_4_net__300_, n_4_net__299_, n_4_net__298_, n_4_net__297_, n_4_net__296_, n_4_net__295_, n_4_net__294_, n_4_net__293_, n_4_net__292_, n_4_net__291_, n_4_net__290_, n_4_net__289_, n_4_net__288_, n_4_net__287_, n_4_net__286_, n_4_net__285_, n_4_net__284_, n_4_net__283_, n_4_net__282_, n_4_net__281_, n_4_net__280_, n_4_net__279_, n_4_net__278_, n_4_net__277_, n_4_net__276_, n_4_net__275_, n_4_net__274_, n_4_net__273_, n_4_net__272_, n_4_net__271_, n_4_net__270_, n_4_net__269_, n_4_net__268_, n_4_net__267_, n_4_net__266_, n_4_net__265_, n_4_net__264_, n_4_net__263_, n_4_net__262_, n_4_net__261_, n_4_net__260_, n_4_net__259_, n_4_net__258_, n_4_net__257_, n_4_net__256_, n_4_net__255_, n_4_net__254_, n_4_net__253_, n_4_net__252_, n_4_net__251_, n_4_net__250_, n_4_net__249_, n_4_net__248_, n_4_net__247_, n_4_net__246_, n_4_net__245_, n_4_net__244_, n_4_net__243_, n_4_net__242_, n_4_net__241_, n_4_net__240_, n_4_net__239_, n_4_net__238_, n_4_net__237_, n_4_net__236_, n_4_net__235_, n_4_net__234_, n_4_net__233_, n_4_net__232_, n_4_net__231_, n_4_net__230_, n_4_net__229_, n_4_net__228_, n_4_net__227_, n_4_net__226_, n_4_net__225_, n_4_net__224_, n_4_net__223_, n_4_net__222_, n_4_net__221_, n_4_net__220_, n_4_net__219_, n_4_net__218_, n_4_net__217_, n_4_net__216_, n_4_net__215_, n_4_net__214_, n_4_net__213_, n_4_net__212_, n_4_net__211_, n_4_net__210_, n_4_net__209_, n_4_net__208_, n_4_net__207_, n_4_net__206_, n_4_net__205_, n_4_net__204_, n_4_net__203_, n_4_net__202_, n_4_net__201_, n_4_net__200_, n_4_net__199_, n_4_net__198_, n_4_net__197_, n_4_net__196_, n_4_net__195_, n_4_net__194_, n_4_net__193_, n_4_net__192_, n_4_net__191_, n_4_net__190_, n_4_net__189_, n_4_net__188_, n_4_net__187_, n_4_net__186_, n_4_net__185_, n_4_net__184_, n_4_net__183_, n_4_net__182_, n_4_net__181_, n_4_net__180_, n_4_net__179_, n_4_net__178_, n_4_net__177_, n_4_net__176_, n_4_net__175_, n_4_net__174_, n_4_net__173_, n_4_net__172_, n_4_net__171_, n_4_net__170_, n_4_net__169_, n_4_net__168_, n_4_net__167_, n_4_net__166_, n_4_net__165_, n_4_net__164_, n_4_net__163_, n_4_net__162_, n_4_net__161_, n_4_net__160_, n_4_net__159_, n_4_net__158_, n_4_net__157_, n_4_net__156_, n_4_net__155_, n_4_net__154_, n_4_net__153_, n_4_net__152_, n_4_net__151_, n_4_net__150_, n_4_net__149_, n_4_net__148_, n_4_net__147_, n_4_net__146_, n_4_net__145_, n_4_net__144_, n_4_net__143_, n_4_net__142_, n_4_net__141_, n_4_net__140_, n_4_net__139_, n_4_net__138_, n_4_net__137_, n_4_net__136_, n_4_net__135_, n_4_net__134_, n_4_net__133_, n_4_net__132_, n_4_net__131_, n_4_net__130_, n_4_net__129_, n_4_net__128_, n_4_net__127_, n_4_net__126_, n_4_net__125_, n_4_net__124_, n_4_net__123_, n_4_net__122_, n_4_net__121_, n_4_net__120_, n_4_net__119_, n_4_net__118_, n_4_net__117_, n_4_net__116_, n_4_net__115_, n_4_net__114_, n_4_net__113_, n_4_net__112_, n_4_net__111_, n_4_net__110_, n_4_net__109_, n_4_net__108_, n_4_net__107_, n_4_net__106_, n_4_net__105_, n_4_net__104_, n_4_net__103_, n_4_net__102_, n_4_net__101_, n_4_net__100_, n_4_net__99_, n_4_net__98_, n_4_net__97_, n_4_net__96_, n_4_net__95_, n_4_net__94_, n_4_net__93_, n_4_net__92_, n_4_net__91_, n_4_net__90_, n_4_net__89_, n_4_net__88_, n_4_net__87_, n_4_net__86_, n_4_net__85_, n_4_net__84_, n_4_net__83_, n_4_net__82_, n_4_net__81_, n_4_net__80_, n_4_net__79_, n_4_net__78_, n_4_net__77_, n_4_net__76_, n_4_net__75_, n_4_net__74_, n_4_net__73_, n_4_net__72_, n_4_net__71_, n_4_net__70_, n_4_net__69_, n_4_net__68_, n_4_net__67_, n_4_net__66_, n_4_net__65_, n_4_net__64_, n_4_net__63_, n_4_net__62_, n_4_net__61_, n_4_net__60_, n_4_net__59_, n_4_net__58_, n_4_net__57_, n_4_net__56_, n_4_net__55_, n_4_net__54_, n_4_net__53_, n_4_net__52_, n_4_net__51_, n_4_net__50_, n_4_net__49_, n_4_net__48_, n_4_net__47_, n_4_net__46_, n_4_net__45_, n_4_net__44_, n_4_net__43_, n_4_net__42_, n_4_net__41_, n_4_net__40_, n_4_net__39_, n_4_net__38_, n_4_net__37_, n_4_net__36_, n_4_net__35_, n_4_net__34_, n_4_net__33_, n_4_net__32_, n_4_net__31_, n_4_net__30_, n_4_net__29_, n_4_net__28_, n_4_net__27_, n_4_net__26_, n_4_net__25_, n_4_net__24_, n_4_net__23_, n_4_net__22_, n_4_net__21_, n_4_net__20_, n_4_net__19_, n_4_net__18_, n_4_net__17_, n_4_net__16_, n_4_net__15_, n_4_net__14_, n_4_net__13_, n_4_net__12_, n_4_net__11_, n_4_net__10_, n_4_net__9_, n_4_net__8_, n_4_net__7_, n_4_net__6_, n_4_net__5_, n_4_net__4_, n_4_net__3_, n_4_net__2_, n_4_net__1_, n_4_net__0_ }),
    .o(oc_9__out_chan_data_head_array)
  );


  bsg_rr_f2f_output_width_p64_num_out_p10_middle_meet_p10
  oc_9__out_chan_bsg_rr_ff_out
  (
    .clk(clk),
    .reset(n_5_net_),
    .ready_i(ready_i),
    .ready_head_o({ ready_head_9__9_, ready_head_9__8_, ready_head_9__7_, ready_head_9__6_, ready_head_9__5_, ready_head_9__4_, ready_head_9__3_, ready_head_9__2_, ready_head_9__1_, ready_head_9__0_ }),
    .go_channels_i(go_channels),
    .go_cnt_i(go_cnt),
    .data_head_i(oc_9__out_chan_data_head_array),
    .valid_o({ valid_int_o_9__9_, valid_int_o_9__8_, valid_int_o_9__7_, valid_int_o_9__6_, valid_int_o_9__5_, valid_int_o_9__4_, valid_int_o_9__3_, valid_int_o_9__2_, valid_int_o_9__1_, valid_int_o_9__0_ }),
    .data_o({ data_int_o_9__639_, data_int_o_9__638_, data_int_o_9__637_, data_int_o_9__636_, data_int_o_9__635_, data_int_o_9__634_, data_int_o_9__633_, data_int_o_9__632_, data_int_o_9__631_, data_int_o_9__630_, data_int_o_9__629_, data_int_o_9__628_, data_int_o_9__627_, data_int_o_9__626_, data_int_o_9__625_, data_int_o_9__624_, data_int_o_9__623_, data_int_o_9__622_, data_int_o_9__621_, data_int_o_9__620_, data_int_o_9__619_, data_int_o_9__618_, data_int_o_9__617_, data_int_o_9__616_, data_int_o_9__615_, data_int_o_9__614_, data_int_o_9__613_, data_int_o_9__612_, data_int_o_9__611_, data_int_o_9__610_, data_int_o_9__609_, data_int_o_9__608_, data_int_o_9__607_, data_int_o_9__606_, data_int_o_9__605_, data_int_o_9__604_, data_int_o_9__603_, data_int_o_9__602_, data_int_o_9__601_, data_int_o_9__600_, data_int_o_9__599_, data_int_o_9__598_, data_int_o_9__597_, data_int_o_9__596_, data_int_o_9__595_, data_int_o_9__594_, data_int_o_9__593_, data_int_o_9__592_, data_int_o_9__591_, data_int_o_9__590_, data_int_o_9__589_, data_int_o_9__588_, data_int_o_9__587_, data_int_o_9__586_, data_int_o_9__585_, data_int_o_9__584_, data_int_o_9__583_, data_int_o_9__582_, data_int_o_9__581_, data_int_o_9__580_, data_int_o_9__579_, data_int_o_9__578_, data_int_o_9__577_, data_int_o_9__576_, data_int_o_9__575_, data_int_o_9__574_, data_int_o_9__573_, data_int_o_9__572_, data_int_o_9__571_, data_int_o_9__570_, data_int_o_9__569_, data_int_o_9__568_, data_int_o_9__567_, data_int_o_9__566_, data_int_o_9__565_, data_int_o_9__564_, data_int_o_9__563_, data_int_o_9__562_, data_int_o_9__561_, data_int_o_9__560_, data_int_o_9__559_, data_int_o_9__558_, data_int_o_9__557_, data_int_o_9__556_, data_int_o_9__555_, data_int_o_9__554_, data_int_o_9__553_, data_int_o_9__552_, data_int_o_9__551_, data_int_o_9__550_, data_int_o_9__549_, data_int_o_9__548_, data_int_o_9__547_, data_int_o_9__546_, data_int_o_9__545_, data_int_o_9__544_, data_int_o_9__543_, data_int_o_9__542_, data_int_o_9__541_, data_int_o_9__540_, data_int_o_9__539_, data_int_o_9__538_, data_int_o_9__537_, data_int_o_9__536_, data_int_o_9__535_, data_int_o_9__534_, data_int_o_9__533_, data_int_o_9__532_, data_int_o_9__531_, data_int_o_9__530_, data_int_o_9__529_, data_int_o_9__528_, data_int_o_9__527_, data_int_o_9__526_, data_int_o_9__525_, data_int_o_9__524_, data_int_o_9__523_, data_int_o_9__522_, data_int_o_9__521_, data_int_o_9__520_, data_int_o_9__519_, data_int_o_9__518_, data_int_o_9__517_, data_int_o_9__516_, data_int_o_9__515_, data_int_o_9__514_, data_int_o_9__513_, data_int_o_9__512_, data_int_o_9__511_, data_int_o_9__510_, data_int_o_9__509_, data_int_o_9__508_, data_int_o_9__507_, data_int_o_9__506_, data_int_o_9__505_, data_int_o_9__504_, data_int_o_9__503_, data_int_o_9__502_, data_int_o_9__501_, data_int_o_9__500_, data_int_o_9__499_, data_int_o_9__498_, data_int_o_9__497_, data_int_o_9__496_, data_int_o_9__495_, data_int_o_9__494_, data_int_o_9__493_, data_int_o_9__492_, data_int_o_9__491_, data_int_o_9__490_, data_int_o_9__489_, data_int_o_9__488_, data_int_o_9__487_, data_int_o_9__486_, data_int_o_9__485_, data_int_o_9__484_, data_int_o_9__483_, data_int_o_9__482_, data_int_o_9__481_, data_int_o_9__480_, data_int_o_9__479_, data_int_o_9__478_, data_int_o_9__477_, data_int_o_9__476_, data_int_o_9__475_, data_int_o_9__474_, data_int_o_9__473_, data_int_o_9__472_, data_int_o_9__471_, data_int_o_9__470_, data_int_o_9__469_, data_int_o_9__468_, data_int_o_9__467_, data_int_o_9__466_, data_int_o_9__465_, data_int_o_9__464_, data_int_o_9__463_, data_int_o_9__462_, data_int_o_9__461_, data_int_o_9__460_, data_int_o_9__459_, data_int_o_9__458_, data_int_o_9__457_, data_int_o_9__456_, data_int_o_9__455_, data_int_o_9__454_, data_int_o_9__453_, data_int_o_9__452_, data_int_o_9__451_, data_int_o_9__450_, data_int_o_9__449_, data_int_o_9__448_, data_int_o_9__447_, data_int_o_9__446_, data_int_o_9__445_, data_int_o_9__444_, data_int_o_9__443_, data_int_o_9__442_, data_int_o_9__441_, data_int_o_9__440_, data_int_o_9__439_, data_int_o_9__438_, data_int_o_9__437_, data_int_o_9__436_, data_int_o_9__435_, data_int_o_9__434_, data_int_o_9__433_, data_int_o_9__432_, data_int_o_9__431_, data_int_o_9__430_, data_int_o_9__429_, data_int_o_9__428_, data_int_o_9__427_, data_int_o_9__426_, data_int_o_9__425_, data_int_o_9__424_, data_int_o_9__423_, data_int_o_9__422_, data_int_o_9__421_, data_int_o_9__420_, data_int_o_9__419_, data_int_o_9__418_, data_int_o_9__417_, data_int_o_9__416_, data_int_o_9__415_, data_int_o_9__414_, data_int_o_9__413_, data_int_o_9__412_, data_int_o_9__411_, data_int_o_9__410_, data_int_o_9__409_, data_int_o_9__408_, data_int_o_9__407_, data_int_o_9__406_, data_int_o_9__405_, data_int_o_9__404_, data_int_o_9__403_, data_int_o_9__402_, data_int_o_9__401_, data_int_o_9__400_, data_int_o_9__399_, data_int_o_9__398_, data_int_o_9__397_, data_int_o_9__396_, data_int_o_9__395_, data_int_o_9__394_, data_int_o_9__393_, data_int_o_9__392_, data_int_o_9__391_, data_int_o_9__390_, data_int_o_9__389_, data_int_o_9__388_, data_int_o_9__387_, data_int_o_9__386_, data_int_o_9__385_, data_int_o_9__384_, data_int_o_9__383_, data_int_o_9__382_, data_int_o_9__381_, data_int_o_9__380_, data_int_o_9__379_, data_int_o_9__378_, data_int_o_9__377_, data_int_o_9__376_, data_int_o_9__375_, data_int_o_9__374_, data_int_o_9__373_, data_int_o_9__372_, data_int_o_9__371_, data_int_o_9__370_, data_int_o_9__369_, data_int_o_9__368_, data_int_o_9__367_, data_int_o_9__366_, data_int_o_9__365_, data_int_o_9__364_, data_int_o_9__363_, data_int_o_9__362_, data_int_o_9__361_, data_int_o_9__360_, data_int_o_9__359_, data_int_o_9__358_, data_int_o_9__357_, data_int_o_9__356_, data_int_o_9__355_, data_int_o_9__354_, data_int_o_9__353_, data_int_o_9__352_, data_int_o_9__351_, data_int_o_9__350_, data_int_o_9__349_, data_int_o_9__348_, data_int_o_9__347_, data_int_o_9__346_, data_int_o_9__345_, data_int_o_9__344_, data_int_o_9__343_, data_int_o_9__342_, data_int_o_9__341_, data_int_o_9__340_, data_int_o_9__339_, data_int_o_9__338_, data_int_o_9__337_, data_int_o_9__336_, data_int_o_9__335_, data_int_o_9__334_, data_int_o_9__333_, data_int_o_9__332_, data_int_o_9__331_, data_int_o_9__330_, data_int_o_9__329_, data_int_o_9__328_, data_int_o_9__327_, data_int_o_9__326_, data_int_o_9__325_, data_int_o_9__324_, data_int_o_9__323_, data_int_o_9__322_, data_int_o_9__321_, data_int_o_9__320_, data_int_o_9__319_, data_int_o_9__318_, data_int_o_9__317_, data_int_o_9__316_, data_int_o_9__315_, data_int_o_9__314_, data_int_o_9__313_, data_int_o_9__312_, data_int_o_9__311_, data_int_o_9__310_, data_int_o_9__309_, data_int_o_9__308_, data_int_o_9__307_, data_int_o_9__306_, data_int_o_9__305_, data_int_o_9__304_, data_int_o_9__303_, data_int_o_9__302_, data_int_o_9__301_, data_int_o_9__300_, data_int_o_9__299_, data_int_o_9__298_, data_int_o_9__297_, data_int_o_9__296_, data_int_o_9__295_, data_int_o_9__294_, data_int_o_9__293_, data_int_o_9__292_, data_int_o_9__291_, data_int_o_9__290_, data_int_o_9__289_, data_int_o_9__288_, data_int_o_9__287_, data_int_o_9__286_, data_int_o_9__285_, data_int_o_9__284_, data_int_o_9__283_, data_int_o_9__282_, data_int_o_9__281_, data_int_o_9__280_, data_int_o_9__279_, data_int_o_9__278_, data_int_o_9__277_, data_int_o_9__276_, data_int_o_9__275_, data_int_o_9__274_, data_int_o_9__273_, data_int_o_9__272_, data_int_o_9__271_, data_int_o_9__270_, data_int_o_9__269_, data_int_o_9__268_, data_int_o_9__267_, data_int_o_9__266_, data_int_o_9__265_, data_int_o_9__264_, data_int_o_9__263_, data_int_o_9__262_, data_int_o_9__261_, data_int_o_9__260_, data_int_o_9__259_, data_int_o_9__258_, data_int_o_9__257_, data_int_o_9__256_, data_int_o_9__255_, data_int_o_9__254_, data_int_o_9__253_, data_int_o_9__252_, data_int_o_9__251_, data_int_o_9__250_, data_int_o_9__249_, data_int_o_9__248_, data_int_o_9__247_, data_int_o_9__246_, data_int_o_9__245_, data_int_o_9__244_, data_int_o_9__243_, data_int_o_9__242_, data_int_o_9__241_, data_int_o_9__240_, data_int_o_9__239_, data_int_o_9__238_, data_int_o_9__237_, data_int_o_9__236_, data_int_o_9__235_, data_int_o_9__234_, data_int_o_9__233_, data_int_o_9__232_, data_int_o_9__231_, data_int_o_9__230_, data_int_o_9__229_, data_int_o_9__228_, data_int_o_9__227_, data_int_o_9__226_, data_int_o_9__225_, data_int_o_9__224_, data_int_o_9__223_, data_int_o_9__222_, data_int_o_9__221_, data_int_o_9__220_, data_int_o_9__219_, data_int_o_9__218_, data_int_o_9__217_, data_int_o_9__216_, data_int_o_9__215_, data_int_o_9__214_, data_int_o_9__213_, data_int_o_9__212_, data_int_o_9__211_, data_int_o_9__210_, data_int_o_9__209_, data_int_o_9__208_, data_int_o_9__207_, data_int_o_9__206_, data_int_o_9__205_, data_int_o_9__204_, data_int_o_9__203_, data_int_o_9__202_, data_int_o_9__201_, data_int_o_9__200_, data_int_o_9__199_, data_int_o_9__198_, data_int_o_9__197_, data_int_o_9__196_, data_int_o_9__195_, data_int_o_9__194_, data_int_o_9__193_, data_int_o_9__192_, data_int_o_9__191_, data_int_o_9__190_, data_int_o_9__189_, data_int_o_9__188_, data_int_o_9__187_, data_int_o_9__186_, data_int_o_9__185_, data_int_o_9__184_, data_int_o_9__183_, data_int_o_9__182_, data_int_o_9__181_, data_int_o_9__180_, data_int_o_9__179_, data_int_o_9__178_, data_int_o_9__177_, data_int_o_9__176_, data_int_o_9__175_, data_int_o_9__174_, data_int_o_9__173_, data_int_o_9__172_, data_int_o_9__171_, data_int_o_9__170_, data_int_o_9__169_, data_int_o_9__168_, data_int_o_9__167_, data_int_o_9__166_, data_int_o_9__165_, data_int_o_9__164_, data_int_o_9__163_, data_int_o_9__162_, data_int_o_9__161_, data_int_o_9__160_, data_int_o_9__159_, data_int_o_9__158_, data_int_o_9__157_, data_int_o_9__156_, data_int_o_9__155_, data_int_o_9__154_, data_int_o_9__153_, data_int_o_9__152_, data_int_o_9__151_, data_int_o_9__150_, data_int_o_9__149_, data_int_o_9__148_, data_int_o_9__147_, data_int_o_9__146_, data_int_o_9__145_, data_int_o_9__144_, data_int_o_9__143_, data_int_o_9__142_, data_int_o_9__141_, data_int_o_9__140_, data_int_o_9__139_, data_int_o_9__138_, data_int_o_9__137_, data_int_o_9__136_, data_int_o_9__135_, data_int_o_9__134_, data_int_o_9__133_, data_int_o_9__132_, data_int_o_9__131_, data_int_o_9__130_, data_int_o_9__129_, data_int_o_9__128_, data_int_o_9__127_, data_int_o_9__126_, data_int_o_9__125_, data_int_o_9__124_, data_int_o_9__123_, data_int_o_9__122_, data_int_o_9__121_, data_int_o_9__120_, data_int_o_9__119_, data_int_o_9__118_, data_int_o_9__117_, data_int_o_9__116_, data_int_o_9__115_, data_int_o_9__114_, data_int_o_9__113_, data_int_o_9__112_, data_int_o_9__111_, data_int_o_9__110_, data_int_o_9__109_, data_int_o_9__108_, data_int_o_9__107_, data_int_o_9__106_, data_int_o_9__105_, data_int_o_9__104_, data_int_o_9__103_, data_int_o_9__102_, data_int_o_9__101_, data_int_o_9__100_, data_int_o_9__99_, data_int_o_9__98_, data_int_o_9__97_, data_int_o_9__96_, data_int_o_9__95_, data_int_o_9__94_, data_int_o_9__93_, data_int_o_9__92_, data_int_o_9__91_, data_int_o_9__90_, data_int_o_9__89_, data_int_o_9__88_, data_int_o_9__87_, data_int_o_9__86_, data_int_o_9__85_, data_int_o_9__84_, data_int_o_9__83_, data_int_o_9__82_, data_int_o_9__81_, data_int_o_9__80_, data_int_o_9__79_, data_int_o_9__78_, data_int_o_9__77_, data_int_o_9__76_, data_int_o_9__75_, data_int_o_9__74_, data_int_o_9__73_, data_int_o_9__72_, data_int_o_9__71_, data_int_o_9__70_, data_int_o_9__69_, data_int_o_9__68_, data_int_o_9__67_, data_int_o_9__66_, data_int_o_9__65_, data_int_o_9__64_, data_int_o_9__63_, data_int_o_9__62_, data_int_o_9__61_, data_int_o_9__60_, data_int_o_9__59_, data_int_o_9__58_, data_int_o_9__57_, data_int_o_9__56_, data_int_o_9__55_, data_int_o_9__54_, data_int_o_9__53_, data_int_o_9__52_, data_int_o_9__51_, data_int_o_9__50_, data_int_o_9__49_, data_int_o_9__48_, data_int_o_9__47_, data_int_o_9__46_, data_int_o_9__45_, data_int_o_9__44_, data_int_o_9__43_, data_int_o_9__42_, data_int_o_9__41_, data_int_o_9__40_, data_int_o_9__39_, data_int_o_9__38_, data_int_o_9__37_, data_int_o_9__36_, data_int_o_9__35_, data_int_o_9__34_, data_int_o_9__33_, data_int_o_9__32_, data_int_o_9__31_, data_int_o_9__30_, data_int_o_9__29_, data_int_o_9__28_, data_int_o_9__27_, data_int_o_9__26_, data_int_o_9__25_, data_int_o_9__24_, data_int_o_9__23_, data_int_o_9__22_, data_int_o_9__21_, data_int_o_9__20_, data_int_o_9__19_, data_int_o_9__18_, data_int_o_9__17_, data_int_o_9__16_, data_int_o_9__15_, data_int_o_9__14_, data_int_o_9__13_, data_int_o_9__12_, data_int_o_9__11_, data_int_o_9__10_, data_int_o_9__9_, data_int_o_9__8_, data_int_o_9__7_, data_int_o_9__6_, data_int_o_9__5_, data_int_o_9__4_, data_int_o_9__3_, data_int_o_9__2_, data_int_o_9__1_, data_int_o_9__0_ })
  );

  assign N175 = ~in_top_channel_i[3];
  assign N176 = ~in_top_channel_i[0];
  assign N177 = in_top_channel_i[2] | N175;
  assign N178 = in_top_channel_i[1] | N177;
  assign N179 = N176 | N178;
  assign N180 = ~out_top_channel_i[3];
  assign N181 = ~out_top_channel_i[0];
  assign N182 = out_top_channel_i[2] | N180;
  assign N183 = out_top_channel_i[1] | N182;
  assign N184 = N181 | N183;
  assign N125 = N0 & N1 & (N2 & N3);
  assign N0 = ~in_top_channel_i[3];
  assign N1 = ~in_top_channel_i[2];
  assign N2 = ~in_top_channel_i[0];
  assign N3 = ~in_top_channel_i[1];
  assign N126 = in_top_channel_i[3] & N4;
  assign N4 = ~in_top_channel_i[0];
  assign N127 = N5 & N6 & (in_top_channel_i[0] & N7);
  assign N5 = ~in_top_channel_i[3];
  assign N6 = ~in_top_channel_i[2];
  assign N7 = ~in_top_channel_i[1];
  assign N129 = N8 & N9 & in_top_channel_i[1];
  assign N8 = ~in_top_channel_i[2];
  assign N9 = ~in_top_channel_i[0];
  assign N130 = N10 & in_top_channel_i[0] & in_top_channel_i[1];
  assign N10 = ~in_top_channel_i[2];
  assign N131 = in_top_channel_i[2] & N11 & N12;
  assign N11 = ~in_top_channel_i[0];
  assign N12 = ~in_top_channel_i[1];
  assign N132 = in_top_channel_i[2] & in_top_channel_i[0] & N13;
  assign N13 = ~in_top_channel_i[1];
  assign N133 = in_top_channel_i[2] & N14 & in_top_channel_i[1];
  assign N14 = ~in_top_channel_i[0];
  assign N134 = in_top_channel_i[2] & in_top_channel_i[0] & in_top_channel_i[1];
  assign N128 = in_top_channel_i[3] & in_top_channel_i[0];
  assign N135 = N15 & N16 & (N17 & N18);
  assign N15 = ~out_top_channel_i[3];
  assign N16 = ~out_top_channel_i[2];
  assign N17 = ~out_top_channel_i[0];
  assign N18 = ~out_top_channel_i[1];
  assign N136 = out_top_channel_i[3] & N19;
  assign N19 = ~out_top_channel_i[0];
  assign N137 = N20 & N21 & (out_top_channel_i[0] & N22);
  assign N20 = ~out_top_channel_i[3];
  assign N21 = ~out_top_channel_i[2];
  assign N22 = ~out_top_channel_i[1];
  assign N139 = N23 & N24 & out_top_channel_i[1];
  assign N23 = ~out_top_channel_i[2];
  assign N24 = ~out_top_channel_i[0];
  assign N140 = N25 & out_top_channel_i[0] & out_top_channel_i[1];
  assign N25 = ~out_top_channel_i[2];
  assign N141 = out_top_channel_i[2] & N26 & N27;
  assign N26 = ~out_top_channel_i[0];
  assign N27 = ~out_top_channel_i[1];
  assign N142 = out_top_channel_i[2] & out_top_channel_i[0] & N28;
  assign N28 = ~out_top_channel_i[1];
  assign N143 = out_top_channel_i[2] & N29 & out_top_channel_i[1];
  assign N29 = ~out_top_channel_i[0];
  assign N144 = out_top_channel_i[2] & out_top_channel_i[0] & out_top_channel_i[1];
  assign N138 = out_top_channel_i[3] & out_top_channel_i[0];
  assign N145 = N30 & N31 & (N32 & N33);
  assign N30 = ~out_top_channel_i[3];
  assign N31 = ~out_top_channel_i[2];
  assign N32 = ~out_top_channel_i[0];
  assign N33 = ~out_top_channel_i[1];
  assign N146 = out_top_channel_i[3] & N34;
  assign N34 = ~out_top_channel_i[0];
  assign N147 = N35 & N36 & (out_top_channel_i[0] & N37);
  assign N35 = ~out_top_channel_i[3];
  assign N36 = ~out_top_channel_i[2];
  assign N37 = ~out_top_channel_i[1];
  assign N149 = N38 & N39 & out_top_channel_i[1];
  assign N38 = ~out_top_channel_i[2];
  assign N39 = ~out_top_channel_i[0];
  assign N150 = N40 & out_top_channel_i[0] & out_top_channel_i[1];
  assign N40 = ~out_top_channel_i[2];
  assign N151 = out_top_channel_i[2] & N41 & N42;
  assign N41 = ~out_top_channel_i[0];
  assign N42 = ~out_top_channel_i[1];
  assign N152 = out_top_channel_i[2] & out_top_channel_i[0] & N43;
  assign N43 = ~out_top_channel_i[1];
  assign N153 = out_top_channel_i[2] & N44 & out_top_channel_i[1];
  assign N44 = ~out_top_channel_i[0];
  assign N154 = out_top_channel_i[2] & out_top_channel_i[0] & out_top_channel_i[1];
  assign N148 = out_top_channel_i[3] & out_top_channel_i[0];
  assign N155 = N45 & N46 & (N47 & N48);
  assign N45 = ~in_top_channel_i[3];
  assign N46 = ~in_top_channel_i[2];
  assign N47 = ~in_top_channel_i[0];
  assign N48 = ~in_top_channel_i[1];
  assign N156 = in_top_channel_i[3] & N49;
  assign N49 = ~in_top_channel_i[0];
  assign N157 = N50 & N51 & (in_top_channel_i[0] & N52);
  assign N50 = ~in_top_channel_i[3];
  assign N51 = ~in_top_channel_i[2];
  assign N52 = ~in_top_channel_i[1];
  assign N159 = N53 & N54 & in_top_channel_i[1];
  assign N53 = ~in_top_channel_i[2];
  assign N54 = ~in_top_channel_i[0];
  assign N160 = N55 & in_top_channel_i[0] & in_top_channel_i[1];
  assign N55 = ~in_top_channel_i[2];
  assign N161 = in_top_channel_i[2] & N56 & N57;
  assign N56 = ~in_top_channel_i[0];
  assign N57 = ~in_top_channel_i[1];
  assign N162 = in_top_channel_i[2] & in_top_channel_i[0] & N58;
  assign N58 = ~in_top_channel_i[1];
  assign N163 = in_top_channel_i[2] & N59 & in_top_channel_i[1];
  assign N59 = ~in_top_channel_i[0];
  assign N164 = in_top_channel_i[2] & in_top_channel_i[0] & in_top_channel_i[1];
  assign N158 = in_top_channel_i[3] & in_top_channel_i[0];
  assign N165 = N60 & N61 & (N62 & N63);
  assign N60 = ~in_top_channel_i[3];
  assign N61 = ~in_top_channel_i[2];
  assign N62 = ~in_top_channel_i[0];
  assign N63 = ~in_top_channel_i[1];
  assign N166 = in_top_channel_i[3] & N64;
  assign N64 = ~in_top_channel_i[0];
  assign N167 = N65 & N66 & (in_top_channel_i[0] & N67);
  assign N65 = ~in_top_channel_i[3];
  assign N66 = ~in_top_channel_i[2];
  assign N67 = ~in_top_channel_i[1];
  assign N169 = N68 & N69 & in_top_channel_i[1];
  assign N68 = ~in_top_channel_i[2];
  assign N69 = ~in_top_channel_i[0];
  assign N170 = N70 & in_top_channel_i[0] & in_top_channel_i[1];
  assign N70 = ~in_top_channel_i[2];
  assign N171 = in_top_channel_i[2] & N71 & N72;
  assign N71 = ~in_top_channel_i[0];
  assign N72 = ~in_top_channel_i[1];
  assign N172 = in_top_channel_i[2] & in_top_channel_i[0] & N73;
  assign N73 = ~in_top_channel_i[1];
  assign N173 = in_top_channel_i[2] & N74 & in_top_channel_i[1];
  assign N74 = ~in_top_channel_i[0];
  assign N174 = in_top_channel_i[2] & in_top_channel_i[0] & in_top_channel_i[1];
  assign N168 = in_top_channel_i[3] & in_top_channel_i[0];
  assign yumi_o[9] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__9_ : 1'b0;
  assign N75 = N125;
  assign N76 = N127;
  assign N77 = N129;
  assign N78 = N130;
  assign N79 = N131;
  assign N80 = N132;
  assign N81 = N133;
  assign N82 = N134;
  assign N83 = N126;
  assign N84 = N128;
  assign yumi_o[8] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__8_ : 1'b0;
  assign yumi_o[7] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__7_ : 1'b0;
  assign yumi_o[6] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__6_ : 1'b0;
  assign yumi_o[5] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__5_ : 1'b0;
  assign yumi_o[4] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__4_ : 1'b0;
  assign yumi_o[3] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__3_ : 1'b0;
  assign yumi_o[2] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__2_ : 1'b0;
  assign yumi_o[1] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__1_ : 1'b0;
  assign yumi_o[0] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__0_ : 1'b0;
  assign valid_o[9] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__9_ : 1'b0;
  assign N85 = N135;
  assign N86 = N137;
  assign N87 = N139;
  assign N88 = N140;
  assign N89 = N141;
  assign N90 = N142;
  assign N91 = N143;
  assign N92 = N144;
  assign N93 = N136;
  assign N94 = N138;
  assign valid_o[8] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__8_ : 1'b0;
  assign valid_o[7] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__7_ : 1'b0;
  assign valid_o[6] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__6_ : 1'b0;
  assign valid_o[5] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__5_ : 1'b0;
  assign valid_o[4] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__4_ : 1'b0;
  assign valid_o[3] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__3_ : 1'b0;
  assign valid_o[2] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__2_ : 1'b0;
  assign valid_o[1] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__1_ : 1'b0;
  assign valid_o[0] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__0_ : 1'b0;
  assign data_o_flat[639] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__639_ : 1'b0;
  assign N95 = N145;
  assign N96 = N147;
  assign N97 = N149;
  assign N98 = N150;
  assign N99 = N151;
  assign N100 = N152;
  assign N101 = N153;
  assign N102 = N154;
  assign N103 = N146;
  assign N104 = N148;
  assign data_o_flat[638] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__638_ : 1'b0;
  assign data_o_flat[637] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__637_ : 1'b0;
  assign data_o_flat[636] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__636_ : 1'b0;
  assign data_o_flat[635] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__635_ : 1'b0;
  assign data_o_flat[634] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__634_ : 1'b0;
  assign data_o_flat[633] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__633_ : 1'b0;
  assign data_o_flat[632] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__632_ : 1'b0;
  assign data_o_flat[631] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__631_ : 1'b0;
  assign data_o_flat[630] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__630_ : 1'b0;
  assign data_o_flat[629] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__629_ : 1'b0;
  assign data_o_flat[628] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__628_ : 1'b0;
  assign data_o_flat[627] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__627_ : 1'b0;
  assign data_o_flat[626] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__626_ : 1'b0;
  assign data_o_flat[625] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__625_ : 1'b0;
  assign data_o_flat[624] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__624_ : 1'b0;
  assign data_o_flat[623] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__623_ : 1'b0;
  assign data_o_flat[622] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__622_ : 1'b0;
  assign data_o_flat[621] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__621_ : 1'b0;
  assign data_o_flat[620] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__620_ : 1'b0;
  assign data_o_flat[619] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__619_ : 1'b0;
  assign data_o_flat[618] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__618_ : 1'b0;
  assign data_o_flat[617] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__617_ : 1'b0;
  assign data_o_flat[616] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__616_ : 1'b0;
  assign data_o_flat[615] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__615_ : 1'b0;
  assign data_o_flat[614] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__614_ : 1'b0;
  assign data_o_flat[613] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__613_ : 1'b0;
  assign data_o_flat[612] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__612_ : 1'b0;
  assign data_o_flat[611] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__611_ : 1'b0;
  assign data_o_flat[610] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__610_ : 1'b0;
  assign data_o_flat[609] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__609_ : 1'b0;
  assign data_o_flat[608] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__608_ : 1'b0;
  assign data_o_flat[607] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__607_ : 1'b0;
  assign data_o_flat[606] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__606_ : 1'b0;
  assign data_o_flat[605] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__605_ : 1'b0;
  assign data_o_flat[604] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__604_ : 1'b0;
  assign data_o_flat[603] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__603_ : 1'b0;
  assign data_o_flat[602] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__602_ : 1'b0;
  assign data_o_flat[601] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__601_ : 1'b0;
  assign data_o_flat[600] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__600_ : 1'b0;
  assign data_o_flat[599] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__599_ : 1'b0;
  assign data_o_flat[598] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__598_ : 1'b0;
  assign data_o_flat[597] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__597_ : 1'b0;
  assign data_o_flat[596] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__596_ : 1'b0;
  assign data_o_flat[595] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__595_ : 1'b0;
  assign data_o_flat[594] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__594_ : 1'b0;
  assign data_o_flat[593] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__593_ : 1'b0;
  assign data_o_flat[592] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__592_ : 1'b0;
  assign data_o_flat[591] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__591_ : 1'b0;
  assign data_o_flat[590] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__590_ : 1'b0;
  assign data_o_flat[589] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__589_ : 1'b0;
  assign data_o_flat[588] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__588_ : 1'b0;
  assign data_o_flat[587] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__587_ : 1'b0;
  assign data_o_flat[586] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__586_ : 1'b0;
  assign data_o_flat[585] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__585_ : 1'b0;
  assign data_o_flat[584] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__584_ : 1'b0;
  assign data_o_flat[583] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__583_ : 1'b0;
  assign data_o_flat[582] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__582_ : 1'b0;
  assign data_o_flat[581] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__581_ : 1'b0;
  assign data_o_flat[580] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__580_ : 1'b0;
  assign data_o_flat[579] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__579_ : 1'b0;
  assign data_o_flat[578] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__578_ : 1'b0;
  assign data_o_flat[577] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__577_ : 1'b0;
  assign data_o_flat[576] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__576_ : 1'b0;
  assign data_o_flat[575] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__575_ : 1'b0;
  assign data_o_flat[574] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__574_ : 1'b0;
  assign data_o_flat[573] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__573_ : 1'b0;
  assign data_o_flat[572] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__572_ : 1'b0;
  assign data_o_flat[571] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__571_ : 1'b0;
  assign data_o_flat[570] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__570_ : 1'b0;
  assign data_o_flat[569] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__569_ : 1'b0;
  assign data_o_flat[568] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__568_ : 1'b0;
  assign data_o_flat[567] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__567_ : 1'b0;
  assign data_o_flat[566] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__566_ : 1'b0;
  assign data_o_flat[565] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__565_ : 1'b0;
  assign data_o_flat[564] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__564_ : 1'b0;
  assign data_o_flat[563] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__563_ : 1'b0;
  assign data_o_flat[562] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__562_ : 1'b0;
  assign data_o_flat[561] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__561_ : 1'b0;
  assign data_o_flat[560] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__560_ : 1'b0;
  assign data_o_flat[559] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__559_ : 1'b0;
  assign data_o_flat[558] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__558_ : 1'b0;
  assign data_o_flat[557] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__557_ : 1'b0;
  assign data_o_flat[556] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__556_ : 1'b0;
  assign data_o_flat[555] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__555_ : 1'b0;
  assign data_o_flat[554] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__554_ : 1'b0;
  assign data_o_flat[553] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__553_ : 1'b0;
  assign data_o_flat[552] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__552_ : 1'b0;
  assign data_o_flat[551] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__551_ : 1'b0;
  assign data_o_flat[550] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__550_ : 1'b0;
  assign data_o_flat[549] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__549_ : 1'b0;
  assign data_o_flat[548] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__548_ : 1'b0;
  assign data_o_flat[547] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__547_ : 1'b0;
  assign data_o_flat[546] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__546_ : 1'b0;
  assign data_o_flat[545] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__545_ : 1'b0;
  assign data_o_flat[544] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__544_ : 1'b0;
  assign data_o_flat[543] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__543_ : 1'b0;
  assign data_o_flat[542] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__542_ : 1'b0;
  assign data_o_flat[541] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__541_ : 1'b0;
  assign data_o_flat[540] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__540_ : 1'b0;
  assign data_o_flat[539] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__539_ : 1'b0;
  assign data_o_flat[538] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__538_ : 1'b0;
  assign data_o_flat[537] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__537_ : 1'b0;
  assign data_o_flat[536] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__536_ : 1'b0;
  assign data_o_flat[535] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__535_ : 1'b0;
  assign data_o_flat[534] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__534_ : 1'b0;
  assign data_o_flat[533] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__533_ : 1'b0;
  assign data_o_flat[532] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__532_ : 1'b0;
  assign data_o_flat[531] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__531_ : 1'b0;
  assign data_o_flat[530] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__530_ : 1'b0;
  assign data_o_flat[529] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__529_ : 1'b0;
  assign data_o_flat[528] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__528_ : 1'b0;
  assign data_o_flat[527] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__527_ : 1'b0;
  assign data_o_flat[526] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__526_ : 1'b0;
  assign data_o_flat[525] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__525_ : 1'b0;
  assign data_o_flat[524] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__524_ : 1'b0;
  assign data_o_flat[523] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__523_ : 1'b0;
  assign data_o_flat[522] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__522_ : 1'b0;
  assign data_o_flat[521] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__521_ : 1'b0;
  assign data_o_flat[520] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__520_ : 1'b0;
  assign data_o_flat[519] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__519_ : 1'b0;
  assign data_o_flat[518] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__518_ : 1'b0;
  assign data_o_flat[517] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__517_ : 1'b0;
  assign data_o_flat[516] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__516_ : 1'b0;
  assign data_o_flat[515] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__515_ : 1'b0;
  assign data_o_flat[514] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__514_ : 1'b0;
  assign data_o_flat[513] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__513_ : 1'b0;
  assign data_o_flat[512] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__512_ : 1'b0;
  assign data_o_flat[511] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__511_ : 1'b0;
  assign data_o_flat[510] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__510_ : 1'b0;
  assign data_o_flat[509] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__509_ : 1'b0;
  assign data_o_flat[508] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__508_ : 1'b0;
  assign data_o_flat[507] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__507_ : 1'b0;
  assign data_o_flat[506] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__506_ : 1'b0;
  assign data_o_flat[505] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__505_ : 1'b0;
  assign data_o_flat[504] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__504_ : 1'b0;
  assign data_o_flat[503] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__503_ : 1'b0;
  assign data_o_flat[502] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__502_ : 1'b0;
  assign data_o_flat[501] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__501_ : 1'b0;
  assign data_o_flat[500] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__500_ : 1'b0;
  assign data_o_flat[499] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__499_ : 1'b0;
  assign data_o_flat[498] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__498_ : 1'b0;
  assign data_o_flat[497] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__497_ : 1'b0;
  assign data_o_flat[496] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__496_ : 1'b0;
  assign data_o_flat[495] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__495_ : 1'b0;
  assign data_o_flat[494] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__494_ : 1'b0;
  assign data_o_flat[493] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__493_ : 1'b0;
  assign data_o_flat[492] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__492_ : 1'b0;
  assign data_o_flat[491] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__491_ : 1'b0;
  assign data_o_flat[490] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__490_ : 1'b0;
  assign data_o_flat[489] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__489_ : 1'b0;
  assign data_o_flat[488] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__488_ : 1'b0;
  assign data_o_flat[487] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__487_ : 1'b0;
  assign data_o_flat[486] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__486_ : 1'b0;
  assign data_o_flat[485] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__485_ : 1'b0;
  assign data_o_flat[484] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__484_ : 1'b0;
  assign data_o_flat[483] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__483_ : 1'b0;
  assign data_o_flat[482] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__482_ : 1'b0;
  assign data_o_flat[481] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__481_ : 1'b0;
  assign data_o_flat[480] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__480_ : 1'b0;
  assign data_o_flat[479] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__479_ : 1'b0;
  assign data_o_flat[478] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__478_ : 1'b0;
  assign data_o_flat[477] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__477_ : 1'b0;
  assign data_o_flat[476] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__476_ : 1'b0;
  assign data_o_flat[475] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__475_ : 1'b0;
  assign data_o_flat[474] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__474_ : 1'b0;
  assign data_o_flat[473] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__473_ : 1'b0;
  assign data_o_flat[472] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__472_ : 1'b0;
  assign data_o_flat[471] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__471_ : 1'b0;
  assign data_o_flat[470] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__470_ : 1'b0;
  assign data_o_flat[469] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__469_ : 1'b0;
  assign data_o_flat[468] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__468_ : 1'b0;
  assign data_o_flat[467] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__467_ : 1'b0;
  assign data_o_flat[466] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__466_ : 1'b0;
  assign data_o_flat[465] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__465_ : 1'b0;
  assign data_o_flat[464] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__464_ : 1'b0;
  assign data_o_flat[463] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__463_ : 1'b0;
  assign data_o_flat[462] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__462_ : 1'b0;
  assign data_o_flat[461] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__461_ : 1'b0;
  assign data_o_flat[460] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__460_ : 1'b0;
  assign data_o_flat[459] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__459_ : 1'b0;
  assign data_o_flat[458] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__458_ : 1'b0;
  assign data_o_flat[457] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__457_ : 1'b0;
  assign data_o_flat[456] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__456_ : 1'b0;
  assign data_o_flat[455] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__455_ : 1'b0;
  assign data_o_flat[454] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__454_ : 1'b0;
  assign data_o_flat[453] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__453_ : 1'b0;
  assign data_o_flat[452] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__452_ : 1'b0;
  assign data_o_flat[451] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__451_ : 1'b0;
  assign data_o_flat[450] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__450_ : 1'b0;
  assign data_o_flat[449] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__449_ : 1'b0;
  assign data_o_flat[448] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__448_ : 1'b0;
  assign data_o_flat[447] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__447_ : 1'b0;
  assign data_o_flat[446] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__446_ : 1'b0;
  assign data_o_flat[445] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__445_ : 1'b0;
  assign data_o_flat[444] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__444_ : 1'b0;
  assign data_o_flat[443] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__443_ : 1'b0;
  assign data_o_flat[442] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__442_ : 1'b0;
  assign data_o_flat[441] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__441_ : 1'b0;
  assign data_o_flat[440] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__440_ : 1'b0;
  assign data_o_flat[439] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__439_ : 1'b0;
  assign data_o_flat[438] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__438_ : 1'b0;
  assign data_o_flat[437] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__437_ : 1'b0;
  assign data_o_flat[436] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__436_ : 1'b0;
  assign data_o_flat[435] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__435_ : 1'b0;
  assign data_o_flat[434] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__434_ : 1'b0;
  assign data_o_flat[433] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__433_ : 1'b0;
  assign data_o_flat[432] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__432_ : 1'b0;
  assign data_o_flat[431] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__431_ : 1'b0;
  assign data_o_flat[430] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__430_ : 1'b0;
  assign data_o_flat[429] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__429_ : 1'b0;
  assign data_o_flat[428] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__428_ : 1'b0;
  assign data_o_flat[427] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__427_ : 1'b0;
  assign data_o_flat[426] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__426_ : 1'b0;
  assign data_o_flat[425] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__425_ : 1'b0;
  assign data_o_flat[424] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__424_ : 1'b0;
  assign data_o_flat[423] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__423_ : 1'b0;
  assign data_o_flat[422] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__422_ : 1'b0;
  assign data_o_flat[421] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__421_ : 1'b0;
  assign data_o_flat[420] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__420_ : 1'b0;
  assign data_o_flat[419] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__419_ : 1'b0;
  assign data_o_flat[418] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__418_ : 1'b0;
  assign data_o_flat[417] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__417_ : 1'b0;
  assign data_o_flat[416] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__416_ : 1'b0;
  assign data_o_flat[415] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__415_ : 1'b0;
  assign data_o_flat[414] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__414_ : 1'b0;
  assign data_o_flat[413] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__413_ : 1'b0;
  assign data_o_flat[412] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__412_ : 1'b0;
  assign data_o_flat[411] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__411_ : 1'b0;
  assign data_o_flat[410] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__410_ : 1'b0;
  assign data_o_flat[409] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__409_ : 1'b0;
  assign data_o_flat[408] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__408_ : 1'b0;
  assign data_o_flat[407] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__407_ : 1'b0;
  assign data_o_flat[406] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__406_ : 1'b0;
  assign data_o_flat[405] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__405_ : 1'b0;
  assign data_o_flat[404] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__404_ : 1'b0;
  assign data_o_flat[403] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__403_ : 1'b0;
  assign data_o_flat[402] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__402_ : 1'b0;
  assign data_o_flat[401] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__401_ : 1'b0;
  assign data_o_flat[400] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__400_ : 1'b0;
  assign data_o_flat[399] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__399_ : 1'b0;
  assign data_o_flat[398] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__398_ : 1'b0;
  assign data_o_flat[397] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__397_ : 1'b0;
  assign data_o_flat[396] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__396_ : 1'b0;
  assign data_o_flat[395] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__395_ : 1'b0;
  assign data_o_flat[394] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__394_ : 1'b0;
  assign data_o_flat[393] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__393_ : 1'b0;
  assign data_o_flat[392] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__392_ : 1'b0;
  assign data_o_flat[391] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__391_ : 1'b0;
  assign data_o_flat[390] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__390_ : 1'b0;
  assign data_o_flat[389] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__389_ : 1'b0;
  assign data_o_flat[388] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__388_ : 1'b0;
  assign data_o_flat[387] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__387_ : 1'b0;
  assign data_o_flat[386] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__386_ : 1'b0;
  assign data_o_flat[385] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__385_ : 1'b0;
  assign data_o_flat[384] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__384_ : 1'b0;
  assign data_o_flat[383] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__383_ : 1'b0;
  assign data_o_flat[382] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__382_ : 1'b0;
  assign data_o_flat[381] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__381_ : 1'b0;
  assign data_o_flat[380] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__380_ : 1'b0;
  assign data_o_flat[379] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__379_ : 1'b0;
  assign data_o_flat[378] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__378_ : 1'b0;
  assign data_o_flat[377] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__377_ : 1'b0;
  assign data_o_flat[376] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__376_ : 1'b0;
  assign data_o_flat[375] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__375_ : 1'b0;
  assign data_o_flat[374] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__374_ : 1'b0;
  assign data_o_flat[373] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__373_ : 1'b0;
  assign data_o_flat[372] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__372_ : 1'b0;
  assign data_o_flat[371] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__371_ : 1'b0;
  assign data_o_flat[370] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__370_ : 1'b0;
  assign data_o_flat[369] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__369_ : 1'b0;
  assign data_o_flat[368] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__368_ : 1'b0;
  assign data_o_flat[367] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__367_ : 1'b0;
  assign data_o_flat[366] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__366_ : 1'b0;
  assign data_o_flat[365] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__365_ : 1'b0;
  assign data_o_flat[364] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__364_ : 1'b0;
  assign data_o_flat[363] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__363_ : 1'b0;
  assign data_o_flat[362] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__362_ : 1'b0;
  assign data_o_flat[361] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__361_ : 1'b0;
  assign data_o_flat[360] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__360_ : 1'b0;
  assign data_o_flat[359] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__359_ : 1'b0;
  assign data_o_flat[358] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__358_ : 1'b0;
  assign data_o_flat[357] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__357_ : 1'b0;
  assign data_o_flat[356] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__356_ : 1'b0;
  assign data_o_flat[355] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__355_ : 1'b0;
  assign data_o_flat[354] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__354_ : 1'b0;
  assign data_o_flat[353] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__353_ : 1'b0;
  assign data_o_flat[352] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__352_ : 1'b0;
  assign data_o_flat[351] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__351_ : 1'b0;
  assign data_o_flat[350] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__350_ : 1'b0;
  assign data_o_flat[349] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__349_ : 1'b0;
  assign data_o_flat[348] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__348_ : 1'b0;
  assign data_o_flat[347] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__347_ : 1'b0;
  assign data_o_flat[346] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__346_ : 1'b0;
  assign data_o_flat[345] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__345_ : 1'b0;
  assign data_o_flat[344] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__344_ : 1'b0;
  assign data_o_flat[343] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__343_ : 1'b0;
  assign data_o_flat[342] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__342_ : 1'b0;
  assign data_o_flat[341] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__341_ : 1'b0;
  assign data_o_flat[340] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__340_ : 1'b0;
  assign data_o_flat[339] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__339_ : 1'b0;
  assign data_o_flat[338] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__338_ : 1'b0;
  assign data_o_flat[337] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__337_ : 1'b0;
  assign data_o_flat[336] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__336_ : 1'b0;
  assign data_o_flat[335] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__335_ : 1'b0;
  assign data_o_flat[334] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__334_ : 1'b0;
  assign data_o_flat[333] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__333_ : 1'b0;
  assign data_o_flat[332] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__332_ : 1'b0;
  assign data_o_flat[331] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__331_ : 1'b0;
  assign data_o_flat[330] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__330_ : 1'b0;
  assign data_o_flat[329] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__329_ : 1'b0;
  assign data_o_flat[328] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__328_ : 1'b0;
  assign data_o_flat[327] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__327_ : 1'b0;
  assign data_o_flat[326] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__326_ : 1'b0;
  assign data_o_flat[325] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__325_ : 1'b0;
  assign data_o_flat[324] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__324_ : 1'b0;
  assign data_o_flat[323] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__323_ : 1'b0;
  assign data_o_flat[322] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__322_ : 1'b0;
  assign data_o_flat[321] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__321_ : 1'b0;
  assign data_o_flat[320] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__320_ : 1'b0;
  assign data_o_flat[319] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__319_ : 1'b0;
  assign data_o_flat[318] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__318_ : 1'b0;
  assign data_o_flat[317] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__317_ : 1'b0;
  assign data_o_flat[316] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__316_ : 1'b0;
  assign data_o_flat[315] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__315_ : 1'b0;
  assign data_o_flat[314] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__314_ : 1'b0;
  assign data_o_flat[313] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__313_ : 1'b0;
  assign data_o_flat[312] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__312_ : 1'b0;
  assign data_o_flat[311] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__311_ : 1'b0;
  assign data_o_flat[310] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__310_ : 1'b0;
  assign data_o_flat[309] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__309_ : 1'b0;
  assign data_o_flat[308] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__308_ : 1'b0;
  assign data_o_flat[307] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__307_ : 1'b0;
  assign data_o_flat[306] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__306_ : 1'b0;
  assign data_o_flat[305] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__305_ : 1'b0;
  assign data_o_flat[304] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__304_ : 1'b0;
  assign data_o_flat[303] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__303_ : 1'b0;
  assign data_o_flat[302] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__302_ : 1'b0;
  assign data_o_flat[301] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__301_ : 1'b0;
  assign data_o_flat[300] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__300_ : 1'b0;
  assign data_o_flat[299] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__299_ : 1'b0;
  assign data_o_flat[298] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__298_ : 1'b0;
  assign data_o_flat[297] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__297_ : 1'b0;
  assign data_o_flat[296] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__296_ : 1'b0;
  assign data_o_flat[295] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__295_ : 1'b0;
  assign data_o_flat[294] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__294_ : 1'b0;
  assign data_o_flat[293] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__293_ : 1'b0;
  assign data_o_flat[292] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__292_ : 1'b0;
  assign data_o_flat[291] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__291_ : 1'b0;
  assign data_o_flat[290] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__290_ : 1'b0;
  assign data_o_flat[289] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__289_ : 1'b0;
  assign data_o_flat[288] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__288_ : 1'b0;
  assign data_o_flat[287] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__287_ : 1'b0;
  assign data_o_flat[286] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__286_ : 1'b0;
  assign data_o_flat[285] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__285_ : 1'b0;
  assign data_o_flat[284] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__284_ : 1'b0;
  assign data_o_flat[283] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__283_ : 1'b0;
  assign data_o_flat[282] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__282_ : 1'b0;
  assign data_o_flat[281] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__281_ : 1'b0;
  assign data_o_flat[280] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__280_ : 1'b0;
  assign data_o_flat[279] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__279_ : 1'b0;
  assign data_o_flat[278] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__278_ : 1'b0;
  assign data_o_flat[277] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__277_ : 1'b0;
  assign data_o_flat[276] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__276_ : 1'b0;
  assign data_o_flat[275] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__275_ : 1'b0;
  assign data_o_flat[274] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__274_ : 1'b0;
  assign data_o_flat[273] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__273_ : 1'b0;
  assign data_o_flat[272] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__272_ : 1'b0;
  assign data_o_flat[271] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__271_ : 1'b0;
  assign data_o_flat[270] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__270_ : 1'b0;
  assign data_o_flat[269] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__269_ : 1'b0;
  assign data_o_flat[268] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__268_ : 1'b0;
  assign data_o_flat[267] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__267_ : 1'b0;
  assign data_o_flat[266] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__266_ : 1'b0;
  assign data_o_flat[265] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__265_ : 1'b0;
  assign data_o_flat[264] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__264_ : 1'b0;
  assign data_o_flat[263] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__263_ : 1'b0;
  assign data_o_flat[262] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__262_ : 1'b0;
  assign data_o_flat[261] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__261_ : 1'b0;
  assign data_o_flat[260] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__260_ : 1'b0;
  assign data_o_flat[259] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__259_ : 1'b0;
  assign data_o_flat[258] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__258_ : 1'b0;
  assign data_o_flat[257] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__257_ : 1'b0;
  assign data_o_flat[256] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__256_ : 1'b0;
  assign data_o_flat[255] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__255_ : 1'b0;
  assign data_o_flat[254] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__254_ : 1'b0;
  assign data_o_flat[253] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__253_ : 1'b0;
  assign data_o_flat[252] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__252_ : 1'b0;
  assign data_o_flat[251] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__251_ : 1'b0;
  assign data_o_flat[250] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__250_ : 1'b0;
  assign data_o_flat[249] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__249_ : 1'b0;
  assign data_o_flat[248] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__248_ : 1'b0;
  assign data_o_flat[247] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__247_ : 1'b0;
  assign data_o_flat[246] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__246_ : 1'b0;
  assign data_o_flat[245] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__245_ : 1'b0;
  assign data_o_flat[244] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__244_ : 1'b0;
  assign data_o_flat[243] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__243_ : 1'b0;
  assign data_o_flat[242] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__242_ : 1'b0;
  assign data_o_flat[241] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__241_ : 1'b0;
  assign data_o_flat[240] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__240_ : 1'b0;
  assign data_o_flat[239] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__239_ : 1'b0;
  assign data_o_flat[238] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__238_ : 1'b0;
  assign data_o_flat[237] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__237_ : 1'b0;
  assign data_o_flat[236] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__236_ : 1'b0;
  assign data_o_flat[235] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__235_ : 1'b0;
  assign data_o_flat[234] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__234_ : 1'b0;
  assign data_o_flat[233] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__233_ : 1'b0;
  assign data_o_flat[232] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__232_ : 1'b0;
  assign data_o_flat[231] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__231_ : 1'b0;
  assign data_o_flat[230] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__230_ : 1'b0;
  assign data_o_flat[229] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__229_ : 1'b0;
  assign data_o_flat[228] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__228_ : 1'b0;
  assign data_o_flat[227] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__227_ : 1'b0;
  assign data_o_flat[226] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__226_ : 1'b0;
  assign data_o_flat[225] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__225_ : 1'b0;
  assign data_o_flat[224] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__224_ : 1'b0;
  assign data_o_flat[223] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__223_ : 1'b0;
  assign data_o_flat[222] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__222_ : 1'b0;
  assign data_o_flat[221] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__221_ : 1'b0;
  assign data_o_flat[220] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__220_ : 1'b0;
  assign data_o_flat[219] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__219_ : 1'b0;
  assign data_o_flat[218] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__218_ : 1'b0;
  assign data_o_flat[217] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__217_ : 1'b0;
  assign data_o_flat[216] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__216_ : 1'b0;
  assign data_o_flat[215] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__215_ : 1'b0;
  assign data_o_flat[214] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__214_ : 1'b0;
  assign data_o_flat[213] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__213_ : 1'b0;
  assign data_o_flat[212] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__212_ : 1'b0;
  assign data_o_flat[211] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__211_ : 1'b0;
  assign data_o_flat[210] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__210_ : 1'b0;
  assign data_o_flat[209] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__209_ : 1'b0;
  assign data_o_flat[208] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__208_ : 1'b0;
  assign data_o_flat[207] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__207_ : 1'b0;
  assign data_o_flat[206] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__206_ : 1'b0;
  assign data_o_flat[205] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__205_ : 1'b0;
  assign data_o_flat[204] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__204_ : 1'b0;
  assign data_o_flat[203] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__203_ : 1'b0;
  assign data_o_flat[202] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__202_ : 1'b0;
  assign data_o_flat[201] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__201_ : 1'b0;
  assign data_o_flat[200] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__200_ : 1'b0;
  assign data_o_flat[199] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__199_ : 1'b0;
  assign data_o_flat[198] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__198_ : 1'b0;
  assign data_o_flat[197] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__197_ : 1'b0;
  assign data_o_flat[196] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__196_ : 1'b0;
  assign data_o_flat[195] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__195_ : 1'b0;
  assign data_o_flat[194] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__194_ : 1'b0;
  assign data_o_flat[193] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__193_ : 1'b0;
  assign data_o_flat[192] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__192_ : 1'b0;
  assign data_o_flat[191] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__191_ : 1'b0;
  assign data_o_flat[190] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__190_ : 1'b0;
  assign data_o_flat[189] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__189_ : 1'b0;
  assign data_o_flat[188] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__188_ : 1'b0;
  assign data_o_flat[187] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__187_ : 1'b0;
  assign data_o_flat[186] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__186_ : 1'b0;
  assign data_o_flat[185] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__185_ : 1'b0;
  assign data_o_flat[184] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__184_ : 1'b0;
  assign data_o_flat[183] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__183_ : 1'b0;
  assign data_o_flat[182] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__182_ : 1'b0;
  assign data_o_flat[181] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__181_ : 1'b0;
  assign data_o_flat[180] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__180_ : 1'b0;
  assign data_o_flat[179] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__179_ : 1'b0;
  assign data_o_flat[178] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__178_ : 1'b0;
  assign data_o_flat[177] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__177_ : 1'b0;
  assign data_o_flat[176] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__176_ : 1'b0;
  assign data_o_flat[175] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__175_ : 1'b0;
  assign data_o_flat[174] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__174_ : 1'b0;
  assign data_o_flat[173] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__173_ : 1'b0;
  assign data_o_flat[172] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__172_ : 1'b0;
  assign data_o_flat[171] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__171_ : 1'b0;
  assign data_o_flat[170] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__170_ : 1'b0;
  assign data_o_flat[169] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__169_ : 1'b0;
  assign data_o_flat[168] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__168_ : 1'b0;
  assign data_o_flat[167] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__167_ : 1'b0;
  assign data_o_flat[166] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__166_ : 1'b0;
  assign data_o_flat[165] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__165_ : 1'b0;
  assign data_o_flat[164] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__164_ : 1'b0;
  assign data_o_flat[163] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__163_ : 1'b0;
  assign data_o_flat[162] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__162_ : 1'b0;
  assign data_o_flat[161] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__161_ : 1'b0;
  assign data_o_flat[160] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__160_ : 1'b0;
  assign data_o_flat[159] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__159_ : 1'b0;
  assign data_o_flat[158] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__158_ : 1'b0;
  assign data_o_flat[157] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__157_ : 1'b0;
  assign data_o_flat[156] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__156_ : 1'b0;
  assign data_o_flat[155] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__155_ : 1'b0;
  assign data_o_flat[154] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__154_ : 1'b0;
  assign data_o_flat[153] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__153_ : 1'b0;
  assign data_o_flat[152] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__152_ : 1'b0;
  assign data_o_flat[151] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__151_ : 1'b0;
  assign data_o_flat[150] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__150_ : 1'b0;
  assign data_o_flat[149] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__149_ : 1'b0;
  assign data_o_flat[148] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__148_ : 1'b0;
  assign data_o_flat[147] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__147_ : 1'b0;
  assign data_o_flat[146] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__146_ : 1'b0;
  assign data_o_flat[145] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__145_ : 1'b0;
  assign data_o_flat[144] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__144_ : 1'b0;
  assign data_o_flat[143] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__143_ : 1'b0;
  assign data_o_flat[142] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__142_ : 1'b0;
  assign data_o_flat[141] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__141_ : 1'b0;
  assign data_o_flat[140] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__140_ : 1'b0;
  assign data_o_flat[139] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__139_ : 1'b0;
  assign data_o_flat[138] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__138_ : 1'b0;
  assign data_o_flat[137] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__137_ : 1'b0;
  assign data_o_flat[136] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__136_ : 1'b0;
  assign data_o_flat[135] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__135_ : 1'b0;
  assign data_o_flat[134] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__134_ : 1'b0;
  assign data_o_flat[133] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__133_ : 1'b0;
  assign data_o_flat[132] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__132_ : 1'b0;
  assign data_o_flat[131] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__131_ : 1'b0;
  assign data_o_flat[130] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__130_ : 1'b0;
  assign data_o_flat[129] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__129_ : 1'b0;
  assign data_o_flat[128] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__128_ : 1'b0;
  assign data_o_flat[127] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__127_ : 1'b0;
  assign data_o_flat[126] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__126_ : 1'b0;
  assign data_o_flat[125] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__125_ : 1'b0;
  assign data_o_flat[124] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__124_ : 1'b0;
  assign data_o_flat[123] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__123_ : 1'b0;
  assign data_o_flat[122] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__122_ : 1'b0;
  assign data_o_flat[121] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__121_ : 1'b0;
  assign data_o_flat[120] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__120_ : 1'b0;
  assign data_o_flat[119] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__119_ : 1'b0;
  assign data_o_flat[118] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__118_ : 1'b0;
  assign data_o_flat[117] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__117_ : 1'b0;
  assign data_o_flat[116] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__116_ : 1'b0;
  assign data_o_flat[115] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__115_ : 1'b0;
  assign data_o_flat[114] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__114_ : 1'b0;
  assign data_o_flat[113] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__113_ : 1'b0;
  assign data_o_flat[112] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__112_ : 1'b0;
  assign data_o_flat[111] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__111_ : 1'b0;
  assign data_o_flat[110] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__110_ : 1'b0;
  assign data_o_flat[109] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__109_ : 1'b0;
  assign data_o_flat[108] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__108_ : 1'b0;
  assign data_o_flat[107] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__107_ : 1'b0;
  assign data_o_flat[106] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__106_ : 1'b0;
  assign data_o_flat[105] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__105_ : 1'b0;
  assign data_o_flat[104] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__104_ : 1'b0;
  assign data_o_flat[103] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__103_ : 1'b0;
  assign data_o_flat[102] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__102_ : 1'b0;
  assign data_o_flat[101] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__101_ : 1'b0;
  assign data_o_flat[100] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__100_ : 1'b0;
  assign data_o_flat[99] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__99_ : 1'b0;
  assign data_o_flat[98] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__98_ : 1'b0;
  assign data_o_flat[97] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__97_ : 1'b0;
  assign data_o_flat[96] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__96_ : 1'b0;
  assign data_o_flat[95] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__95_ : 1'b0;
  assign data_o_flat[94] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__94_ : 1'b0;
  assign data_o_flat[93] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__93_ : 1'b0;
  assign data_o_flat[92] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__92_ : 1'b0;
  assign data_o_flat[91] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__91_ : 1'b0;
  assign data_o_flat[90] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__90_ : 1'b0;
  assign data_o_flat[89] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__89_ : 1'b0;
  assign data_o_flat[88] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__88_ : 1'b0;
  assign data_o_flat[87] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__87_ : 1'b0;
  assign data_o_flat[86] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__86_ : 1'b0;
  assign data_o_flat[85] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__85_ : 1'b0;
  assign data_o_flat[84] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__84_ : 1'b0;
  assign data_o_flat[83] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__83_ : 1'b0;
  assign data_o_flat[82] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__82_ : 1'b0;
  assign data_o_flat[81] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__81_ : 1'b0;
  assign data_o_flat[80] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__80_ : 1'b0;
  assign data_o_flat[79] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__79_ : 1'b0;
  assign data_o_flat[78] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__78_ : 1'b0;
  assign data_o_flat[77] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__77_ : 1'b0;
  assign data_o_flat[76] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__76_ : 1'b0;
  assign data_o_flat[75] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__75_ : 1'b0;
  assign data_o_flat[74] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__74_ : 1'b0;
  assign data_o_flat[73] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__73_ : 1'b0;
  assign data_o_flat[72] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__72_ : 1'b0;
  assign data_o_flat[71] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__71_ : 1'b0;
  assign data_o_flat[70] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__70_ : 1'b0;
  assign data_o_flat[69] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__69_ : 1'b0;
  assign data_o_flat[68] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__68_ : 1'b0;
  assign data_o_flat[67] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__67_ : 1'b0;
  assign data_o_flat[66] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__66_ : 1'b0;
  assign data_o_flat[65] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__65_ : 1'b0;
  assign data_o_flat[64] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__64_ : 1'b0;
  assign data_o_flat[63] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__63_ : 1'b0;
  assign data_o_flat[62] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__62_ : 1'b0;
  assign data_o_flat[61] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__61_ : 1'b0;
  assign data_o_flat[60] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__60_ : 1'b0;
  assign data_o_flat[59] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__59_ : 1'b0;
  assign data_o_flat[58] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__58_ : 1'b0;
  assign data_o_flat[57] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__57_ : 1'b0;
  assign data_o_flat[56] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__56_ : 1'b0;
  assign data_o_flat[55] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__55_ : 1'b0;
  assign data_o_flat[54] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__54_ : 1'b0;
  assign data_o_flat[53] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__53_ : 1'b0;
  assign data_o_flat[52] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__52_ : 1'b0;
  assign data_o_flat[51] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__51_ : 1'b0;
  assign data_o_flat[50] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__50_ : 1'b0;
  assign data_o_flat[49] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__49_ : 1'b0;
  assign data_o_flat[48] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__48_ : 1'b0;
  assign data_o_flat[47] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__47_ : 1'b0;
  assign data_o_flat[46] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__46_ : 1'b0;
  assign data_o_flat[45] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__45_ : 1'b0;
  assign data_o_flat[44] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__44_ : 1'b0;
  assign data_o_flat[43] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__43_ : 1'b0;
  assign data_o_flat[42] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__42_ : 1'b0;
  assign data_o_flat[41] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__41_ : 1'b0;
  assign data_o_flat[40] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__40_ : 1'b0;
  assign data_o_flat[39] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__39_ : 1'b0;
  assign data_o_flat[38] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__38_ : 1'b0;
  assign data_o_flat[37] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__37_ : 1'b0;
  assign data_o_flat[36] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__36_ : 1'b0;
  assign data_o_flat[35] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__35_ : 1'b0;
  assign data_o_flat[34] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__34_ : 1'b0;
  assign data_o_flat[33] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__33_ : 1'b0;
  assign data_o_flat[32] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__32_ : 1'b0;
  assign data_o_flat[31] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__31_ : 1'b0;
  assign data_o_flat[30] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__30_ : 1'b0;
  assign data_o_flat[29] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__29_ : 1'b0;
  assign data_o_flat[28] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__28_ : 1'b0;
  assign data_o_flat[27] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__27_ : 1'b0;
  assign data_o_flat[26] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__26_ : 1'b0;
  assign data_o_flat[25] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__25_ : 1'b0;
  assign data_o_flat[24] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__24_ : 1'b0;
  assign data_o_flat[23] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__23_ : 1'b0;
  assign data_o_flat[22] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__22_ : 1'b0;
  assign data_o_flat[21] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__21_ : 1'b0;
  assign data_o_flat[20] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__20_ : 1'b0;
  assign data_o_flat[19] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__19_ : 1'b0;
  assign data_o_flat[18] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__18_ : 1'b0;
  assign data_o_flat[17] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__17_ : 1'b0;
  assign data_o_flat[16] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__16_ : 1'b0;
  assign data_o_flat[15] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__15_ : 1'b0;
  assign data_o_flat[14] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__14_ : 1'b0;
  assign data_o_flat[13] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__13_ : 1'b0;
  assign data_o_flat[12] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__12_ : 1'b0;
  assign data_o_flat[11] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__11_ : 1'b0;
  assign data_o_flat[10] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__10_ : 1'b0;
  assign data_o_flat[9] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__9_ : 1'b0;
  assign data_o_flat[8] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__8_ : 1'b0;
  assign data_o_flat[7] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__7_ : 1'b0;
  assign data_o_flat[6] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__6_ : 1'b0;
  assign data_o_flat[5] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__5_ : 1'b0;
  assign data_o_flat[4] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__4_ : 1'b0;
  assign data_o_flat[3] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__3_ : 1'b0;
  assign data_o_flat[2] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__2_ : 1'b0;
  assign data_o_flat[1] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__1_ : 1'b0;
  assign data_o_flat[0] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__0_ : 1'b0;
  assign n_2_net__9_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__9_ : 1'b0;
  assign N105 = N155;
  assign N106 = N157;
  assign N107 = N159;
  assign N108 = N160;
  assign N109 = N161;
  assign N110 = N162;
  assign N111 = N163;
  assign N112 = N164;
  assign N113 = N156;
  assign N114 = N158;
  assign n_2_net__8_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__8_ : 1'b0;
  assign n_2_net__7_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__7_ : 1'b0;
  assign n_2_net__6_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__6_ : 1'b0;
  assign n_2_net__5_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__5_ : 1'b0;
  assign n_2_net__4_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__4_ : 1'b0;
  assign n_2_net__3_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__3_ : 1'b0;
  assign n_2_net__2_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__2_ : 1'b0;
  assign n_2_net__1_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__1_ : 1'b0;
  assign n_2_net__0_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__0_ : 1'b0;
  assign n_3_net__9_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__9_ : 1'b0;
  assign n_3_net__8_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__8_ : 1'b0;
  assign n_3_net__7_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__7_ : 1'b0;
  assign n_3_net__6_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__6_ : 1'b0;
  assign n_3_net__5_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__5_ : 1'b0;
  assign n_3_net__4_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__4_ : 1'b0;
  assign n_3_net__3_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__3_ : 1'b0;
  assign n_3_net__2_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__2_ : 1'b0;
  assign n_3_net__1_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__1_ : 1'b0;
  assign n_3_net__0_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__0_ : 1'b0;
  assign n_4_net__639_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__639_ : 1'b0;
  assign N115 = N165;
  assign N116 = N167;
  assign N117 = N169;
  assign N118 = N170;
  assign N119 = N171;
  assign N120 = N172;
  assign N121 = N173;
  assign N122 = N174;
  assign N123 = N166;
  assign N124 = N168;
  assign n_4_net__638_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__638_ : 1'b0;
  assign n_4_net__637_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__637_ : 1'b0;
  assign n_4_net__636_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__636_ : 1'b0;
  assign n_4_net__635_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__635_ : 1'b0;
  assign n_4_net__634_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__634_ : 1'b0;
  assign n_4_net__633_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__633_ : 1'b0;
  assign n_4_net__632_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__632_ : 1'b0;
  assign n_4_net__631_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__631_ : 1'b0;
  assign n_4_net__630_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__630_ : 1'b0;
  assign n_4_net__629_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__629_ : 1'b0;
  assign n_4_net__628_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__628_ : 1'b0;
  assign n_4_net__627_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__627_ : 1'b0;
  assign n_4_net__626_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__626_ : 1'b0;
  assign n_4_net__625_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__625_ : 1'b0;
  assign n_4_net__624_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__624_ : 1'b0;
  assign n_4_net__623_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__623_ : 1'b0;
  assign n_4_net__622_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__622_ : 1'b0;
  assign n_4_net__621_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__621_ : 1'b0;
  assign n_4_net__620_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__620_ : 1'b0;
  assign n_4_net__619_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__619_ : 1'b0;
  assign n_4_net__618_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__618_ : 1'b0;
  assign n_4_net__617_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__617_ : 1'b0;
  assign n_4_net__616_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__616_ : 1'b0;
  assign n_4_net__615_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__615_ : 1'b0;
  assign n_4_net__614_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__614_ : 1'b0;
  assign n_4_net__613_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__613_ : 1'b0;
  assign n_4_net__612_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__612_ : 1'b0;
  assign n_4_net__611_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__611_ : 1'b0;
  assign n_4_net__610_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__610_ : 1'b0;
  assign n_4_net__609_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__609_ : 1'b0;
  assign n_4_net__608_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__608_ : 1'b0;
  assign n_4_net__607_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__607_ : 1'b0;
  assign n_4_net__606_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__606_ : 1'b0;
  assign n_4_net__605_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__605_ : 1'b0;
  assign n_4_net__604_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__604_ : 1'b0;
  assign n_4_net__603_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__603_ : 1'b0;
  assign n_4_net__602_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__602_ : 1'b0;
  assign n_4_net__601_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__601_ : 1'b0;
  assign n_4_net__600_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__600_ : 1'b0;
  assign n_4_net__599_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__599_ : 1'b0;
  assign n_4_net__598_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__598_ : 1'b0;
  assign n_4_net__597_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__597_ : 1'b0;
  assign n_4_net__596_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__596_ : 1'b0;
  assign n_4_net__595_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__595_ : 1'b0;
  assign n_4_net__594_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__594_ : 1'b0;
  assign n_4_net__593_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__593_ : 1'b0;
  assign n_4_net__592_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__592_ : 1'b0;
  assign n_4_net__591_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__591_ : 1'b0;
  assign n_4_net__590_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__590_ : 1'b0;
  assign n_4_net__589_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__589_ : 1'b0;
  assign n_4_net__588_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__588_ : 1'b0;
  assign n_4_net__587_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__587_ : 1'b0;
  assign n_4_net__586_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__586_ : 1'b0;
  assign n_4_net__585_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__585_ : 1'b0;
  assign n_4_net__584_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__584_ : 1'b0;
  assign n_4_net__583_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__583_ : 1'b0;
  assign n_4_net__582_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__582_ : 1'b0;
  assign n_4_net__581_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__581_ : 1'b0;
  assign n_4_net__580_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__580_ : 1'b0;
  assign n_4_net__579_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__579_ : 1'b0;
  assign n_4_net__578_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__578_ : 1'b0;
  assign n_4_net__577_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__577_ : 1'b0;
  assign n_4_net__576_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__576_ : 1'b0;
  assign n_4_net__575_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__575_ : 1'b0;
  assign n_4_net__574_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__574_ : 1'b0;
  assign n_4_net__573_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__573_ : 1'b0;
  assign n_4_net__572_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__572_ : 1'b0;
  assign n_4_net__571_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__571_ : 1'b0;
  assign n_4_net__570_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__570_ : 1'b0;
  assign n_4_net__569_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__569_ : 1'b0;
  assign n_4_net__568_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__568_ : 1'b0;
  assign n_4_net__567_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__567_ : 1'b0;
  assign n_4_net__566_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__566_ : 1'b0;
  assign n_4_net__565_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__565_ : 1'b0;
  assign n_4_net__564_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__564_ : 1'b0;
  assign n_4_net__563_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__563_ : 1'b0;
  assign n_4_net__562_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__562_ : 1'b0;
  assign n_4_net__561_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__561_ : 1'b0;
  assign n_4_net__560_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__560_ : 1'b0;
  assign n_4_net__559_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__559_ : 1'b0;
  assign n_4_net__558_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__558_ : 1'b0;
  assign n_4_net__557_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__557_ : 1'b0;
  assign n_4_net__556_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__556_ : 1'b0;
  assign n_4_net__555_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__555_ : 1'b0;
  assign n_4_net__554_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__554_ : 1'b0;
  assign n_4_net__553_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__553_ : 1'b0;
  assign n_4_net__552_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__552_ : 1'b0;
  assign n_4_net__551_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__551_ : 1'b0;
  assign n_4_net__550_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__550_ : 1'b0;
  assign n_4_net__549_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__549_ : 1'b0;
  assign n_4_net__548_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__548_ : 1'b0;
  assign n_4_net__547_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__547_ : 1'b0;
  assign n_4_net__546_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__546_ : 1'b0;
  assign n_4_net__545_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__545_ : 1'b0;
  assign n_4_net__544_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__544_ : 1'b0;
  assign n_4_net__543_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__543_ : 1'b0;
  assign n_4_net__542_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__542_ : 1'b0;
  assign n_4_net__541_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__541_ : 1'b0;
  assign n_4_net__540_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__540_ : 1'b0;
  assign n_4_net__539_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__539_ : 1'b0;
  assign n_4_net__538_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__538_ : 1'b0;
  assign n_4_net__537_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__537_ : 1'b0;
  assign n_4_net__536_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__536_ : 1'b0;
  assign n_4_net__535_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__535_ : 1'b0;
  assign n_4_net__534_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__534_ : 1'b0;
  assign n_4_net__533_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__533_ : 1'b0;
  assign n_4_net__532_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__532_ : 1'b0;
  assign n_4_net__531_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__531_ : 1'b0;
  assign n_4_net__530_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__530_ : 1'b0;
  assign n_4_net__529_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__529_ : 1'b0;
  assign n_4_net__528_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__528_ : 1'b0;
  assign n_4_net__527_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__527_ : 1'b0;
  assign n_4_net__526_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__526_ : 1'b0;
  assign n_4_net__525_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__525_ : 1'b0;
  assign n_4_net__524_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__524_ : 1'b0;
  assign n_4_net__523_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__523_ : 1'b0;
  assign n_4_net__522_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__522_ : 1'b0;
  assign n_4_net__521_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__521_ : 1'b0;
  assign n_4_net__520_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__520_ : 1'b0;
  assign n_4_net__519_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__519_ : 1'b0;
  assign n_4_net__518_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__518_ : 1'b0;
  assign n_4_net__517_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__517_ : 1'b0;
  assign n_4_net__516_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__516_ : 1'b0;
  assign n_4_net__515_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__515_ : 1'b0;
  assign n_4_net__514_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__514_ : 1'b0;
  assign n_4_net__513_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__513_ : 1'b0;
  assign n_4_net__512_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__512_ : 1'b0;
  assign n_4_net__511_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__511_ : 1'b0;
  assign n_4_net__510_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__510_ : 1'b0;
  assign n_4_net__509_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__509_ : 1'b0;
  assign n_4_net__508_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__508_ : 1'b0;
  assign n_4_net__507_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__507_ : 1'b0;
  assign n_4_net__506_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__506_ : 1'b0;
  assign n_4_net__505_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__505_ : 1'b0;
  assign n_4_net__504_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__504_ : 1'b0;
  assign n_4_net__503_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__503_ : 1'b0;
  assign n_4_net__502_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__502_ : 1'b0;
  assign n_4_net__501_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__501_ : 1'b0;
  assign n_4_net__500_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__500_ : 1'b0;
  assign n_4_net__499_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__499_ : 1'b0;
  assign n_4_net__498_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__498_ : 1'b0;
  assign n_4_net__497_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__497_ : 1'b0;
  assign n_4_net__496_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__496_ : 1'b0;
  assign n_4_net__495_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__495_ : 1'b0;
  assign n_4_net__494_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__494_ : 1'b0;
  assign n_4_net__493_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__493_ : 1'b0;
  assign n_4_net__492_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__492_ : 1'b0;
  assign n_4_net__491_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__491_ : 1'b0;
  assign n_4_net__490_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__490_ : 1'b0;
  assign n_4_net__489_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__489_ : 1'b0;
  assign n_4_net__488_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__488_ : 1'b0;
  assign n_4_net__487_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__487_ : 1'b0;
  assign n_4_net__486_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__486_ : 1'b0;
  assign n_4_net__485_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__485_ : 1'b0;
  assign n_4_net__484_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__484_ : 1'b0;
  assign n_4_net__483_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__483_ : 1'b0;
  assign n_4_net__482_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__482_ : 1'b0;
  assign n_4_net__481_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__481_ : 1'b0;
  assign n_4_net__480_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__480_ : 1'b0;
  assign n_4_net__479_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__479_ : 1'b0;
  assign n_4_net__478_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__478_ : 1'b0;
  assign n_4_net__477_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__477_ : 1'b0;
  assign n_4_net__476_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__476_ : 1'b0;
  assign n_4_net__475_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__475_ : 1'b0;
  assign n_4_net__474_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__474_ : 1'b0;
  assign n_4_net__473_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__473_ : 1'b0;
  assign n_4_net__472_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__472_ : 1'b0;
  assign n_4_net__471_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__471_ : 1'b0;
  assign n_4_net__470_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__470_ : 1'b0;
  assign n_4_net__469_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__469_ : 1'b0;
  assign n_4_net__468_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__468_ : 1'b0;
  assign n_4_net__467_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__467_ : 1'b0;
  assign n_4_net__466_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__466_ : 1'b0;
  assign n_4_net__465_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__465_ : 1'b0;
  assign n_4_net__464_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__464_ : 1'b0;
  assign n_4_net__463_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__463_ : 1'b0;
  assign n_4_net__462_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__462_ : 1'b0;
  assign n_4_net__461_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__461_ : 1'b0;
  assign n_4_net__460_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__460_ : 1'b0;
  assign n_4_net__459_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__459_ : 1'b0;
  assign n_4_net__458_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__458_ : 1'b0;
  assign n_4_net__457_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__457_ : 1'b0;
  assign n_4_net__456_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__456_ : 1'b0;
  assign n_4_net__455_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__455_ : 1'b0;
  assign n_4_net__454_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__454_ : 1'b0;
  assign n_4_net__453_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__453_ : 1'b0;
  assign n_4_net__452_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__452_ : 1'b0;
  assign n_4_net__451_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__451_ : 1'b0;
  assign n_4_net__450_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__450_ : 1'b0;
  assign n_4_net__449_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__449_ : 1'b0;
  assign n_4_net__448_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__448_ : 1'b0;
  assign n_4_net__447_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__447_ : 1'b0;
  assign n_4_net__446_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__446_ : 1'b0;
  assign n_4_net__445_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__445_ : 1'b0;
  assign n_4_net__444_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__444_ : 1'b0;
  assign n_4_net__443_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__443_ : 1'b0;
  assign n_4_net__442_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__442_ : 1'b0;
  assign n_4_net__441_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__441_ : 1'b0;
  assign n_4_net__440_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__440_ : 1'b0;
  assign n_4_net__439_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__439_ : 1'b0;
  assign n_4_net__438_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__438_ : 1'b0;
  assign n_4_net__437_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__437_ : 1'b0;
  assign n_4_net__436_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__436_ : 1'b0;
  assign n_4_net__435_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__435_ : 1'b0;
  assign n_4_net__434_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__434_ : 1'b0;
  assign n_4_net__433_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__433_ : 1'b0;
  assign n_4_net__432_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__432_ : 1'b0;
  assign n_4_net__431_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__431_ : 1'b0;
  assign n_4_net__430_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__430_ : 1'b0;
  assign n_4_net__429_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__429_ : 1'b0;
  assign n_4_net__428_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__428_ : 1'b0;
  assign n_4_net__427_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__427_ : 1'b0;
  assign n_4_net__426_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__426_ : 1'b0;
  assign n_4_net__425_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__425_ : 1'b0;
  assign n_4_net__424_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__424_ : 1'b0;
  assign n_4_net__423_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__423_ : 1'b0;
  assign n_4_net__422_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__422_ : 1'b0;
  assign n_4_net__421_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__421_ : 1'b0;
  assign n_4_net__420_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__420_ : 1'b0;
  assign n_4_net__419_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__419_ : 1'b0;
  assign n_4_net__418_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__418_ : 1'b0;
  assign n_4_net__417_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__417_ : 1'b0;
  assign n_4_net__416_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__416_ : 1'b0;
  assign n_4_net__415_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__415_ : 1'b0;
  assign n_4_net__414_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__414_ : 1'b0;
  assign n_4_net__413_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__413_ : 1'b0;
  assign n_4_net__412_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__412_ : 1'b0;
  assign n_4_net__411_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__411_ : 1'b0;
  assign n_4_net__410_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__410_ : 1'b0;
  assign n_4_net__409_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__409_ : 1'b0;
  assign n_4_net__408_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__408_ : 1'b0;
  assign n_4_net__407_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__407_ : 1'b0;
  assign n_4_net__406_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__406_ : 1'b0;
  assign n_4_net__405_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__405_ : 1'b0;
  assign n_4_net__404_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__404_ : 1'b0;
  assign n_4_net__403_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__403_ : 1'b0;
  assign n_4_net__402_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__402_ : 1'b0;
  assign n_4_net__401_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__401_ : 1'b0;
  assign n_4_net__400_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__400_ : 1'b0;
  assign n_4_net__399_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__399_ : 1'b0;
  assign n_4_net__398_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__398_ : 1'b0;
  assign n_4_net__397_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__397_ : 1'b0;
  assign n_4_net__396_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__396_ : 1'b0;
  assign n_4_net__395_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__395_ : 1'b0;
  assign n_4_net__394_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__394_ : 1'b0;
  assign n_4_net__393_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__393_ : 1'b0;
  assign n_4_net__392_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__392_ : 1'b0;
  assign n_4_net__391_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__391_ : 1'b0;
  assign n_4_net__390_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__390_ : 1'b0;
  assign n_4_net__389_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__389_ : 1'b0;
  assign n_4_net__388_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__388_ : 1'b0;
  assign n_4_net__387_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__387_ : 1'b0;
  assign n_4_net__386_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__386_ : 1'b0;
  assign n_4_net__385_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__385_ : 1'b0;
  assign n_4_net__384_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__384_ : 1'b0;
  assign n_4_net__383_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__383_ : 1'b0;
  assign n_4_net__382_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__382_ : 1'b0;
  assign n_4_net__381_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__381_ : 1'b0;
  assign n_4_net__380_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__380_ : 1'b0;
  assign n_4_net__379_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__379_ : 1'b0;
  assign n_4_net__378_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__378_ : 1'b0;
  assign n_4_net__377_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__377_ : 1'b0;
  assign n_4_net__376_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__376_ : 1'b0;
  assign n_4_net__375_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__375_ : 1'b0;
  assign n_4_net__374_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__374_ : 1'b0;
  assign n_4_net__373_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__373_ : 1'b0;
  assign n_4_net__372_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__372_ : 1'b0;
  assign n_4_net__371_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__371_ : 1'b0;
  assign n_4_net__370_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__370_ : 1'b0;
  assign n_4_net__369_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__369_ : 1'b0;
  assign n_4_net__368_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__368_ : 1'b0;
  assign n_4_net__367_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__367_ : 1'b0;
  assign n_4_net__366_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__366_ : 1'b0;
  assign n_4_net__365_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__365_ : 1'b0;
  assign n_4_net__364_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__364_ : 1'b0;
  assign n_4_net__363_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__363_ : 1'b0;
  assign n_4_net__362_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__362_ : 1'b0;
  assign n_4_net__361_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__361_ : 1'b0;
  assign n_4_net__360_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__360_ : 1'b0;
  assign n_4_net__359_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__359_ : 1'b0;
  assign n_4_net__358_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__358_ : 1'b0;
  assign n_4_net__357_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__357_ : 1'b0;
  assign n_4_net__356_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__356_ : 1'b0;
  assign n_4_net__355_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__355_ : 1'b0;
  assign n_4_net__354_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__354_ : 1'b0;
  assign n_4_net__353_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__353_ : 1'b0;
  assign n_4_net__352_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__352_ : 1'b0;
  assign n_4_net__351_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__351_ : 1'b0;
  assign n_4_net__350_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__350_ : 1'b0;
  assign n_4_net__349_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__349_ : 1'b0;
  assign n_4_net__348_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__348_ : 1'b0;
  assign n_4_net__347_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__347_ : 1'b0;
  assign n_4_net__346_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__346_ : 1'b0;
  assign n_4_net__345_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__345_ : 1'b0;
  assign n_4_net__344_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__344_ : 1'b0;
  assign n_4_net__343_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__343_ : 1'b0;
  assign n_4_net__342_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__342_ : 1'b0;
  assign n_4_net__341_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__341_ : 1'b0;
  assign n_4_net__340_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__340_ : 1'b0;
  assign n_4_net__339_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__339_ : 1'b0;
  assign n_4_net__338_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__338_ : 1'b0;
  assign n_4_net__337_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__337_ : 1'b0;
  assign n_4_net__336_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__336_ : 1'b0;
  assign n_4_net__335_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__335_ : 1'b0;
  assign n_4_net__334_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__334_ : 1'b0;
  assign n_4_net__333_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__333_ : 1'b0;
  assign n_4_net__332_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__332_ : 1'b0;
  assign n_4_net__331_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__331_ : 1'b0;
  assign n_4_net__330_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__330_ : 1'b0;
  assign n_4_net__329_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__329_ : 1'b0;
  assign n_4_net__328_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__328_ : 1'b0;
  assign n_4_net__327_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__327_ : 1'b0;
  assign n_4_net__326_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__326_ : 1'b0;
  assign n_4_net__325_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__325_ : 1'b0;
  assign n_4_net__324_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__324_ : 1'b0;
  assign n_4_net__323_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__323_ : 1'b0;
  assign n_4_net__322_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__322_ : 1'b0;
  assign n_4_net__321_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__321_ : 1'b0;
  assign n_4_net__320_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__320_ : 1'b0;
  assign n_4_net__319_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__319_ : 1'b0;
  assign n_4_net__318_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__318_ : 1'b0;
  assign n_4_net__317_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__317_ : 1'b0;
  assign n_4_net__316_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__316_ : 1'b0;
  assign n_4_net__315_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__315_ : 1'b0;
  assign n_4_net__314_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__314_ : 1'b0;
  assign n_4_net__313_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__313_ : 1'b0;
  assign n_4_net__312_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__312_ : 1'b0;
  assign n_4_net__311_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__311_ : 1'b0;
  assign n_4_net__310_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__310_ : 1'b0;
  assign n_4_net__309_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__309_ : 1'b0;
  assign n_4_net__308_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__308_ : 1'b0;
  assign n_4_net__307_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__307_ : 1'b0;
  assign n_4_net__306_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__306_ : 1'b0;
  assign n_4_net__305_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__305_ : 1'b0;
  assign n_4_net__304_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__304_ : 1'b0;
  assign n_4_net__303_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__303_ : 1'b0;
  assign n_4_net__302_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__302_ : 1'b0;
  assign n_4_net__301_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__301_ : 1'b0;
  assign n_4_net__300_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__300_ : 1'b0;
  assign n_4_net__299_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__299_ : 1'b0;
  assign n_4_net__298_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__298_ : 1'b0;
  assign n_4_net__297_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__297_ : 1'b0;
  assign n_4_net__296_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__296_ : 1'b0;
  assign n_4_net__295_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__295_ : 1'b0;
  assign n_4_net__294_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__294_ : 1'b0;
  assign n_4_net__293_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__293_ : 1'b0;
  assign n_4_net__292_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__292_ : 1'b0;
  assign n_4_net__291_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__291_ : 1'b0;
  assign n_4_net__290_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__290_ : 1'b0;
  assign n_4_net__289_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__289_ : 1'b0;
  assign n_4_net__288_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__288_ : 1'b0;
  assign n_4_net__287_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__287_ : 1'b0;
  assign n_4_net__286_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__286_ : 1'b0;
  assign n_4_net__285_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__285_ : 1'b0;
  assign n_4_net__284_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__284_ : 1'b0;
  assign n_4_net__283_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__283_ : 1'b0;
  assign n_4_net__282_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__282_ : 1'b0;
  assign n_4_net__281_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__281_ : 1'b0;
  assign n_4_net__280_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__280_ : 1'b0;
  assign n_4_net__279_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__279_ : 1'b0;
  assign n_4_net__278_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__278_ : 1'b0;
  assign n_4_net__277_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__277_ : 1'b0;
  assign n_4_net__276_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__276_ : 1'b0;
  assign n_4_net__275_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__275_ : 1'b0;
  assign n_4_net__274_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__274_ : 1'b0;
  assign n_4_net__273_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__273_ : 1'b0;
  assign n_4_net__272_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__272_ : 1'b0;
  assign n_4_net__271_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__271_ : 1'b0;
  assign n_4_net__270_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__270_ : 1'b0;
  assign n_4_net__269_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__269_ : 1'b0;
  assign n_4_net__268_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__268_ : 1'b0;
  assign n_4_net__267_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__267_ : 1'b0;
  assign n_4_net__266_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__266_ : 1'b0;
  assign n_4_net__265_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__265_ : 1'b0;
  assign n_4_net__264_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__264_ : 1'b0;
  assign n_4_net__263_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__263_ : 1'b0;
  assign n_4_net__262_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__262_ : 1'b0;
  assign n_4_net__261_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__261_ : 1'b0;
  assign n_4_net__260_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__260_ : 1'b0;
  assign n_4_net__259_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__259_ : 1'b0;
  assign n_4_net__258_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__258_ : 1'b0;
  assign n_4_net__257_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__257_ : 1'b0;
  assign n_4_net__256_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__256_ : 1'b0;
  assign n_4_net__255_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__255_ : 1'b0;
  assign n_4_net__254_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__254_ : 1'b0;
  assign n_4_net__253_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__253_ : 1'b0;
  assign n_4_net__252_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__252_ : 1'b0;
  assign n_4_net__251_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__251_ : 1'b0;
  assign n_4_net__250_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__250_ : 1'b0;
  assign n_4_net__249_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__249_ : 1'b0;
  assign n_4_net__248_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__248_ : 1'b0;
  assign n_4_net__247_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__247_ : 1'b0;
  assign n_4_net__246_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__246_ : 1'b0;
  assign n_4_net__245_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__245_ : 1'b0;
  assign n_4_net__244_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__244_ : 1'b0;
  assign n_4_net__243_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__243_ : 1'b0;
  assign n_4_net__242_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__242_ : 1'b0;
  assign n_4_net__241_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__241_ : 1'b0;
  assign n_4_net__240_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__240_ : 1'b0;
  assign n_4_net__239_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__239_ : 1'b0;
  assign n_4_net__238_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__238_ : 1'b0;
  assign n_4_net__237_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__237_ : 1'b0;
  assign n_4_net__236_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__236_ : 1'b0;
  assign n_4_net__235_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__235_ : 1'b0;
  assign n_4_net__234_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__234_ : 1'b0;
  assign n_4_net__233_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__233_ : 1'b0;
  assign n_4_net__232_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__232_ : 1'b0;
  assign n_4_net__231_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__231_ : 1'b0;
  assign n_4_net__230_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__230_ : 1'b0;
  assign n_4_net__229_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__229_ : 1'b0;
  assign n_4_net__228_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__228_ : 1'b0;
  assign n_4_net__227_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__227_ : 1'b0;
  assign n_4_net__226_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__226_ : 1'b0;
  assign n_4_net__225_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__225_ : 1'b0;
  assign n_4_net__224_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__224_ : 1'b0;
  assign n_4_net__223_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__223_ : 1'b0;
  assign n_4_net__222_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__222_ : 1'b0;
  assign n_4_net__221_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__221_ : 1'b0;
  assign n_4_net__220_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__220_ : 1'b0;
  assign n_4_net__219_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__219_ : 1'b0;
  assign n_4_net__218_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__218_ : 1'b0;
  assign n_4_net__217_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__217_ : 1'b0;
  assign n_4_net__216_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__216_ : 1'b0;
  assign n_4_net__215_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__215_ : 1'b0;
  assign n_4_net__214_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__214_ : 1'b0;
  assign n_4_net__213_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__213_ : 1'b0;
  assign n_4_net__212_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__212_ : 1'b0;
  assign n_4_net__211_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__211_ : 1'b0;
  assign n_4_net__210_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__210_ : 1'b0;
  assign n_4_net__209_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__209_ : 1'b0;
  assign n_4_net__208_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__208_ : 1'b0;
  assign n_4_net__207_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__207_ : 1'b0;
  assign n_4_net__206_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__206_ : 1'b0;
  assign n_4_net__205_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__205_ : 1'b0;
  assign n_4_net__204_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__204_ : 1'b0;
  assign n_4_net__203_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__203_ : 1'b0;
  assign n_4_net__202_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__202_ : 1'b0;
  assign n_4_net__201_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__201_ : 1'b0;
  assign n_4_net__200_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__200_ : 1'b0;
  assign n_4_net__199_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__199_ : 1'b0;
  assign n_4_net__198_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__198_ : 1'b0;
  assign n_4_net__197_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__197_ : 1'b0;
  assign n_4_net__196_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__196_ : 1'b0;
  assign n_4_net__195_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__195_ : 1'b0;
  assign n_4_net__194_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__194_ : 1'b0;
  assign n_4_net__193_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__193_ : 1'b0;
  assign n_4_net__192_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__192_ : 1'b0;
  assign n_4_net__191_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__191_ : 1'b0;
  assign n_4_net__190_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__190_ : 1'b0;
  assign n_4_net__189_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__189_ : 1'b0;
  assign n_4_net__188_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__188_ : 1'b0;
  assign n_4_net__187_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__187_ : 1'b0;
  assign n_4_net__186_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__186_ : 1'b0;
  assign n_4_net__185_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__185_ : 1'b0;
  assign n_4_net__184_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__184_ : 1'b0;
  assign n_4_net__183_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__183_ : 1'b0;
  assign n_4_net__182_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__182_ : 1'b0;
  assign n_4_net__181_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__181_ : 1'b0;
  assign n_4_net__180_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__180_ : 1'b0;
  assign n_4_net__179_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__179_ : 1'b0;
  assign n_4_net__178_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__178_ : 1'b0;
  assign n_4_net__177_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__177_ : 1'b0;
  assign n_4_net__176_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__176_ : 1'b0;
  assign n_4_net__175_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__175_ : 1'b0;
  assign n_4_net__174_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__174_ : 1'b0;
  assign n_4_net__173_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__173_ : 1'b0;
  assign n_4_net__172_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__172_ : 1'b0;
  assign n_4_net__171_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__171_ : 1'b0;
  assign n_4_net__170_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__170_ : 1'b0;
  assign n_4_net__169_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__169_ : 1'b0;
  assign n_4_net__168_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__168_ : 1'b0;
  assign n_4_net__167_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__167_ : 1'b0;
  assign n_4_net__166_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__166_ : 1'b0;
  assign n_4_net__165_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__165_ : 1'b0;
  assign n_4_net__164_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__164_ : 1'b0;
  assign n_4_net__163_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__163_ : 1'b0;
  assign n_4_net__162_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__162_ : 1'b0;
  assign n_4_net__161_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__161_ : 1'b0;
  assign n_4_net__160_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__160_ : 1'b0;
  assign n_4_net__159_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__159_ : 1'b0;
  assign n_4_net__158_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__158_ : 1'b0;
  assign n_4_net__157_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__157_ : 1'b0;
  assign n_4_net__156_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__156_ : 1'b0;
  assign n_4_net__155_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__155_ : 1'b0;
  assign n_4_net__154_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__154_ : 1'b0;
  assign n_4_net__153_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__153_ : 1'b0;
  assign n_4_net__152_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__152_ : 1'b0;
  assign n_4_net__151_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__151_ : 1'b0;
  assign n_4_net__150_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__150_ : 1'b0;
  assign n_4_net__149_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__149_ : 1'b0;
  assign n_4_net__148_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__148_ : 1'b0;
  assign n_4_net__147_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__147_ : 1'b0;
  assign n_4_net__146_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__146_ : 1'b0;
  assign n_4_net__145_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__145_ : 1'b0;
  assign n_4_net__144_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__144_ : 1'b0;
  assign n_4_net__143_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__143_ : 1'b0;
  assign n_4_net__142_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__142_ : 1'b0;
  assign n_4_net__141_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__141_ : 1'b0;
  assign n_4_net__140_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__140_ : 1'b0;
  assign n_4_net__139_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__139_ : 1'b0;
  assign n_4_net__138_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__138_ : 1'b0;
  assign n_4_net__137_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__137_ : 1'b0;
  assign n_4_net__136_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__136_ : 1'b0;
  assign n_4_net__135_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__135_ : 1'b0;
  assign n_4_net__134_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__134_ : 1'b0;
  assign n_4_net__133_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__133_ : 1'b0;
  assign n_4_net__132_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__132_ : 1'b0;
  assign n_4_net__131_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__131_ : 1'b0;
  assign n_4_net__130_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__130_ : 1'b0;
  assign n_4_net__129_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__129_ : 1'b0;
  assign n_4_net__128_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__128_ : 1'b0;
  assign n_4_net__127_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__127_ : 1'b0;
  assign n_4_net__126_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__126_ : 1'b0;
  assign n_4_net__125_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__125_ : 1'b0;
  assign n_4_net__124_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__124_ : 1'b0;
  assign n_4_net__123_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__123_ : 1'b0;
  assign n_4_net__122_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__122_ : 1'b0;
  assign n_4_net__121_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__121_ : 1'b0;
  assign n_4_net__120_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__120_ : 1'b0;
  assign n_4_net__119_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__119_ : 1'b0;
  assign n_4_net__118_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__118_ : 1'b0;
  assign n_4_net__117_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__117_ : 1'b0;
  assign n_4_net__116_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__116_ : 1'b0;
  assign n_4_net__115_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__115_ : 1'b0;
  assign n_4_net__114_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__114_ : 1'b0;
  assign n_4_net__113_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__113_ : 1'b0;
  assign n_4_net__112_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__112_ : 1'b0;
  assign n_4_net__111_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__111_ : 1'b0;
  assign n_4_net__110_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__110_ : 1'b0;
  assign n_4_net__109_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__109_ : 1'b0;
  assign n_4_net__108_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__108_ : 1'b0;
  assign n_4_net__107_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__107_ : 1'b0;
  assign n_4_net__106_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__106_ : 1'b0;
  assign n_4_net__105_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__105_ : 1'b0;
  assign n_4_net__104_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__104_ : 1'b0;
  assign n_4_net__103_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__103_ : 1'b0;
  assign n_4_net__102_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__102_ : 1'b0;
  assign n_4_net__101_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__101_ : 1'b0;
  assign n_4_net__100_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__100_ : 1'b0;
  assign n_4_net__99_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__99_ : 1'b0;
  assign n_4_net__98_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__98_ : 1'b0;
  assign n_4_net__97_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__97_ : 1'b0;
  assign n_4_net__96_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__96_ : 1'b0;
  assign n_4_net__95_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__95_ : 1'b0;
  assign n_4_net__94_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__94_ : 1'b0;
  assign n_4_net__93_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__93_ : 1'b0;
  assign n_4_net__92_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__92_ : 1'b0;
  assign n_4_net__91_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__91_ : 1'b0;
  assign n_4_net__90_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__90_ : 1'b0;
  assign n_4_net__89_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__89_ : 1'b0;
  assign n_4_net__88_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__88_ : 1'b0;
  assign n_4_net__87_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__87_ : 1'b0;
  assign n_4_net__86_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__86_ : 1'b0;
  assign n_4_net__85_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__85_ : 1'b0;
  assign n_4_net__84_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__84_ : 1'b0;
  assign n_4_net__83_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__83_ : 1'b0;
  assign n_4_net__82_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__82_ : 1'b0;
  assign n_4_net__81_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__81_ : 1'b0;
  assign n_4_net__80_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__80_ : 1'b0;
  assign n_4_net__79_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__79_ : 1'b0;
  assign n_4_net__78_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__78_ : 1'b0;
  assign n_4_net__77_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__77_ : 1'b0;
  assign n_4_net__76_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__76_ : 1'b0;
  assign n_4_net__75_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__75_ : 1'b0;
  assign n_4_net__74_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__74_ : 1'b0;
  assign n_4_net__73_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__73_ : 1'b0;
  assign n_4_net__72_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__72_ : 1'b0;
  assign n_4_net__71_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__71_ : 1'b0;
  assign n_4_net__70_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__70_ : 1'b0;
  assign n_4_net__69_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__69_ : 1'b0;
  assign n_4_net__68_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__68_ : 1'b0;
  assign n_4_net__67_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__67_ : 1'b0;
  assign n_4_net__66_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__66_ : 1'b0;
  assign n_4_net__65_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__65_ : 1'b0;
  assign n_4_net__64_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__64_ : 1'b0;
  assign n_4_net__63_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__63_ : 1'b0;
  assign n_4_net__62_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__62_ : 1'b0;
  assign n_4_net__61_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__61_ : 1'b0;
  assign n_4_net__60_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__60_ : 1'b0;
  assign n_4_net__59_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__59_ : 1'b0;
  assign n_4_net__58_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__58_ : 1'b0;
  assign n_4_net__57_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__57_ : 1'b0;
  assign n_4_net__56_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__56_ : 1'b0;
  assign n_4_net__55_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__55_ : 1'b0;
  assign n_4_net__54_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__54_ : 1'b0;
  assign n_4_net__53_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__53_ : 1'b0;
  assign n_4_net__52_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__52_ : 1'b0;
  assign n_4_net__51_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__51_ : 1'b0;
  assign n_4_net__50_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__50_ : 1'b0;
  assign n_4_net__49_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__49_ : 1'b0;
  assign n_4_net__48_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__48_ : 1'b0;
  assign n_4_net__47_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__47_ : 1'b0;
  assign n_4_net__46_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__46_ : 1'b0;
  assign n_4_net__45_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__45_ : 1'b0;
  assign n_4_net__44_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__44_ : 1'b0;
  assign n_4_net__43_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__43_ : 1'b0;
  assign n_4_net__42_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__42_ : 1'b0;
  assign n_4_net__41_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__41_ : 1'b0;
  assign n_4_net__40_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__40_ : 1'b0;
  assign n_4_net__39_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__39_ : 1'b0;
  assign n_4_net__38_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__38_ : 1'b0;
  assign n_4_net__37_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__37_ : 1'b0;
  assign n_4_net__36_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__36_ : 1'b0;
  assign n_4_net__35_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__35_ : 1'b0;
  assign n_4_net__34_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__34_ : 1'b0;
  assign n_4_net__33_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__33_ : 1'b0;
  assign n_4_net__32_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__32_ : 1'b0;
  assign n_4_net__31_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__31_ : 1'b0;
  assign n_4_net__30_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__30_ : 1'b0;
  assign n_4_net__29_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__29_ : 1'b0;
  assign n_4_net__28_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__28_ : 1'b0;
  assign n_4_net__27_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__27_ : 1'b0;
  assign n_4_net__26_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__26_ : 1'b0;
  assign n_4_net__25_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__25_ : 1'b0;
  assign n_4_net__24_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__24_ : 1'b0;
  assign n_4_net__23_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__23_ : 1'b0;
  assign n_4_net__22_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__22_ : 1'b0;
  assign n_4_net__21_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__21_ : 1'b0;
  assign n_4_net__20_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__20_ : 1'b0;
  assign n_4_net__19_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__19_ : 1'b0;
  assign n_4_net__18_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__18_ : 1'b0;
  assign n_4_net__17_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__17_ : 1'b0;
  assign n_4_net__16_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__16_ : 1'b0;
  assign n_4_net__15_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__15_ : 1'b0;
  assign n_4_net__14_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__14_ : 1'b0;
  assign n_4_net__13_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__13_ : 1'b0;
  assign n_4_net__12_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__12_ : 1'b0;
  assign n_4_net__11_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__11_ : 1'b0;
  assign n_4_net__10_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__10_ : 1'b0;
  assign n_4_net__9_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__9_ : 1'b0;
  assign n_4_net__8_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__8_ : 1'b0;
  assign n_4_net__7_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__7_ : 1'b0;
  assign n_4_net__6_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__6_ : 1'b0;
  assign n_4_net__5_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__5_ : 1'b0;
  assign n_4_net__4_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__4_ : 1'b0;
  assign n_4_net__3_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__3_ : 1'b0;
  assign n_4_net__2_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__2_ : 1'b0;
  assign n_4_net__1_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__1_ : 1'b0;
  assign n_4_net__0_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__0_ : 1'b0;
  assign n_0_net_ = reset | N179;
  assign n_5_net_ = reset | N184;

endmodule



module bsg_assembler_out
(
  clk,
  reset,
  calibration_done_i,
  valid_i,
  data_i,
  ready_o,
  in_top_channel_i,
  out_top_channel_i,
  valid_o,
  data_o,
  ready_i
);

  input [639:0] data_i;
  input [3:0] in_top_channel_i;
  input [3:0] out_top_channel_i;
  output [9:0] valid_o;
  output [639:0] data_o;
  input [9:0] ready_i;
  input clk;
  input reset;
  input calibration_done_i;
  input valid_i;
  output ready_o;
  wire [9:0] valid_o,fifo_not_full_vec,fifo_valid_vec,fifo_deq_vec;
  wire [639:0] data_o,fifo_data_vec;
  wire ready_o,n_0_net_,n_1_net_,n_2_net_,n_3_net_,n_4_net_,n_5_net_,n_6_net_,n_7_net_,
  n_8_net_,n_9_net_,N0,N1,N2,N3,N4,N5,N6,N7,N8;

  bsg_two_fifo_width_p64_ready_THEN_valid_p1
  fifos_0__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[0]),
    .data_i(data_i[63:0]),
    .v_i(n_0_net_),
    .v_o(fifo_valid_vec[0]),
    .data_o(fifo_data_vec[63:0]),
    .yumi_i(fifo_deq_vec[0])
  );


  bsg_two_fifo_width_p64_ready_THEN_valid_p1
  fifos_1__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[1]),
    .data_i(data_i[127:64]),
    .v_i(n_1_net_),
    .v_o(fifo_valid_vec[1]),
    .data_o(fifo_data_vec[127:64]),
    .yumi_i(fifo_deq_vec[1])
  );


  bsg_two_fifo_width_p64_ready_THEN_valid_p1
  fifos_2__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[2]),
    .data_i(data_i[191:128]),
    .v_i(n_2_net_),
    .v_o(fifo_valid_vec[2]),
    .data_o(fifo_data_vec[191:128]),
    .yumi_i(fifo_deq_vec[2])
  );


  bsg_two_fifo_width_p64_ready_THEN_valid_p1
  fifos_3__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[3]),
    .data_i(data_i[255:192]),
    .v_i(n_3_net_),
    .v_o(fifo_valid_vec[3]),
    .data_o(fifo_data_vec[255:192]),
    .yumi_i(fifo_deq_vec[3])
  );


  bsg_two_fifo_width_p64_ready_THEN_valid_p1
  fifos_4__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[4]),
    .data_i(data_i[319:256]),
    .v_i(n_4_net_),
    .v_o(fifo_valid_vec[4]),
    .data_o(fifo_data_vec[319:256]),
    .yumi_i(fifo_deq_vec[4])
  );


  bsg_two_fifo_width_p64_ready_THEN_valid_p1
  fifos_5__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[5]),
    .data_i(data_i[383:320]),
    .v_i(n_5_net_),
    .v_o(fifo_valid_vec[5]),
    .data_o(fifo_data_vec[383:320]),
    .yumi_i(fifo_deq_vec[5])
  );


  bsg_two_fifo_width_p64_ready_THEN_valid_p1
  fifos_6__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[6]),
    .data_i(data_i[447:384]),
    .v_i(n_6_net_),
    .v_o(fifo_valid_vec[6]),
    .data_o(fifo_data_vec[447:384]),
    .yumi_i(fifo_deq_vec[6])
  );


  bsg_two_fifo_width_p64_ready_THEN_valid_p1
  fifos_7__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[7]),
    .data_i(data_i[511:448]),
    .v_i(n_7_net_),
    .v_o(fifo_valid_vec[7]),
    .data_o(fifo_data_vec[511:448]),
    .yumi_i(fifo_deq_vec[7])
  );


  bsg_two_fifo_width_p64_ready_THEN_valid_p1
  fifos_8__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[8]),
    .data_i(data_i[575:512]),
    .v_i(n_8_net_),
    .v_o(fifo_valid_vec[8]),
    .data_o(fifo_data_vec[575:512]),
    .yumi_i(fifo_deq_vec[8])
  );


  bsg_two_fifo_width_p64_ready_THEN_valid_p1
  fifos_9__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[9]),
    .data_i(data_i[639:576]),
    .v_i(n_9_net_),
    .v_o(fifo_valid_vec[9]),
    .data_o(fifo_data_vec[639:576]),
    .yumi_i(fifo_deq_vec[9])
  );


  bsg_round_robin_fifo_to_fifo_width_p64_num_in_p10_num_out_p10_out_channel_count_mask_p512
  rr_fifo_to_fifo
  (
    .clk(clk),
    .reset(reset),
    .valid_i(fifo_valid_vec),
    .data_i(fifo_data_vec),
    .yumi_o(fifo_deq_vec),
    .in_top_channel_i(in_top_channel_i),
    .out_top_channel_i(out_top_channel_i),
    .valid_o(valid_o),
    .data_o(data_o),
    .ready_i(ready_i)
  );

  assign ready_o = N8 & calibration_done_i;
  assign N8 = N7 & fifo_not_full_vec[0];
  assign N7 = N6 & fifo_not_full_vec[1];
  assign N6 = N5 & fifo_not_full_vec[2];
  assign N5 = N4 & fifo_not_full_vec[3];
  assign N4 = N3 & fifo_not_full_vec[4];
  assign N3 = N2 & fifo_not_full_vec[5];
  assign N2 = N1 & fifo_not_full_vec[6];
  assign N1 = N0 & fifo_not_full_vec[7];
  assign N0 = fifo_not_full_vec[9] & fifo_not_full_vec[8];
  assign n_0_net_ = valid_i & ready_o;
  assign n_1_net_ = valid_i & ready_o;
  assign n_2_net_ = valid_i & ready_o;
  assign n_3_net_ = valid_i & ready_o;
  assign n_4_net_ = valid_i & ready_o;
  assign n_5_net_ = valid_i & ready_o;
  assign n_6_net_ = valid_i & ready_o;
  assign n_7_net_ = valid_i & ready_o;
  assign n_8_net_ = valid_i & ready_o;
  assign n_9_net_ = valid_i & ready_o;

endmodule

