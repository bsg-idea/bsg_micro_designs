

module top
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  o
);

  input [127:0] a_i;
  input [127:0] b_i;
  output [255:0] o;
  input clk_i;
  input rst_i;
  input v_i;

  bsg_mul_array
  wrapper
  (
    .a_i(a_i),
    .b_i(b_i),
    .o(o),
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i)
  );


endmodule



module bsg_and_width_p128
(
  a_i,
  b_i,
  o
);

  input [127:0] a_i;
  input [127:0] b_i;
  output [127:0] o;
  wire [127:0] o;
  assign o[127] = a_i[127] & b_i[127];
  assign o[126] = a_i[126] & b_i[126];
  assign o[125] = a_i[125] & b_i[125];
  assign o[124] = a_i[124] & b_i[124];
  assign o[123] = a_i[123] & b_i[123];
  assign o[122] = a_i[122] & b_i[122];
  assign o[121] = a_i[121] & b_i[121];
  assign o[120] = a_i[120] & b_i[120];
  assign o[119] = a_i[119] & b_i[119];
  assign o[118] = a_i[118] & b_i[118];
  assign o[117] = a_i[117] & b_i[117];
  assign o[116] = a_i[116] & b_i[116];
  assign o[115] = a_i[115] & b_i[115];
  assign o[114] = a_i[114] & b_i[114];
  assign o[113] = a_i[113] & b_i[113];
  assign o[112] = a_i[112] & b_i[112];
  assign o[111] = a_i[111] & b_i[111];
  assign o[110] = a_i[110] & b_i[110];
  assign o[109] = a_i[109] & b_i[109];
  assign o[108] = a_i[108] & b_i[108];
  assign o[107] = a_i[107] & b_i[107];
  assign o[106] = a_i[106] & b_i[106];
  assign o[105] = a_i[105] & b_i[105];
  assign o[104] = a_i[104] & b_i[104];
  assign o[103] = a_i[103] & b_i[103];
  assign o[102] = a_i[102] & b_i[102];
  assign o[101] = a_i[101] & b_i[101];
  assign o[100] = a_i[100] & b_i[100];
  assign o[99] = a_i[99] & b_i[99];
  assign o[98] = a_i[98] & b_i[98];
  assign o[97] = a_i[97] & b_i[97];
  assign o[96] = a_i[96] & b_i[96];
  assign o[95] = a_i[95] & b_i[95];
  assign o[94] = a_i[94] & b_i[94];
  assign o[93] = a_i[93] & b_i[93];
  assign o[92] = a_i[92] & b_i[92];
  assign o[91] = a_i[91] & b_i[91];
  assign o[90] = a_i[90] & b_i[90];
  assign o[89] = a_i[89] & b_i[89];
  assign o[88] = a_i[88] & b_i[88];
  assign o[87] = a_i[87] & b_i[87];
  assign o[86] = a_i[86] & b_i[86];
  assign o[85] = a_i[85] & b_i[85];
  assign o[84] = a_i[84] & b_i[84];
  assign o[83] = a_i[83] & b_i[83];
  assign o[82] = a_i[82] & b_i[82];
  assign o[81] = a_i[81] & b_i[81];
  assign o[80] = a_i[80] & b_i[80];
  assign o[79] = a_i[79] & b_i[79];
  assign o[78] = a_i[78] & b_i[78];
  assign o[77] = a_i[77] & b_i[77];
  assign o[76] = a_i[76] & b_i[76];
  assign o[75] = a_i[75] & b_i[75];
  assign o[74] = a_i[74] & b_i[74];
  assign o[73] = a_i[73] & b_i[73];
  assign o[72] = a_i[72] & b_i[72];
  assign o[71] = a_i[71] & b_i[71];
  assign o[70] = a_i[70] & b_i[70];
  assign o[69] = a_i[69] & b_i[69];
  assign o[68] = a_i[68] & b_i[68];
  assign o[67] = a_i[67] & b_i[67];
  assign o[66] = a_i[66] & b_i[66];
  assign o[65] = a_i[65] & b_i[65];
  assign o[64] = a_i[64] & b_i[64];
  assign o[63] = a_i[63] & b_i[63];
  assign o[62] = a_i[62] & b_i[62];
  assign o[61] = a_i[61] & b_i[61];
  assign o[60] = a_i[60] & b_i[60];
  assign o[59] = a_i[59] & b_i[59];
  assign o[58] = a_i[58] & b_i[58];
  assign o[57] = a_i[57] & b_i[57];
  assign o[56] = a_i[56] & b_i[56];
  assign o[55] = a_i[55] & b_i[55];
  assign o[54] = a_i[54] & b_i[54];
  assign o[53] = a_i[53] & b_i[53];
  assign o[52] = a_i[52] & b_i[52];
  assign o[51] = a_i[51] & b_i[51];
  assign o[50] = a_i[50] & b_i[50];
  assign o[49] = a_i[49] & b_i[49];
  assign o[48] = a_i[48] & b_i[48];
  assign o[47] = a_i[47] & b_i[47];
  assign o[46] = a_i[46] & b_i[46];
  assign o[45] = a_i[45] & b_i[45];
  assign o[44] = a_i[44] & b_i[44];
  assign o[43] = a_i[43] & b_i[43];
  assign o[42] = a_i[42] & b_i[42];
  assign o[41] = a_i[41] & b_i[41];
  assign o[40] = a_i[40] & b_i[40];
  assign o[39] = a_i[39] & b_i[39];
  assign o[38] = a_i[38] & b_i[38];
  assign o[37] = a_i[37] & b_i[37];
  assign o[36] = a_i[36] & b_i[36];
  assign o[35] = a_i[35] & b_i[35];
  assign o[34] = a_i[34] & b_i[34];
  assign o[33] = a_i[33] & b_i[33];
  assign o[32] = a_i[32] & b_i[32];
  assign o[31] = a_i[31] & b_i[31];
  assign o[30] = a_i[30] & b_i[30];
  assign o[29] = a_i[29] & b_i[29];
  assign o[28] = a_i[28] & b_i[28];
  assign o[27] = a_i[27] & b_i[27];
  assign o[26] = a_i[26] & b_i[26];
  assign o[25] = a_i[25] & b_i[25];
  assign o[24] = a_i[24] & b_i[24];
  assign o[23] = a_i[23] & b_i[23];
  assign o[22] = a_i[22] & b_i[22];
  assign o[21] = a_i[21] & b_i[21];
  assign o[20] = a_i[20] & b_i[20];
  assign o[19] = a_i[19] & b_i[19];
  assign o[18] = a_i[18] & b_i[18];
  assign o[17] = a_i[17] & b_i[17];
  assign o[16] = a_i[16] & b_i[16];
  assign o[15] = a_i[15] & b_i[15];
  assign o[14] = a_i[14] & b_i[14];
  assign o[13] = a_i[13] & b_i[13];
  assign o[12] = a_i[12] & b_i[12];
  assign o[11] = a_i[11] & b_i[11];
  assign o[10] = a_i[10] & b_i[10];
  assign o[9] = a_i[9] & b_i[9];
  assign o[8] = a_i[8] & b_i[8];
  assign o[7] = a_i[7] & b_i[7];
  assign o[6] = a_i[6] & b_i[6];
  assign o[5] = a_i[5] & b_i[5];
  assign o[4] = a_i[4] & b_i[4];
  assign o[3] = a_i[3] & b_i[3];
  assign o[2] = a_i[2] & b_i[2];
  assign o[1] = a_i[1] & b_i[1];
  assign o[0] = a_i[0] & b_i[0];

endmodule



module bsg_adder_ripple_carry_width_p128
(
  a_i,
  b_i,
  s_o,
  c_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  output [127:0] s_o;
  output c_o;
  wire [127:0] s_o;
  wire c_o;
  assign { c_o, s_o } = a_i + b_i;

endmodule



module bsg_mul_array_row_128_0_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [0:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [1:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [1:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[1] = s_o[0];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1], b_i[1:1] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_1_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [1:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [2:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [2:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[2] = s_o[0];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2], b_i[2:2] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_2_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [2:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [3:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [3:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[3] = s_o[0];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3], b_i[3:3] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_3_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [3:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [4:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [4:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[4] = s_o[0];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4], b_i[4:4] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_4_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [4:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [5:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [5:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[5] = s_o[0];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5], b_i[5:5] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_5_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [5:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [6:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [6:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[6] = s_o[0];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6], b_i[6:6] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_6_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [6:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [7:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [7:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[7] = s_o[0];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7], b_i[7:7] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_7_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [7:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [8:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [8:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[8] = s_o[0];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8], b_i[8:8] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_8_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [8:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [9:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [9:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[9] = s_o[0];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9], b_i[9:9] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_9_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [9:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [10:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [10:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[10] = s_o[0];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10], b_i[10:10] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_10_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [10:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [11:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [11:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[11] = s_o[0];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11], b_i[11:11] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_11_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [11:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [12:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [12:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[12] = s_o[0];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12], b_i[12:12] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_12_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [12:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [13:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [13:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[13] = s_o[0];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13], b_i[13:13] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_13_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [13:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [14:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [14:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[14] = s_o[0];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14], b_i[14:14] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_14_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [14:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [15:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [15:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[15] = s_o[0];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15], b_i[15:15] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_15_1
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [15:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [16:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire N0,N1,pc,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,
  N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,
  N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,
  N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,
  N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,
  N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,
  N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,
  N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
  N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,
  N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,
  N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,
  N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,
  N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,
  N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,
  N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,
  N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,
  N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,
  N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,
  N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,
  N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,
  N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,
  N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415;
  wire [127:0] pp,ps;
  reg [16:0] prod_accum_o;
  reg [127:0] a_o,b_o,s_o;
  reg c_o;

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16], b_i[16:16] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(ps),
    .c_o(pc)
  );

  assign { N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N1)? a_i : 1'b0;
  assign N0 = rst_i;
  assign N1 = N2;
  assign { N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1)? b_i : 1'b0;
  assign { N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1)? ps : 1'b0;
  assign N387 = (N0)? 1'b0 : 
                (N1)? pc : 1'b0;
  assign { N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                    (N1)? { ps[0:0], prod_accum_i } : 1'b0;
  assign N2 = ~rst_i;
  assign N405 = ~v_i;
  assign N406 = N405 & N2;
  assign N407 = ~N406;
  assign N408 = N405 & N2;
  assign N409 = ~N408;
  assign N410 = N405 & N2;
  assign N411 = ~N410;
  assign N412 = N405 & N2;
  assign N413 = ~N412;
  assign N414 = N405 & N2;
  assign N415 = ~N414;

  always @(posedge clk_i) begin
    if(N407) begin
      { prod_accum_o[16:16] } <= { N404 };
      { s_o[97:0] } <= { N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259 };
      c_o <= N387;
    end 
    if(N409) begin
      { prod_accum_o[15:15] } <= { N403 };
      { b_o[68:0] } <= { N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131 };
      { s_o[127:98] } <= { N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357 };
    end 
    if(N411) begin
      { prod_accum_o[14:14] } <= { N402 };
      { a_o[39:0] } <= { N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3 };
      { b_o[127:69] } <= { N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200 };
    end 
    if(N413) begin
      { prod_accum_o[13:13], prod_accum_o[10:0] } <= { N401, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388 };
      { a_o[127:40] } <= { N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43 };
    end 
    if(N415) begin
      { prod_accum_o[12:11] } <= { N400, N399 };
    end 
  end


endmodule



module bsg_mul_array_row_128_16_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [16:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [17:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [17:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[17] = s_o[0];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17], b_i[17:17] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_17_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [17:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [18:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [18:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[18] = s_o[0];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18], b_i[18:18] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_18_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [18:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [19:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [19:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[19] = s_o[0];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19], b_i[19:19] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_19_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [19:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [20:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [20:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[20] = s_o[0];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20], b_i[20:20] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_20_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [20:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [21:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [21:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[21] = s_o[0];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21], b_i[21:21] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_21_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [21:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [22:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [22:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[22] = s_o[0];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22], b_i[22:22] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_22_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [22:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [23:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [23:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[23] = s_o[0];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23], b_i[23:23] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_23_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [23:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [24:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [24:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[24] = s_o[0];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24], b_i[24:24] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_24_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [24:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [25:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [25:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[25] = s_o[0];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25], b_i[25:25] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_25_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [25:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [26:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [26:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[26] = s_o[0];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26], b_i[26:26] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_26_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [26:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [27:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [27:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[27] = s_o[0];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27], b_i[27:27] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_27_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [27:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [28:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [28:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[28] = s_o[0];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28], b_i[28:28] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_28_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [28:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [29:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [29:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[29] = s_o[0];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29], b_i[29:29] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_29_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [29:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [30:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [30:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[30] = s_o[0];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30], b_i[30:30] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_30_0
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [30:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [31:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [31:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[31] = s_o[0];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31], b_i[31:31] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_31_1
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [31:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [32:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire N0,N1,pc,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,
  N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,
  N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,
  N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,
  N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,
  N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,
  N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,
  N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
  N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,
  N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,
  N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,
  N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,
  N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,
  N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,
  N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,
  N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,
  N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,
  N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,
  N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,
  N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,
  N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,
  N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,
  N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431;
  wire [127:0] pp,ps;
  reg [32:0] prod_accum_o;
  reg [127:0] a_o,b_o,s_o;
  reg c_o;

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32], b_i[32:32] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(ps),
    .c_o(pc)
  );

  assign { N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N1)? a_i : 1'b0;
  assign N0 = rst_i;
  assign N1 = N2;
  assign { N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1)? b_i : 1'b0;
  assign { N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1)? ps : 1'b0;
  assign N387 = (N0)? 1'b0 : 
                (N1)? pc : 1'b0;
  assign { N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                    (N1)? { ps[0:0], prod_accum_i } : 1'b0;
  assign N2 = ~rst_i;
  assign N421 = ~v_i;
  assign N422 = N421 & N2;
  assign N423 = ~N422;
  assign N424 = N421 & N2;
  assign N425 = ~N424;
  assign N426 = N421 & N2;
  assign N427 = ~N426;
  assign N428 = N421 & N2;
  assign N429 = ~N428;
  assign N430 = N421 & N2;
  assign N431 = ~N430;

  always @(posedge clk_i) begin
    if(N423) begin
      { prod_accum_o[32:32] } <= { N420 };
      { s_o[97:0] } <= { N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259 };
      c_o <= N387;
    end 
    if(N425) begin
      { prod_accum_o[31:31] } <= { N419 };
      { b_o[68:0] } <= { N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131 };
      { s_o[127:98] } <= { N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357 };
    end 
    if(N427) begin
      { prod_accum_o[30:30] } <= { N418 };
      { a_o[39:0] } <= { N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3 };
      { b_o[127:69] } <= { N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200 };
    end 
    if(N429) begin
      { prod_accum_o[29:29], prod_accum_o[10:0] } <= { N417, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388 };
      { a_o[127:40] } <= { N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43 };
    end 
    if(N431) begin
      { prod_accum_o[28:11] } <= { N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399 };
    end 
  end


endmodule



module bsg_mul_array_row_128_32_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [32:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [33:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [33:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[33] = s_o[0];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33], b_i[33:33] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_33_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [33:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [34:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [34:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[34] = s_o[0];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34], b_i[34:34] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_34_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [34:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [35:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [35:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[35] = s_o[0];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35], b_i[35:35] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_35_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [35:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [36:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [36:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[36] = s_o[0];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36], b_i[36:36] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_36_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [36:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [37:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [37:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[37] = s_o[0];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37], b_i[37:37] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_37_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [37:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [38:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [38:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[38] = s_o[0];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38], b_i[38:38] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_38_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [38:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [39:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [39:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[39] = s_o[0];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39], b_i[39:39] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_39_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [39:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [40:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [40:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[40] = s_o[0];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40], b_i[40:40] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_40_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [40:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [41:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [41:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[41] = s_o[0];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41], b_i[41:41] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_41_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [41:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [42:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [42:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[42] = s_o[0];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42], b_i[42:42] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_42_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [42:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [43:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [43:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[43] = s_o[0];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43], b_i[43:43] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_43_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [43:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [44:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [44:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[44] = s_o[0];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44], b_i[44:44] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_44_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [44:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [45:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [45:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[45] = s_o[0];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45], b_i[45:45] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_45_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [45:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [46:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [46:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[46] = s_o[0];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46], b_i[46:46] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_46_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [46:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [47:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [47:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[47] = s_o[0];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47], b_i[47:47] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_47_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [47:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [48:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [48:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[48] = s_o[0];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48], b_i[48:48] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_48_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [48:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [49:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [49:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[49] = s_o[0];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49], b_i[49:49] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_49_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [49:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [50:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [50:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[50] = s_o[0];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50], b_i[50:50] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_50_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [50:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [51:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [51:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[51] = s_o[0];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51], b_i[51:51] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_51_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [51:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [52:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [52:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[52] = s_o[0];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52], b_i[52:52] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_52_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [52:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [53:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [53:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[53] = s_o[0];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53], b_i[53:53] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_53_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [53:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [54:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [54:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[54] = s_o[0];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54], b_i[54:54] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_54_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [54:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [55:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [55:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[55] = s_o[0];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55], b_i[55:55] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_55_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [55:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [56:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [56:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[56] = s_o[0];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56], b_i[56:56] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_56_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [56:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [57:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [57:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[57] = s_o[0];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57], b_i[57:57] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_57_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [57:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [58:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [58:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[58] = s_o[0];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58], b_i[58:58] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_58_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [58:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [59:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [59:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[59] = s_o[0];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59], b_i[59:59] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_59_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [59:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [60:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [60:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[60] = s_o[0];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60], b_i[60:60] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_60_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [60:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [61:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [61:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[61] = s_o[0];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61], b_i[61:61] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_61_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [61:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [62:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [62:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[62] = s_o[0];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62], b_i[62:62] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_62_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [62:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [63:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [63:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[63] = s_o[0];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63], b_i[63:63] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_63_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [63:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [64:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [64:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[64] = s_o[0];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64], b_i[64:64] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_64_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [64:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [65:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [65:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[65] = s_o[0];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65], b_i[65:65] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_65_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [65:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [66:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [66:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[66] = s_o[0];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66], b_i[66:66] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_66_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [66:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [67:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [67:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[67] = s_o[0];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67], b_i[67:67] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_67_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [67:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [68:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [68:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[68] = s_o[0];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68], b_i[68:68] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_68_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [68:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [69:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [69:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[69] = s_o[0];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69], b_i[69:69] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_69_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [69:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [70:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [70:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[70] = s_o[0];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70], b_i[70:70] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_70_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [70:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [71:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [71:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[71] = s_o[0];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71], b_i[71:71] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_71_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [71:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [72:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [72:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[72] = s_o[0];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72], b_i[72:72] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_72_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [72:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [73:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [73:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[73] = s_o[0];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73], b_i[73:73] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_73_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [73:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [74:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [74:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[74] = s_o[0];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74], b_i[74:74] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_74_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [74:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [75:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [75:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[75] = s_o[0];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75], b_i[75:75] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_75_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [75:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [76:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [76:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[76] = s_o[0];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76], b_i[76:76] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_76_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [76:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [77:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [77:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[77] = s_o[0];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77], b_i[77:77] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_77_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [77:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [78:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [78:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[78] = s_o[0];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78], b_i[78:78] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_78_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [78:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [79:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [79:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[79] = s_o[0];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79], b_i[79:79] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_79_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [79:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [80:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [80:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[80] = s_o[0];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80], b_i[80:80] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_80_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [80:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [81:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [81:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[81] = s_o[0];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81], b_i[81:81] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_81_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [81:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [82:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [82:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[82] = s_o[0];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82], b_i[82:82] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_82_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [82:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [83:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [83:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[83] = s_o[0];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83], b_i[83:83] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_83_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [83:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [84:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [84:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[84] = s_o[0];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84], b_i[84:84] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_84_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [84:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [85:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [85:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[85] = s_o[0];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85], b_i[85:85] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_85_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [85:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [86:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [86:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[86] = s_o[0];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86], b_i[86:86] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_86_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [86:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [87:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [87:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[87] = s_o[0];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87], b_i[87:87] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_87_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [87:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [88:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [88:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[88] = s_o[0];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88], b_i[88:88] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_88_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [88:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [89:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [89:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[89] = s_o[0];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89], b_i[89:89] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_89_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [89:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [90:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [90:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[90] = s_o[0];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90], b_i[90:90] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_90_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [90:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [91:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [91:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[91] = s_o[0];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91], b_i[91:91] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_91_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [91:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [92:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [92:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[92] = s_o[0];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92], b_i[92:92] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_92_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [92:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [93:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [93:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[93] = s_o[0];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93], b_i[93:93] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_93_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [93:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [94:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [94:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[94] = s_o[0];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94], b_i[94:94] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_94_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [94:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [95:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [95:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[95] = s_o[0];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95], b_i[95:95] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_95_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [95:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [96:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [96:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[96] = s_o[0];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96], b_i[96:96] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_96_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [96:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [97:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [97:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[97] = s_o[0];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97], b_i[97:97] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_97_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [97:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [98:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [98:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[98] = s_o[0];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98], b_i[98:98] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_98_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [98:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [99:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [99:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[99] = s_o[0];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99], b_i[99:99] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_99_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [99:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [100:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [100:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[100] = s_o[0];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100], b_i[100:100] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_100_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [100:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [101:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [101:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[101] = s_o[0];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101], b_i[101:101] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_101_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [101:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [102:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [102:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[102] = s_o[0];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102], b_i[102:102] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_102_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [102:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [103:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [103:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[103] = s_o[0];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103], b_i[103:103] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_103_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [103:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [104:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [104:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[104] = s_o[0];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104], b_i[104:104] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_104_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [104:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [105:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [105:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[105] = s_o[0];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105], b_i[105:105] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_105_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [105:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [106:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [106:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[106] = s_o[0];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106], b_i[106:106] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_106_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [106:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [107:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [107:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[107] = s_o[0];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107], b_i[107:107] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_107_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [107:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [108:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [108:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[108] = s_o[0];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108], b_i[108:108] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_108_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [108:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [109:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [109:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[109] = s_o[0];
  assign prod_accum_o[108] = prod_accum_i[108];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109], b_i[109:109] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_109_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [109:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [110:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [110:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[110] = s_o[0];
  assign prod_accum_o[109] = prod_accum_i[109];
  assign prod_accum_o[108] = prod_accum_i[108];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110], b_i[110:110] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_110_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [110:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [111:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [111:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[111] = s_o[0];
  assign prod_accum_o[110] = prod_accum_i[110];
  assign prod_accum_o[109] = prod_accum_i[109];
  assign prod_accum_o[108] = prod_accum_i[108];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111], b_i[111:111] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_111_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [111:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [112:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [112:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[112] = s_o[0];
  assign prod_accum_o[111] = prod_accum_i[111];
  assign prod_accum_o[110] = prod_accum_i[110];
  assign prod_accum_o[109] = prod_accum_i[109];
  assign prod_accum_o[108] = prod_accum_i[108];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112], b_i[112:112] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_112_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [112:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [113:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [113:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[113] = s_o[0];
  assign prod_accum_o[112] = prod_accum_i[112];
  assign prod_accum_o[111] = prod_accum_i[111];
  assign prod_accum_o[110] = prod_accum_i[110];
  assign prod_accum_o[109] = prod_accum_i[109];
  assign prod_accum_o[108] = prod_accum_i[108];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113], b_i[113:113] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_113_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [113:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [114:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [114:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[114] = s_o[0];
  assign prod_accum_o[113] = prod_accum_i[113];
  assign prod_accum_o[112] = prod_accum_i[112];
  assign prod_accum_o[111] = prod_accum_i[111];
  assign prod_accum_o[110] = prod_accum_i[110];
  assign prod_accum_o[109] = prod_accum_i[109];
  assign prod_accum_o[108] = prod_accum_i[108];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114], b_i[114:114] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_114_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [114:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [115:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [115:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[115] = s_o[0];
  assign prod_accum_o[114] = prod_accum_i[114];
  assign prod_accum_o[113] = prod_accum_i[113];
  assign prod_accum_o[112] = prod_accum_i[112];
  assign prod_accum_o[111] = prod_accum_i[111];
  assign prod_accum_o[110] = prod_accum_i[110];
  assign prod_accum_o[109] = prod_accum_i[109];
  assign prod_accum_o[108] = prod_accum_i[108];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115], b_i[115:115] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_115_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [115:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [116:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [116:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[116] = s_o[0];
  assign prod_accum_o[115] = prod_accum_i[115];
  assign prod_accum_o[114] = prod_accum_i[114];
  assign prod_accum_o[113] = prod_accum_i[113];
  assign prod_accum_o[112] = prod_accum_i[112];
  assign prod_accum_o[111] = prod_accum_i[111];
  assign prod_accum_o[110] = prod_accum_i[110];
  assign prod_accum_o[109] = prod_accum_i[109];
  assign prod_accum_o[108] = prod_accum_i[108];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116], b_i[116:116] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_116_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [116:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [117:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [117:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[117] = s_o[0];
  assign prod_accum_o[116] = prod_accum_i[116];
  assign prod_accum_o[115] = prod_accum_i[115];
  assign prod_accum_o[114] = prod_accum_i[114];
  assign prod_accum_o[113] = prod_accum_i[113];
  assign prod_accum_o[112] = prod_accum_i[112];
  assign prod_accum_o[111] = prod_accum_i[111];
  assign prod_accum_o[110] = prod_accum_i[110];
  assign prod_accum_o[109] = prod_accum_i[109];
  assign prod_accum_o[108] = prod_accum_i[108];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117], b_i[117:117] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_117_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [117:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [118:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [118:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[118] = s_o[0];
  assign prod_accum_o[117] = prod_accum_i[117];
  assign prod_accum_o[116] = prod_accum_i[116];
  assign prod_accum_o[115] = prod_accum_i[115];
  assign prod_accum_o[114] = prod_accum_i[114];
  assign prod_accum_o[113] = prod_accum_i[113];
  assign prod_accum_o[112] = prod_accum_i[112];
  assign prod_accum_o[111] = prod_accum_i[111];
  assign prod_accum_o[110] = prod_accum_i[110];
  assign prod_accum_o[109] = prod_accum_i[109];
  assign prod_accum_o[108] = prod_accum_i[108];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118], b_i[118:118] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_118_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [118:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [119:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [119:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[119] = s_o[0];
  assign prod_accum_o[118] = prod_accum_i[118];
  assign prod_accum_o[117] = prod_accum_i[117];
  assign prod_accum_o[116] = prod_accum_i[116];
  assign prod_accum_o[115] = prod_accum_i[115];
  assign prod_accum_o[114] = prod_accum_i[114];
  assign prod_accum_o[113] = prod_accum_i[113];
  assign prod_accum_o[112] = prod_accum_i[112];
  assign prod_accum_o[111] = prod_accum_i[111];
  assign prod_accum_o[110] = prod_accum_i[110];
  assign prod_accum_o[109] = prod_accum_i[109];
  assign prod_accum_o[108] = prod_accum_i[108];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119], b_i[119:119] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_119_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [119:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [120:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [120:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[120] = s_o[0];
  assign prod_accum_o[119] = prod_accum_i[119];
  assign prod_accum_o[118] = prod_accum_i[118];
  assign prod_accum_o[117] = prod_accum_i[117];
  assign prod_accum_o[116] = prod_accum_i[116];
  assign prod_accum_o[115] = prod_accum_i[115];
  assign prod_accum_o[114] = prod_accum_i[114];
  assign prod_accum_o[113] = prod_accum_i[113];
  assign prod_accum_o[112] = prod_accum_i[112];
  assign prod_accum_o[111] = prod_accum_i[111];
  assign prod_accum_o[110] = prod_accum_i[110];
  assign prod_accum_o[109] = prod_accum_i[109];
  assign prod_accum_o[108] = prod_accum_i[108];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120], b_i[120:120] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_120_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [120:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [121:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [121:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[121] = s_o[0];
  assign prod_accum_o[120] = prod_accum_i[120];
  assign prod_accum_o[119] = prod_accum_i[119];
  assign prod_accum_o[118] = prod_accum_i[118];
  assign prod_accum_o[117] = prod_accum_i[117];
  assign prod_accum_o[116] = prod_accum_i[116];
  assign prod_accum_o[115] = prod_accum_i[115];
  assign prod_accum_o[114] = prod_accum_i[114];
  assign prod_accum_o[113] = prod_accum_i[113];
  assign prod_accum_o[112] = prod_accum_i[112];
  assign prod_accum_o[111] = prod_accum_i[111];
  assign prod_accum_o[110] = prod_accum_i[110];
  assign prod_accum_o[109] = prod_accum_i[109];
  assign prod_accum_o[108] = prod_accum_i[108];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121], b_i[121:121] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_121_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [121:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [122:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [122:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[122] = s_o[0];
  assign prod_accum_o[121] = prod_accum_i[121];
  assign prod_accum_o[120] = prod_accum_i[120];
  assign prod_accum_o[119] = prod_accum_i[119];
  assign prod_accum_o[118] = prod_accum_i[118];
  assign prod_accum_o[117] = prod_accum_i[117];
  assign prod_accum_o[116] = prod_accum_i[116];
  assign prod_accum_o[115] = prod_accum_i[115];
  assign prod_accum_o[114] = prod_accum_i[114];
  assign prod_accum_o[113] = prod_accum_i[113];
  assign prod_accum_o[112] = prod_accum_i[112];
  assign prod_accum_o[111] = prod_accum_i[111];
  assign prod_accum_o[110] = prod_accum_i[110];
  assign prod_accum_o[109] = prod_accum_i[109];
  assign prod_accum_o[108] = prod_accum_i[108];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122], b_i[122:122] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_122_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [122:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [123:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [123:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[123] = s_o[0];
  assign prod_accum_o[122] = prod_accum_i[122];
  assign prod_accum_o[121] = prod_accum_i[121];
  assign prod_accum_o[120] = prod_accum_i[120];
  assign prod_accum_o[119] = prod_accum_i[119];
  assign prod_accum_o[118] = prod_accum_i[118];
  assign prod_accum_o[117] = prod_accum_i[117];
  assign prod_accum_o[116] = prod_accum_i[116];
  assign prod_accum_o[115] = prod_accum_i[115];
  assign prod_accum_o[114] = prod_accum_i[114];
  assign prod_accum_o[113] = prod_accum_i[113];
  assign prod_accum_o[112] = prod_accum_i[112];
  assign prod_accum_o[111] = prod_accum_i[111];
  assign prod_accum_o[110] = prod_accum_i[110];
  assign prod_accum_o[109] = prod_accum_i[109];
  assign prod_accum_o[108] = prod_accum_i[108];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123], b_i[123:123] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_123_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [123:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [124:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [124:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[124] = s_o[0];
  assign prod_accum_o[123] = prod_accum_i[123];
  assign prod_accum_o[122] = prod_accum_i[122];
  assign prod_accum_o[121] = prod_accum_i[121];
  assign prod_accum_o[120] = prod_accum_i[120];
  assign prod_accum_o[119] = prod_accum_i[119];
  assign prod_accum_o[118] = prod_accum_i[118];
  assign prod_accum_o[117] = prod_accum_i[117];
  assign prod_accum_o[116] = prod_accum_i[116];
  assign prod_accum_o[115] = prod_accum_i[115];
  assign prod_accum_o[114] = prod_accum_i[114];
  assign prod_accum_o[113] = prod_accum_i[113];
  assign prod_accum_o[112] = prod_accum_i[112];
  assign prod_accum_o[111] = prod_accum_i[111];
  assign prod_accum_o[110] = prod_accum_i[110];
  assign prod_accum_o[109] = prod_accum_i[109];
  assign prod_accum_o[108] = prod_accum_i[108];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124], b_i[124:124] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_124_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [124:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [125:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [125:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[125] = s_o[0];
  assign prod_accum_o[124] = prod_accum_i[124];
  assign prod_accum_o[123] = prod_accum_i[123];
  assign prod_accum_o[122] = prod_accum_i[122];
  assign prod_accum_o[121] = prod_accum_i[121];
  assign prod_accum_o[120] = prod_accum_i[120];
  assign prod_accum_o[119] = prod_accum_i[119];
  assign prod_accum_o[118] = prod_accum_i[118];
  assign prod_accum_o[117] = prod_accum_i[117];
  assign prod_accum_o[116] = prod_accum_i[116];
  assign prod_accum_o[115] = prod_accum_i[115];
  assign prod_accum_o[114] = prod_accum_i[114];
  assign prod_accum_o[113] = prod_accum_i[113];
  assign prod_accum_o[112] = prod_accum_i[112];
  assign prod_accum_o[111] = prod_accum_i[111];
  assign prod_accum_o[110] = prod_accum_i[110];
  assign prod_accum_o[109] = prod_accum_i[109];
  assign prod_accum_o[108] = prod_accum_i[108];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125], b_i[125:125] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_125_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [125:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [126:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,pp;
  wire [126:0] prod_accum_o;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[126] = s_o[0];
  assign prod_accum_o[125] = prod_accum_i[125];
  assign prod_accum_o[124] = prod_accum_i[124];
  assign prod_accum_o[123] = prod_accum_i[123];
  assign prod_accum_o[122] = prod_accum_i[122];
  assign prod_accum_o[121] = prod_accum_i[121];
  assign prod_accum_o[120] = prod_accum_i[120];
  assign prod_accum_o[119] = prod_accum_i[119];
  assign prod_accum_o[118] = prod_accum_i[118];
  assign prod_accum_o[117] = prod_accum_i[117];
  assign prod_accum_o[116] = prod_accum_i[116];
  assign prod_accum_o[115] = prod_accum_i[115];
  assign prod_accum_o[114] = prod_accum_i[114];
  assign prod_accum_o[113] = prod_accum_i[113];
  assign prod_accum_o[112] = prod_accum_i[112];
  assign prod_accum_o[111] = prod_accum_i[111];
  assign prod_accum_o[110] = prod_accum_i[110];
  assign prod_accum_o[109] = prod_accum_i[109];
  assign prod_accum_o[108] = prod_accum_i[108];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126], b_i[126:126] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array_row_128_126_x
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  s_i,
  c_i,
  prod_accum_i,
  a_o,
  b_o,
  s_o,
  c_o,
  prod_accum_o
);

  input [127:0] a_i;
  input [127:0] b_i;
  input [127:0] s_i;
  input [126:0] prod_accum_i;
  output [127:0] a_o;
  output [127:0] b_o;
  output [127:0] s_o;
  output [127:0] prod_accum_o;
  input clk_i;
  input rst_i;
  input v_i;
  input c_i;
  output c_o;
  wire [127:0] a_o,b_o,s_o,prod_accum_o,pp;
  wire c_o;
  assign a_o[127] = a_i[127];
  assign a_o[126] = a_i[126];
  assign a_o[125] = a_i[125];
  assign a_o[124] = a_i[124];
  assign a_o[123] = a_i[123];
  assign a_o[122] = a_i[122];
  assign a_o[121] = a_i[121];
  assign a_o[120] = a_i[120];
  assign a_o[119] = a_i[119];
  assign a_o[118] = a_i[118];
  assign a_o[117] = a_i[117];
  assign a_o[116] = a_i[116];
  assign a_o[115] = a_i[115];
  assign a_o[114] = a_i[114];
  assign a_o[113] = a_i[113];
  assign a_o[112] = a_i[112];
  assign a_o[111] = a_i[111];
  assign a_o[110] = a_i[110];
  assign a_o[109] = a_i[109];
  assign a_o[108] = a_i[108];
  assign a_o[107] = a_i[107];
  assign a_o[106] = a_i[106];
  assign a_o[105] = a_i[105];
  assign a_o[104] = a_i[104];
  assign a_o[103] = a_i[103];
  assign a_o[102] = a_i[102];
  assign a_o[101] = a_i[101];
  assign a_o[100] = a_i[100];
  assign a_o[99] = a_i[99];
  assign a_o[98] = a_i[98];
  assign a_o[97] = a_i[97];
  assign a_o[96] = a_i[96];
  assign a_o[95] = a_i[95];
  assign a_o[94] = a_i[94];
  assign a_o[93] = a_i[93];
  assign a_o[92] = a_i[92];
  assign a_o[91] = a_i[91];
  assign a_o[90] = a_i[90];
  assign a_o[89] = a_i[89];
  assign a_o[88] = a_i[88];
  assign a_o[87] = a_i[87];
  assign a_o[86] = a_i[86];
  assign a_o[85] = a_i[85];
  assign a_o[84] = a_i[84];
  assign a_o[83] = a_i[83];
  assign a_o[82] = a_i[82];
  assign a_o[81] = a_i[81];
  assign a_o[80] = a_i[80];
  assign a_o[79] = a_i[79];
  assign a_o[78] = a_i[78];
  assign a_o[77] = a_i[77];
  assign a_o[76] = a_i[76];
  assign a_o[75] = a_i[75];
  assign a_o[74] = a_i[74];
  assign a_o[73] = a_i[73];
  assign a_o[72] = a_i[72];
  assign a_o[71] = a_i[71];
  assign a_o[70] = a_i[70];
  assign a_o[69] = a_i[69];
  assign a_o[68] = a_i[68];
  assign a_o[67] = a_i[67];
  assign a_o[66] = a_i[66];
  assign a_o[65] = a_i[65];
  assign a_o[64] = a_i[64];
  assign a_o[63] = a_i[63];
  assign a_o[62] = a_i[62];
  assign a_o[61] = a_i[61];
  assign a_o[60] = a_i[60];
  assign a_o[59] = a_i[59];
  assign a_o[58] = a_i[58];
  assign a_o[57] = a_i[57];
  assign a_o[56] = a_i[56];
  assign a_o[55] = a_i[55];
  assign a_o[54] = a_i[54];
  assign a_o[53] = a_i[53];
  assign a_o[52] = a_i[52];
  assign a_o[51] = a_i[51];
  assign a_o[50] = a_i[50];
  assign a_o[49] = a_i[49];
  assign a_o[48] = a_i[48];
  assign a_o[47] = a_i[47];
  assign a_o[46] = a_i[46];
  assign a_o[45] = a_i[45];
  assign a_o[44] = a_i[44];
  assign a_o[43] = a_i[43];
  assign a_o[42] = a_i[42];
  assign a_o[41] = a_i[41];
  assign a_o[40] = a_i[40];
  assign a_o[39] = a_i[39];
  assign a_o[38] = a_i[38];
  assign a_o[37] = a_i[37];
  assign a_o[36] = a_i[36];
  assign a_o[35] = a_i[35];
  assign a_o[34] = a_i[34];
  assign a_o[33] = a_i[33];
  assign a_o[32] = a_i[32];
  assign a_o[31] = a_i[31];
  assign a_o[30] = a_i[30];
  assign a_o[29] = a_i[29];
  assign a_o[28] = a_i[28];
  assign a_o[27] = a_i[27];
  assign a_o[26] = a_i[26];
  assign a_o[25] = a_i[25];
  assign a_o[24] = a_i[24];
  assign a_o[23] = a_i[23];
  assign a_o[22] = a_i[22];
  assign a_o[21] = a_i[21];
  assign a_o[20] = a_i[20];
  assign a_o[19] = a_i[19];
  assign a_o[18] = a_i[18];
  assign a_o[17] = a_i[17];
  assign a_o[16] = a_i[16];
  assign a_o[15] = a_i[15];
  assign a_o[14] = a_i[14];
  assign a_o[13] = a_i[13];
  assign a_o[12] = a_i[12];
  assign a_o[11] = a_i[11];
  assign a_o[10] = a_i[10];
  assign a_o[9] = a_i[9];
  assign a_o[8] = a_i[8];
  assign a_o[7] = a_i[7];
  assign a_o[6] = a_i[6];
  assign a_o[5] = a_i[5];
  assign a_o[4] = a_i[4];
  assign a_o[3] = a_i[3];
  assign a_o[2] = a_i[2];
  assign a_o[1] = a_i[1];
  assign a_o[0] = a_i[0];
  assign b_o[127] = b_i[127];
  assign b_o[126] = b_i[126];
  assign b_o[125] = b_i[125];
  assign b_o[124] = b_i[124];
  assign b_o[123] = b_i[123];
  assign b_o[122] = b_i[122];
  assign b_o[121] = b_i[121];
  assign b_o[120] = b_i[120];
  assign b_o[119] = b_i[119];
  assign b_o[118] = b_i[118];
  assign b_o[117] = b_i[117];
  assign b_o[116] = b_i[116];
  assign b_o[115] = b_i[115];
  assign b_o[114] = b_i[114];
  assign b_o[113] = b_i[113];
  assign b_o[112] = b_i[112];
  assign b_o[111] = b_i[111];
  assign b_o[110] = b_i[110];
  assign b_o[109] = b_i[109];
  assign b_o[108] = b_i[108];
  assign b_o[107] = b_i[107];
  assign b_o[106] = b_i[106];
  assign b_o[105] = b_i[105];
  assign b_o[104] = b_i[104];
  assign b_o[103] = b_i[103];
  assign b_o[102] = b_i[102];
  assign b_o[101] = b_i[101];
  assign b_o[100] = b_i[100];
  assign b_o[99] = b_i[99];
  assign b_o[98] = b_i[98];
  assign b_o[97] = b_i[97];
  assign b_o[96] = b_i[96];
  assign b_o[95] = b_i[95];
  assign b_o[94] = b_i[94];
  assign b_o[93] = b_i[93];
  assign b_o[92] = b_i[92];
  assign b_o[91] = b_i[91];
  assign b_o[90] = b_i[90];
  assign b_o[89] = b_i[89];
  assign b_o[88] = b_i[88];
  assign b_o[87] = b_i[87];
  assign b_o[86] = b_i[86];
  assign b_o[85] = b_i[85];
  assign b_o[84] = b_i[84];
  assign b_o[83] = b_i[83];
  assign b_o[82] = b_i[82];
  assign b_o[81] = b_i[81];
  assign b_o[80] = b_i[80];
  assign b_o[79] = b_i[79];
  assign b_o[78] = b_i[78];
  assign b_o[77] = b_i[77];
  assign b_o[76] = b_i[76];
  assign b_o[75] = b_i[75];
  assign b_o[74] = b_i[74];
  assign b_o[73] = b_i[73];
  assign b_o[72] = b_i[72];
  assign b_o[71] = b_i[71];
  assign b_o[70] = b_i[70];
  assign b_o[69] = b_i[69];
  assign b_o[68] = b_i[68];
  assign b_o[67] = b_i[67];
  assign b_o[66] = b_i[66];
  assign b_o[65] = b_i[65];
  assign b_o[64] = b_i[64];
  assign b_o[63] = b_i[63];
  assign b_o[62] = b_i[62];
  assign b_o[61] = b_i[61];
  assign b_o[60] = b_i[60];
  assign b_o[59] = b_i[59];
  assign b_o[58] = b_i[58];
  assign b_o[57] = b_i[57];
  assign b_o[56] = b_i[56];
  assign b_o[55] = b_i[55];
  assign b_o[54] = b_i[54];
  assign b_o[53] = b_i[53];
  assign b_o[52] = b_i[52];
  assign b_o[51] = b_i[51];
  assign b_o[50] = b_i[50];
  assign b_o[49] = b_i[49];
  assign b_o[48] = b_i[48];
  assign b_o[47] = b_i[47];
  assign b_o[46] = b_i[46];
  assign b_o[45] = b_i[45];
  assign b_o[44] = b_i[44];
  assign b_o[43] = b_i[43];
  assign b_o[42] = b_i[42];
  assign b_o[41] = b_i[41];
  assign b_o[40] = b_i[40];
  assign b_o[39] = b_i[39];
  assign b_o[38] = b_i[38];
  assign b_o[37] = b_i[37];
  assign b_o[36] = b_i[36];
  assign b_o[35] = b_i[35];
  assign b_o[34] = b_i[34];
  assign b_o[33] = b_i[33];
  assign b_o[32] = b_i[32];
  assign b_o[31] = b_i[31];
  assign b_o[30] = b_i[30];
  assign b_o[29] = b_i[29];
  assign b_o[28] = b_i[28];
  assign b_o[27] = b_i[27];
  assign b_o[26] = b_i[26];
  assign b_o[25] = b_i[25];
  assign b_o[24] = b_i[24];
  assign b_o[23] = b_i[23];
  assign b_o[22] = b_i[22];
  assign b_o[21] = b_i[21];
  assign b_o[20] = b_i[20];
  assign b_o[19] = b_i[19];
  assign b_o[18] = b_i[18];
  assign b_o[17] = b_i[17];
  assign b_o[16] = b_i[16];
  assign b_o[15] = b_i[15];
  assign b_o[14] = b_i[14];
  assign b_o[13] = b_i[13];
  assign b_o[12] = b_i[12];
  assign b_o[11] = b_i[11];
  assign b_o[10] = b_i[10];
  assign b_o[9] = b_i[9];
  assign b_o[8] = b_i[8];
  assign b_o[7] = b_i[7];
  assign b_o[6] = b_i[6];
  assign b_o[5] = b_i[5];
  assign b_o[4] = b_i[4];
  assign b_o[3] = b_i[3];
  assign b_o[2] = b_i[2];
  assign b_o[1] = b_i[1];
  assign b_o[0] = b_i[0];
  assign prod_accum_o[127] = s_o[0];
  assign prod_accum_o[126] = prod_accum_i[126];
  assign prod_accum_o[125] = prod_accum_i[125];
  assign prod_accum_o[124] = prod_accum_i[124];
  assign prod_accum_o[123] = prod_accum_i[123];
  assign prod_accum_o[122] = prod_accum_i[122];
  assign prod_accum_o[121] = prod_accum_i[121];
  assign prod_accum_o[120] = prod_accum_i[120];
  assign prod_accum_o[119] = prod_accum_i[119];
  assign prod_accum_o[118] = prod_accum_i[118];
  assign prod_accum_o[117] = prod_accum_i[117];
  assign prod_accum_o[116] = prod_accum_i[116];
  assign prod_accum_o[115] = prod_accum_i[115];
  assign prod_accum_o[114] = prod_accum_i[114];
  assign prod_accum_o[113] = prod_accum_i[113];
  assign prod_accum_o[112] = prod_accum_i[112];
  assign prod_accum_o[111] = prod_accum_i[111];
  assign prod_accum_o[110] = prod_accum_i[110];
  assign prod_accum_o[109] = prod_accum_i[109];
  assign prod_accum_o[108] = prod_accum_i[108];
  assign prod_accum_o[107] = prod_accum_i[107];
  assign prod_accum_o[106] = prod_accum_i[106];
  assign prod_accum_o[105] = prod_accum_i[105];
  assign prod_accum_o[104] = prod_accum_i[104];
  assign prod_accum_o[103] = prod_accum_i[103];
  assign prod_accum_o[102] = prod_accum_i[102];
  assign prod_accum_o[101] = prod_accum_i[101];
  assign prod_accum_o[100] = prod_accum_i[100];
  assign prod_accum_o[99] = prod_accum_i[99];
  assign prod_accum_o[98] = prod_accum_i[98];
  assign prod_accum_o[97] = prod_accum_i[97];
  assign prod_accum_o[96] = prod_accum_i[96];
  assign prod_accum_o[95] = prod_accum_i[95];
  assign prod_accum_o[94] = prod_accum_i[94];
  assign prod_accum_o[93] = prod_accum_i[93];
  assign prod_accum_o[92] = prod_accum_i[92];
  assign prod_accum_o[91] = prod_accum_i[91];
  assign prod_accum_o[90] = prod_accum_i[90];
  assign prod_accum_o[89] = prod_accum_i[89];
  assign prod_accum_o[88] = prod_accum_i[88];
  assign prod_accum_o[87] = prod_accum_i[87];
  assign prod_accum_o[86] = prod_accum_i[86];
  assign prod_accum_o[85] = prod_accum_i[85];
  assign prod_accum_o[84] = prod_accum_i[84];
  assign prod_accum_o[83] = prod_accum_i[83];
  assign prod_accum_o[82] = prod_accum_i[82];
  assign prod_accum_o[81] = prod_accum_i[81];
  assign prod_accum_o[80] = prod_accum_i[80];
  assign prod_accum_o[79] = prod_accum_i[79];
  assign prod_accum_o[78] = prod_accum_i[78];
  assign prod_accum_o[77] = prod_accum_i[77];
  assign prod_accum_o[76] = prod_accum_i[76];
  assign prod_accum_o[75] = prod_accum_i[75];
  assign prod_accum_o[74] = prod_accum_i[74];
  assign prod_accum_o[73] = prod_accum_i[73];
  assign prod_accum_o[72] = prod_accum_i[72];
  assign prod_accum_o[71] = prod_accum_i[71];
  assign prod_accum_o[70] = prod_accum_i[70];
  assign prod_accum_o[69] = prod_accum_i[69];
  assign prod_accum_o[68] = prod_accum_i[68];
  assign prod_accum_o[67] = prod_accum_i[67];
  assign prod_accum_o[66] = prod_accum_i[66];
  assign prod_accum_o[65] = prod_accum_i[65];
  assign prod_accum_o[64] = prod_accum_i[64];
  assign prod_accum_o[63] = prod_accum_i[63];
  assign prod_accum_o[62] = prod_accum_i[62];
  assign prod_accum_o[61] = prod_accum_i[61];
  assign prod_accum_o[60] = prod_accum_i[60];
  assign prod_accum_o[59] = prod_accum_i[59];
  assign prod_accum_o[58] = prod_accum_i[58];
  assign prod_accum_o[57] = prod_accum_i[57];
  assign prod_accum_o[56] = prod_accum_i[56];
  assign prod_accum_o[55] = prod_accum_i[55];
  assign prod_accum_o[54] = prod_accum_i[54];
  assign prod_accum_o[53] = prod_accum_i[53];
  assign prod_accum_o[52] = prod_accum_i[52];
  assign prod_accum_o[51] = prod_accum_i[51];
  assign prod_accum_o[50] = prod_accum_i[50];
  assign prod_accum_o[49] = prod_accum_i[49];
  assign prod_accum_o[48] = prod_accum_i[48];
  assign prod_accum_o[47] = prod_accum_i[47];
  assign prod_accum_o[46] = prod_accum_i[46];
  assign prod_accum_o[45] = prod_accum_i[45];
  assign prod_accum_o[44] = prod_accum_i[44];
  assign prod_accum_o[43] = prod_accum_i[43];
  assign prod_accum_o[42] = prod_accum_i[42];
  assign prod_accum_o[41] = prod_accum_i[41];
  assign prod_accum_o[40] = prod_accum_i[40];
  assign prod_accum_o[39] = prod_accum_i[39];
  assign prod_accum_o[38] = prod_accum_i[38];
  assign prod_accum_o[37] = prod_accum_i[37];
  assign prod_accum_o[36] = prod_accum_i[36];
  assign prod_accum_o[35] = prod_accum_i[35];
  assign prod_accum_o[34] = prod_accum_i[34];
  assign prod_accum_o[33] = prod_accum_i[33];
  assign prod_accum_o[32] = prod_accum_i[32];
  assign prod_accum_o[31] = prod_accum_i[31];
  assign prod_accum_o[30] = prod_accum_i[30];
  assign prod_accum_o[29] = prod_accum_i[29];
  assign prod_accum_o[28] = prod_accum_i[28];
  assign prod_accum_o[27] = prod_accum_i[27];
  assign prod_accum_o[26] = prod_accum_i[26];
  assign prod_accum_o[25] = prod_accum_i[25];
  assign prod_accum_o[24] = prod_accum_i[24];
  assign prod_accum_o[23] = prod_accum_i[23];
  assign prod_accum_o[22] = prod_accum_i[22];
  assign prod_accum_o[21] = prod_accum_i[21];
  assign prod_accum_o[20] = prod_accum_i[20];
  assign prod_accum_o[19] = prod_accum_i[19];
  assign prod_accum_o[18] = prod_accum_i[18];
  assign prod_accum_o[17] = prod_accum_i[17];
  assign prod_accum_o[16] = prod_accum_i[16];
  assign prod_accum_o[15] = prod_accum_i[15];
  assign prod_accum_o[14] = prod_accum_i[14];
  assign prod_accum_o[13] = prod_accum_i[13];
  assign prod_accum_o[12] = prod_accum_i[12];
  assign prod_accum_o[11] = prod_accum_i[11];
  assign prod_accum_o[10] = prod_accum_i[10];
  assign prod_accum_o[9] = prod_accum_i[9];
  assign prod_accum_o[8] = prod_accum_i[8];
  assign prod_accum_o[7] = prod_accum_i[7];
  assign prod_accum_o[6] = prod_accum_i[6];
  assign prod_accum_o[5] = prod_accum_i[5];
  assign prod_accum_o[4] = prod_accum_i[4];
  assign prod_accum_o[3] = prod_accum_i[3];
  assign prod_accum_o[2] = prod_accum_i[2];
  assign prod_accum_o[1] = prod_accum_i[1];
  assign prod_accum_o[0] = prod_accum_i[0];

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127], b_i[127:127] }),
    .o(pp)
  );


  bsg_adder_ripple_carry_width_p128
  adder0
  (
    .a_i(pp),
    .b_i({ c_i, s_i[127:1] }),
    .s_o(s_o),
    .c_o(c_o)
  );


endmodule



module bsg_mul_array
(
  clk_i,
  rst_i,
  v_i,
  a_i,
  b_i,
  o
);

  input [127:0] a_i;
  input [127:0] b_i;
  output [255:0] o;
  input clk_i;
  input rst_i;
  input v_i;
  wire [255:0] o;
  wire s_r_2__127_,s_r_2__126_,s_r_2__125_,s_r_2__124_,s_r_2__123_,s_r_2__122_,
  s_r_2__121_,s_r_2__120_,s_r_2__119_,s_r_2__118_,s_r_2__117_,s_r_2__116_,s_r_2__115_,
  s_r_2__114_,s_r_2__113_,s_r_2__112_,s_r_2__111_,s_r_2__110_,s_r_2__109_,s_r_2__108_,
  s_r_2__107_,s_r_2__106_,s_r_2__105_,s_r_2__104_,s_r_2__103_,s_r_2__102_,
  s_r_2__101_,s_r_2__100_,s_r_2__99_,s_r_2__98_,s_r_2__97_,s_r_2__96_,s_r_2__95_,
  s_r_2__94_,s_r_2__93_,s_r_2__92_,s_r_2__91_,s_r_2__90_,s_r_2__89_,s_r_2__88_,s_r_2__87_,
  s_r_2__86_,s_r_2__85_,s_r_2__84_,s_r_2__83_,s_r_2__82_,s_r_2__81_,s_r_2__80_,
  s_r_2__79_,s_r_2__78_,s_r_2__77_,s_r_2__76_,s_r_2__75_,s_r_2__74_,s_r_2__73_,
  s_r_2__72_,s_r_2__71_,s_r_2__70_,s_r_2__69_,s_r_2__68_,s_r_2__67_,s_r_2__66_,
  s_r_2__65_,s_r_2__64_,s_r_2__63_,s_r_2__62_,s_r_2__61_,s_r_2__60_,s_r_2__59_,s_r_2__58_,
  s_r_2__57_,s_r_2__56_,s_r_2__55_,s_r_2__54_,s_r_2__53_,s_r_2__52_,s_r_2__51_,
  s_r_2__50_,s_r_2__49_,s_r_2__48_,s_r_2__47_,s_r_2__46_,s_r_2__45_,s_r_2__44_,
  s_r_2__43_,s_r_2__42_,s_r_2__41_,s_r_2__40_,s_r_2__39_,s_r_2__38_,s_r_2__37_,s_r_2__36_,
  s_r_2__35_,s_r_2__34_,s_r_2__33_,s_r_2__32_,s_r_2__31_,s_r_2__30_,s_r_2__29_,
  s_r_2__28_,s_r_2__27_,s_r_2__26_,s_r_2__25_,s_r_2__24_,s_r_2__23_,s_r_2__22_,
  s_r_2__21_,s_r_2__20_,s_r_2__19_,s_r_2__18_,s_r_2__17_,s_r_2__16_,s_r_2__15_,
  s_r_2__14_,s_r_2__13_,s_r_2__12_,s_r_2__11_,s_r_2__10_,s_r_2__9_,s_r_2__8_,s_r_2__7_,
  s_r_2__6_,s_r_2__5_,s_r_2__4_,s_r_2__3_,s_r_2__2_,s_r_2__1_,s_r_2__0_,s_r_1__127_,
  s_r_1__126_,s_r_1__125_,s_r_1__124_,s_r_1__123_,s_r_1__122_,s_r_1__121_,
  s_r_1__120_,s_r_1__119_,s_r_1__118_,s_r_1__117_,s_r_1__116_,s_r_1__115_,s_r_1__114_,
  s_r_1__113_,s_r_1__112_,s_r_1__111_,s_r_1__110_,s_r_1__109_,s_r_1__108_,s_r_1__107_,
  s_r_1__106_,s_r_1__105_,s_r_1__104_,s_r_1__103_,s_r_1__102_,s_r_1__101_,
  s_r_1__100_,s_r_1__99_,s_r_1__98_,s_r_1__97_,s_r_1__96_,s_r_1__95_,s_r_1__94_,s_r_1__93_,
  s_r_1__92_,s_r_1__91_,s_r_1__90_,s_r_1__89_,s_r_1__88_,s_r_1__87_,s_r_1__86_,
  s_r_1__85_,s_r_1__84_,s_r_1__83_,s_r_1__82_,s_r_1__81_,s_r_1__80_,s_r_1__79_,
  s_r_1__78_,s_r_1__77_,s_r_1__76_,s_r_1__75_,s_r_1__74_,s_r_1__73_,s_r_1__72_,
  s_r_1__71_,s_r_1__70_,s_r_1__69_,s_r_1__68_,s_r_1__67_,s_r_1__66_,s_r_1__65_,s_r_1__64_,
  s_r_1__63_,s_r_1__62_,s_r_1__61_,s_r_1__60_,s_r_1__59_,s_r_1__58_,s_r_1__57_,
  s_r_1__56_,s_r_1__55_,s_r_1__54_,s_r_1__53_,s_r_1__52_,s_r_1__51_,s_r_1__50_,
  s_r_1__49_,s_r_1__48_,s_r_1__47_,s_r_1__46_,s_r_1__45_,s_r_1__44_,s_r_1__43_,s_r_1__42_,
  s_r_1__41_,s_r_1__40_,s_r_1__39_,s_r_1__38_,s_r_1__37_,s_r_1__36_,s_r_1__35_,
  s_r_1__34_,s_r_1__33_,s_r_1__32_,s_r_1__31_,s_r_1__30_,s_r_1__29_,s_r_1__28_,
  s_r_1__27_,s_r_1__26_,s_r_1__25_,s_r_1__24_,s_r_1__23_,s_r_1__22_,s_r_1__21_,
  s_r_1__20_,s_r_1__19_,s_r_1__18_,s_r_1__17_,s_r_1__16_,s_r_1__15_,s_r_1__14_,s_r_1__13_,
  s_r_1__12_,s_r_1__11_,s_r_1__10_,s_r_1__9_,s_r_1__8_,s_r_1__7_,s_r_1__6_,
  s_r_1__5_,s_r_1__4_,s_r_1__3_,s_r_1__2_,s_r_1__1_,s_r_1__0_,s_r_0__127_,s_r_0__126_,
  s_r_0__125_,s_r_0__124_,s_r_0__123_,s_r_0__122_,s_r_0__121_,s_r_0__120_,s_r_0__119_,
  s_r_0__118_,s_r_0__117_,s_r_0__116_,s_r_0__115_,s_r_0__114_,s_r_0__113_,
  s_r_0__112_,s_r_0__111_,s_r_0__110_,s_r_0__109_,s_r_0__108_,s_r_0__107_,s_r_0__106_,
  s_r_0__105_,s_r_0__104_,s_r_0__103_,s_r_0__102_,s_r_0__101_,s_r_0__100_,s_r_0__99_,
  s_r_0__98_,s_r_0__97_,s_r_0__96_,s_r_0__95_,s_r_0__94_,s_r_0__93_,s_r_0__92_,
  s_r_0__91_,s_r_0__90_,s_r_0__89_,s_r_0__88_,s_r_0__87_,s_r_0__86_,s_r_0__85_,
  s_r_0__84_,s_r_0__83_,s_r_0__82_,s_r_0__81_,s_r_0__80_,s_r_0__79_,s_r_0__78_,
  s_r_0__77_,s_r_0__76_,s_r_0__75_,s_r_0__74_,s_r_0__73_,s_r_0__72_,s_r_0__71_,s_r_0__70_,
  s_r_0__69_,s_r_0__68_,s_r_0__67_,s_r_0__66_,s_r_0__65_,s_r_0__64_,s_r_0__63_,
  s_r_0__62_,s_r_0__61_,s_r_0__60_,s_r_0__59_,s_r_0__58_,s_r_0__57_,s_r_0__56_,
  s_r_0__55_,s_r_0__54_,s_r_0__53_,s_r_0__52_,s_r_0__51_,s_r_0__50_,s_r_0__49_,s_r_0__48_,
  s_r_0__47_,s_r_0__46_,s_r_0__45_,s_r_0__44_,s_r_0__43_,s_r_0__42_,s_r_0__41_,
  s_r_0__40_,s_r_0__39_,s_r_0__38_,s_r_0__37_,s_r_0__36_,s_r_0__35_,s_r_0__34_,
  s_r_0__33_,s_r_0__32_,s_r_0__31_,s_r_0__30_,s_r_0__29_,s_r_0__28_,s_r_0__27_,
  s_r_0__26_,s_r_0__25_,s_r_0__24_,s_r_0__23_,s_r_0__22_,s_r_0__21_,s_r_0__20_,s_r_0__19_,
  s_r_0__18_,s_r_0__17_,s_r_0__16_,s_r_0__15_,s_r_0__14_,s_r_0__13_,s_r_0__12_,
  s_r_0__11_,s_r_0__10_,s_r_0__9_,s_r_0__8_,s_r_0__7_,s_r_0__6_,s_r_0__5_,s_r_0__4_,
  s_r_0__3_,s_r_0__2_,s_r_0__1_,s_r_0__0_,prod_accum_2__3_,prod_accum_2__2_,
  prod_accum_2__1_,prod_accum_2__0_,prod_accum_1__2_,prod_accum_1__1_,prod_accum_1__0_,
  prod_accum_0__1_,prod_accum_0__0_,s_r_6__127_,s_r_6__126_,s_r_6__125_,s_r_6__124_,
  s_r_6__123_,s_r_6__122_,s_r_6__121_,s_r_6__120_,s_r_6__119_,s_r_6__118_,
  s_r_6__117_,s_r_6__116_,s_r_6__115_,s_r_6__114_,s_r_6__113_,s_r_6__112_,s_r_6__111_,
  s_r_6__110_,s_r_6__109_,s_r_6__108_,s_r_6__107_,s_r_6__106_,s_r_6__105_,s_r_6__104_,
  s_r_6__103_,s_r_6__102_,s_r_6__101_,s_r_6__100_,s_r_6__99_,s_r_6__98_,s_r_6__97_,
  s_r_6__96_,s_r_6__95_,s_r_6__94_,s_r_6__93_,s_r_6__92_,s_r_6__91_,s_r_6__90_,
  s_r_6__89_,s_r_6__88_,s_r_6__87_,s_r_6__86_,s_r_6__85_,s_r_6__84_,s_r_6__83_,
  s_r_6__82_,s_r_6__81_,s_r_6__80_,s_r_6__79_,s_r_6__78_,s_r_6__77_,s_r_6__76_,
  s_r_6__75_,s_r_6__74_,s_r_6__73_,s_r_6__72_,s_r_6__71_,s_r_6__70_,s_r_6__69_,s_r_6__68_,
  s_r_6__67_,s_r_6__66_,s_r_6__65_,s_r_6__64_,s_r_6__63_,s_r_6__62_,s_r_6__61_,
  s_r_6__60_,s_r_6__59_,s_r_6__58_,s_r_6__57_,s_r_6__56_,s_r_6__55_,s_r_6__54_,
  s_r_6__53_,s_r_6__52_,s_r_6__51_,s_r_6__50_,s_r_6__49_,s_r_6__48_,s_r_6__47_,
  s_r_6__46_,s_r_6__45_,s_r_6__44_,s_r_6__43_,s_r_6__42_,s_r_6__41_,s_r_6__40_,s_r_6__39_,
  s_r_6__38_,s_r_6__37_,s_r_6__36_,s_r_6__35_,s_r_6__34_,s_r_6__33_,s_r_6__32_,
  s_r_6__31_,s_r_6__30_,s_r_6__29_,s_r_6__28_,s_r_6__27_,s_r_6__26_,s_r_6__25_,
  s_r_6__24_,s_r_6__23_,s_r_6__22_,s_r_6__21_,s_r_6__20_,s_r_6__19_,s_r_6__18_,s_r_6__17_,
  s_r_6__16_,s_r_6__15_,s_r_6__14_,s_r_6__13_,s_r_6__12_,s_r_6__11_,s_r_6__10_,
  s_r_6__9_,s_r_6__8_,s_r_6__7_,s_r_6__6_,s_r_6__5_,s_r_6__4_,s_r_6__3_,s_r_6__2_,
  s_r_6__1_,s_r_6__0_,s_r_5__127_,s_r_5__126_,s_r_5__125_,s_r_5__124_,s_r_5__123_,
  s_r_5__122_,s_r_5__121_,s_r_5__120_,s_r_5__119_,s_r_5__118_,s_r_5__117_,
  s_r_5__116_,s_r_5__115_,s_r_5__114_,s_r_5__113_,s_r_5__112_,s_r_5__111_,s_r_5__110_,
  s_r_5__109_,s_r_5__108_,s_r_5__107_,s_r_5__106_,s_r_5__105_,s_r_5__104_,s_r_5__103_,
  s_r_5__102_,s_r_5__101_,s_r_5__100_,s_r_5__99_,s_r_5__98_,s_r_5__97_,s_r_5__96_,
  s_r_5__95_,s_r_5__94_,s_r_5__93_,s_r_5__92_,s_r_5__91_,s_r_5__90_,s_r_5__89_,
  s_r_5__88_,s_r_5__87_,s_r_5__86_,s_r_5__85_,s_r_5__84_,s_r_5__83_,s_r_5__82_,
  s_r_5__81_,s_r_5__80_,s_r_5__79_,s_r_5__78_,s_r_5__77_,s_r_5__76_,s_r_5__75_,s_r_5__74_,
  s_r_5__73_,s_r_5__72_,s_r_5__71_,s_r_5__70_,s_r_5__69_,s_r_5__68_,s_r_5__67_,
  s_r_5__66_,s_r_5__65_,s_r_5__64_,s_r_5__63_,s_r_5__62_,s_r_5__61_,s_r_5__60_,
  s_r_5__59_,s_r_5__58_,s_r_5__57_,s_r_5__56_,s_r_5__55_,s_r_5__54_,s_r_5__53_,
  s_r_5__52_,s_r_5__51_,s_r_5__50_,s_r_5__49_,s_r_5__48_,s_r_5__47_,s_r_5__46_,s_r_5__45_,
  s_r_5__44_,s_r_5__43_,s_r_5__42_,s_r_5__41_,s_r_5__40_,s_r_5__39_,s_r_5__38_,
  s_r_5__37_,s_r_5__36_,s_r_5__35_,s_r_5__34_,s_r_5__33_,s_r_5__32_,s_r_5__31_,
  s_r_5__30_,s_r_5__29_,s_r_5__28_,s_r_5__27_,s_r_5__26_,s_r_5__25_,s_r_5__24_,s_r_5__23_,
  s_r_5__22_,s_r_5__21_,s_r_5__20_,s_r_5__19_,s_r_5__18_,s_r_5__17_,s_r_5__16_,
  s_r_5__15_,s_r_5__14_,s_r_5__13_,s_r_5__12_,s_r_5__11_,s_r_5__10_,s_r_5__9_,
  s_r_5__8_,s_r_5__7_,s_r_5__6_,s_r_5__5_,s_r_5__4_,s_r_5__3_,s_r_5__2_,s_r_5__1_,
  s_r_5__0_,s_r_4__127_,s_r_4__126_,s_r_4__125_,s_r_4__124_,s_r_4__123_,s_r_4__122_,
  s_r_4__121_,s_r_4__120_,s_r_4__119_,s_r_4__118_,s_r_4__117_,s_r_4__116_,s_r_4__115_,
  s_r_4__114_,s_r_4__113_,s_r_4__112_,s_r_4__111_,s_r_4__110_,s_r_4__109_,
  s_r_4__108_,s_r_4__107_,s_r_4__106_,s_r_4__105_,s_r_4__104_,s_r_4__103_,s_r_4__102_,
  s_r_4__101_,s_r_4__100_,s_r_4__99_,s_r_4__98_,s_r_4__97_,s_r_4__96_,s_r_4__95_,
  s_r_4__94_,s_r_4__93_,s_r_4__92_,s_r_4__91_,s_r_4__90_,s_r_4__89_,s_r_4__88_,
  s_r_4__87_,s_r_4__86_,s_r_4__85_,s_r_4__84_,s_r_4__83_,s_r_4__82_,s_r_4__81_,s_r_4__80_,
  s_r_4__79_,s_r_4__78_,s_r_4__77_,s_r_4__76_,s_r_4__75_,s_r_4__74_,s_r_4__73_,
  s_r_4__72_,s_r_4__71_,s_r_4__70_,s_r_4__69_,s_r_4__68_,s_r_4__67_,s_r_4__66_,
  s_r_4__65_,s_r_4__64_,s_r_4__63_,s_r_4__62_,s_r_4__61_,s_r_4__60_,s_r_4__59_,
  s_r_4__58_,s_r_4__57_,s_r_4__56_,s_r_4__55_,s_r_4__54_,s_r_4__53_,s_r_4__52_,s_r_4__51_,
  s_r_4__50_,s_r_4__49_,s_r_4__48_,s_r_4__47_,s_r_4__46_,s_r_4__45_,s_r_4__44_,
  s_r_4__43_,s_r_4__42_,s_r_4__41_,s_r_4__40_,s_r_4__39_,s_r_4__38_,s_r_4__37_,
  s_r_4__36_,s_r_4__35_,s_r_4__34_,s_r_4__33_,s_r_4__32_,s_r_4__31_,s_r_4__30_,s_r_4__29_,
  s_r_4__28_,s_r_4__27_,s_r_4__26_,s_r_4__25_,s_r_4__24_,s_r_4__23_,s_r_4__22_,
  s_r_4__21_,s_r_4__20_,s_r_4__19_,s_r_4__18_,s_r_4__17_,s_r_4__16_,s_r_4__15_,
  s_r_4__14_,s_r_4__13_,s_r_4__12_,s_r_4__11_,s_r_4__10_,s_r_4__9_,s_r_4__8_,s_r_4__7_,
  s_r_4__6_,s_r_4__5_,s_r_4__4_,s_r_4__3_,s_r_4__2_,s_r_4__1_,s_r_4__0_,
  s_r_3__127_,s_r_3__126_,s_r_3__125_,s_r_3__124_,s_r_3__123_,s_r_3__122_,s_r_3__121_,
  s_r_3__120_,s_r_3__119_,s_r_3__118_,s_r_3__117_,s_r_3__116_,s_r_3__115_,s_r_3__114_,
  s_r_3__113_,s_r_3__112_,s_r_3__111_,s_r_3__110_,s_r_3__109_,s_r_3__108_,
  s_r_3__107_,s_r_3__106_,s_r_3__105_,s_r_3__104_,s_r_3__103_,s_r_3__102_,s_r_3__101_,
  s_r_3__100_,s_r_3__99_,s_r_3__98_,s_r_3__97_,s_r_3__96_,s_r_3__95_,s_r_3__94_,
  s_r_3__93_,s_r_3__92_,s_r_3__91_,s_r_3__90_,s_r_3__89_,s_r_3__88_,s_r_3__87_,s_r_3__86_,
  s_r_3__85_,s_r_3__84_,s_r_3__83_,s_r_3__82_,s_r_3__81_,s_r_3__80_,s_r_3__79_,
  s_r_3__78_,s_r_3__77_,s_r_3__76_,s_r_3__75_,s_r_3__74_,s_r_3__73_,s_r_3__72_,
  s_r_3__71_,s_r_3__70_,s_r_3__69_,s_r_3__68_,s_r_3__67_,s_r_3__66_,s_r_3__65_,
  s_r_3__64_,s_r_3__63_,s_r_3__62_,s_r_3__61_,s_r_3__60_,s_r_3__59_,s_r_3__58_,s_r_3__57_,
  s_r_3__56_,s_r_3__55_,s_r_3__54_,s_r_3__53_,s_r_3__52_,s_r_3__51_,s_r_3__50_,
  s_r_3__49_,s_r_3__48_,s_r_3__47_,s_r_3__46_,s_r_3__45_,s_r_3__44_,s_r_3__43_,
  s_r_3__42_,s_r_3__41_,s_r_3__40_,s_r_3__39_,s_r_3__38_,s_r_3__37_,s_r_3__36_,s_r_3__35_,
  s_r_3__34_,s_r_3__33_,s_r_3__32_,s_r_3__31_,s_r_3__30_,s_r_3__29_,s_r_3__28_,
  s_r_3__27_,s_r_3__26_,s_r_3__25_,s_r_3__24_,s_r_3__23_,s_r_3__22_,s_r_3__21_,
  s_r_3__20_,s_r_3__19_,s_r_3__18_,s_r_3__17_,s_r_3__16_,s_r_3__15_,s_r_3__14_,
  s_r_3__13_,s_r_3__12_,s_r_3__11_,s_r_3__10_,s_r_3__9_,s_r_3__8_,s_r_3__7_,s_r_3__6_,
  s_r_3__5_,s_r_3__4_,s_r_3__3_,s_r_3__2_,s_r_3__1_,s_r_3__0_,prod_accum_6__7_,
  prod_accum_6__6_,prod_accum_6__5_,prod_accum_6__4_,prod_accum_6__3_,prod_accum_6__2_,
  prod_accum_6__1_,prod_accum_6__0_,prod_accum_5__6_,prod_accum_5__5_,
  prod_accum_5__4_,prod_accum_5__3_,prod_accum_5__2_,prod_accum_5__1_,prod_accum_5__0_,
  prod_accum_4__5_,prod_accum_4__4_,prod_accum_4__3_,prod_accum_4__2_,prod_accum_4__1_,
  prod_accum_4__0_,prod_accum_3__4_,prod_accum_3__3_,prod_accum_3__2_,prod_accum_3__1_,
  prod_accum_3__0_,s_r_10__127_,s_r_10__126_,s_r_10__125_,s_r_10__124_,
  s_r_10__123_,s_r_10__122_,s_r_10__121_,s_r_10__120_,s_r_10__119_,s_r_10__118_,s_r_10__117_,
  s_r_10__116_,s_r_10__115_,s_r_10__114_,s_r_10__113_,s_r_10__112_,s_r_10__111_,
  s_r_10__110_,s_r_10__109_,s_r_10__108_,s_r_10__107_,s_r_10__106_,s_r_10__105_,
  s_r_10__104_,s_r_10__103_,s_r_10__102_,s_r_10__101_,s_r_10__100_,s_r_10__99_,
  s_r_10__98_,s_r_10__97_,s_r_10__96_,s_r_10__95_,s_r_10__94_,s_r_10__93_,s_r_10__92_,
  s_r_10__91_,s_r_10__90_,s_r_10__89_,s_r_10__88_,s_r_10__87_,s_r_10__86_,
  s_r_10__85_,s_r_10__84_,s_r_10__83_,s_r_10__82_,s_r_10__81_,s_r_10__80_,s_r_10__79_,
  s_r_10__78_,s_r_10__77_,s_r_10__76_,s_r_10__75_,s_r_10__74_,s_r_10__73_,s_r_10__72_,
  s_r_10__71_,s_r_10__70_,s_r_10__69_,s_r_10__68_,s_r_10__67_,s_r_10__66_,
  s_r_10__65_,s_r_10__64_,s_r_10__63_,s_r_10__62_,s_r_10__61_,s_r_10__60_,s_r_10__59_,
  s_r_10__58_,s_r_10__57_,s_r_10__56_,s_r_10__55_,s_r_10__54_,s_r_10__53_,s_r_10__52_,
  s_r_10__51_,s_r_10__50_,s_r_10__49_,s_r_10__48_,s_r_10__47_,s_r_10__46_,
  s_r_10__45_,s_r_10__44_,s_r_10__43_,s_r_10__42_,s_r_10__41_,s_r_10__40_,s_r_10__39_,
  s_r_10__38_,s_r_10__37_,s_r_10__36_,s_r_10__35_,s_r_10__34_,s_r_10__33_,s_r_10__32_,
  s_r_10__31_,s_r_10__30_,s_r_10__29_,s_r_10__28_,s_r_10__27_,s_r_10__26_,
  s_r_10__25_,s_r_10__24_,s_r_10__23_,s_r_10__22_,s_r_10__21_,s_r_10__20_,s_r_10__19_,
  s_r_10__18_,s_r_10__17_,s_r_10__16_,s_r_10__15_,s_r_10__14_,s_r_10__13_,s_r_10__12_,
  s_r_10__11_,s_r_10__10_,s_r_10__9_,s_r_10__8_,s_r_10__7_,s_r_10__6_,s_r_10__5_,
  s_r_10__4_,s_r_10__3_,s_r_10__2_,s_r_10__1_,s_r_10__0_,s_r_9__127_,s_r_9__126_,
  s_r_9__125_,s_r_9__124_,s_r_9__123_,s_r_9__122_,s_r_9__121_,s_r_9__120_,s_r_9__119_,
  s_r_9__118_,s_r_9__117_,s_r_9__116_,s_r_9__115_,s_r_9__114_,s_r_9__113_,
  s_r_9__112_,s_r_9__111_,s_r_9__110_,s_r_9__109_,s_r_9__108_,s_r_9__107_,s_r_9__106_,
  s_r_9__105_,s_r_9__104_,s_r_9__103_,s_r_9__102_,s_r_9__101_,s_r_9__100_,s_r_9__99_,
  s_r_9__98_,s_r_9__97_,s_r_9__96_,s_r_9__95_,s_r_9__94_,s_r_9__93_,s_r_9__92_,
  s_r_9__91_,s_r_9__90_,s_r_9__89_,s_r_9__88_,s_r_9__87_,s_r_9__86_,s_r_9__85_,
  s_r_9__84_,s_r_9__83_,s_r_9__82_,s_r_9__81_,s_r_9__80_,s_r_9__79_,s_r_9__78_,s_r_9__77_,
  s_r_9__76_,s_r_9__75_,s_r_9__74_,s_r_9__73_,s_r_9__72_,s_r_9__71_,s_r_9__70_,
  s_r_9__69_,s_r_9__68_,s_r_9__67_,s_r_9__66_,s_r_9__65_,s_r_9__64_,s_r_9__63_,
  s_r_9__62_,s_r_9__61_,s_r_9__60_,s_r_9__59_,s_r_9__58_,s_r_9__57_,s_r_9__56_,
  s_r_9__55_,s_r_9__54_,s_r_9__53_,s_r_9__52_,s_r_9__51_,s_r_9__50_,s_r_9__49_,s_r_9__48_,
  s_r_9__47_,s_r_9__46_,s_r_9__45_,s_r_9__44_,s_r_9__43_,s_r_9__42_,s_r_9__41_,
  s_r_9__40_,s_r_9__39_,s_r_9__38_,s_r_9__37_,s_r_9__36_,s_r_9__35_,s_r_9__34_,
  s_r_9__33_,s_r_9__32_,s_r_9__31_,s_r_9__30_,s_r_9__29_,s_r_9__28_,s_r_9__27_,
  s_r_9__26_,s_r_9__25_,s_r_9__24_,s_r_9__23_,s_r_9__22_,s_r_9__21_,s_r_9__20_,s_r_9__19_,
  s_r_9__18_,s_r_9__17_,s_r_9__16_,s_r_9__15_,s_r_9__14_,s_r_9__13_,s_r_9__12_,
  s_r_9__11_,s_r_9__10_,s_r_9__9_,s_r_9__8_,s_r_9__7_,s_r_9__6_,s_r_9__5_,s_r_9__4_,
  s_r_9__3_,s_r_9__2_,s_r_9__1_,s_r_9__0_,s_r_8__127_,s_r_8__126_,s_r_8__125_,
  s_r_8__124_,s_r_8__123_,s_r_8__122_,s_r_8__121_,s_r_8__120_,s_r_8__119_,s_r_8__118_,
  s_r_8__117_,s_r_8__116_,s_r_8__115_,s_r_8__114_,s_r_8__113_,s_r_8__112_,
  s_r_8__111_,s_r_8__110_,s_r_8__109_,s_r_8__108_,s_r_8__107_,s_r_8__106_,s_r_8__105_,
  s_r_8__104_,s_r_8__103_,s_r_8__102_,s_r_8__101_,s_r_8__100_,s_r_8__99_,s_r_8__98_,
  s_r_8__97_,s_r_8__96_,s_r_8__95_,s_r_8__94_,s_r_8__93_,s_r_8__92_,s_r_8__91_,
  s_r_8__90_,s_r_8__89_,s_r_8__88_,s_r_8__87_,s_r_8__86_,s_r_8__85_,s_r_8__84_,s_r_8__83_,
  s_r_8__82_,s_r_8__81_,s_r_8__80_,s_r_8__79_,s_r_8__78_,s_r_8__77_,s_r_8__76_,
  s_r_8__75_,s_r_8__74_,s_r_8__73_,s_r_8__72_,s_r_8__71_,s_r_8__70_,s_r_8__69_,
  s_r_8__68_,s_r_8__67_,s_r_8__66_,s_r_8__65_,s_r_8__64_,s_r_8__63_,s_r_8__62_,
  s_r_8__61_,s_r_8__60_,s_r_8__59_,s_r_8__58_,s_r_8__57_,s_r_8__56_,s_r_8__55_,s_r_8__54_,
  s_r_8__53_,s_r_8__52_,s_r_8__51_,s_r_8__50_,s_r_8__49_,s_r_8__48_,s_r_8__47_,
  s_r_8__46_,s_r_8__45_,s_r_8__44_,s_r_8__43_,s_r_8__42_,s_r_8__41_,s_r_8__40_,
  s_r_8__39_,s_r_8__38_,s_r_8__37_,s_r_8__36_,s_r_8__35_,s_r_8__34_,s_r_8__33_,
  s_r_8__32_,s_r_8__31_,s_r_8__30_,s_r_8__29_,s_r_8__28_,s_r_8__27_,s_r_8__26_,s_r_8__25_,
  s_r_8__24_,s_r_8__23_,s_r_8__22_,s_r_8__21_,s_r_8__20_,s_r_8__19_,s_r_8__18_,
  s_r_8__17_,s_r_8__16_,s_r_8__15_,s_r_8__14_,s_r_8__13_,s_r_8__12_,s_r_8__11_,
  s_r_8__10_,s_r_8__9_,s_r_8__8_,s_r_8__7_,s_r_8__6_,s_r_8__5_,s_r_8__4_,s_r_8__3_,
  s_r_8__2_,s_r_8__1_,s_r_8__0_,s_r_7__127_,s_r_7__126_,s_r_7__125_,s_r_7__124_,
  s_r_7__123_,s_r_7__122_,s_r_7__121_,s_r_7__120_,s_r_7__119_,s_r_7__118_,s_r_7__117_,
  s_r_7__116_,s_r_7__115_,s_r_7__114_,s_r_7__113_,s_r_7__112_,s_r_7__111_,s_r_7__110_,
  s_r_7__109_,s_r_7__108_,s_r_7__107_,s_r_7__106_,s_r_7__105_,s_r_7__104_,
  s_r_7__103_,s_r_7__102_,s_r_7__101_,s_r_7__100_,s_r_7__99_,s_r_7__98_,s_r_7__97_,
  s_r_7__96_,s_r_7__95_,s_r_7__94_,s_r_7__93_,s_r_7__92_,s_r_7__91_,s_r_7__90_,s_r_7__89_,
  s_r_7__88_,s_r_7__87_,s_r_7__86_,s_r_7__85_,s_r_7__84_,s_r_7__83_,s_r_7__82_,
  s_r_7__81_,s_r_7__80_,s_r_7__79_,s_r_7__78_,s_r_7__77_,s_r_7__76_,s_r_7__75_,
  s_r_7__74_,s_r_7__73_,s_r_7__72_,s_r_7__71_,s_r_7__70_,s_r_7__69_,s_r_7__68_,
  s_r_7__67_,s_r_7__66_,s_r_7__65_,s_r_7__64_,s_r_7__63_,s_r_7__62_,s_r_7__61_,s_r_7__60_,
  s_r_7__59_,s_r_7__58_,s_r_7__57_,s_r_7__56_,s_r_7__55_,s_r_7__54_,s_r_7__53_,
  s_r_7__52_,s_r_7__51_,s_r_7__50_,s_r_7__49_,s_r_7__48_,s_r_7__47_,s_r_7__46_,
  s_r_7__45_,s_r_7__44_,s_r_7__43_,s_r_7__42_,s_r_7__41_,s_r_7__40_,s_r_7__39_,
  s_r_7__38_,s_r_7__37_,s_r_7__36_,s_r_7__35_,s_r_7__34_,s_r_7__33_,s_r_7__32_,s_r_7__31_,
  s_r_7__30_,s_r_7__29_,s_r_7__28_,s_r_7__27_,s_r_7__26_,s_r_7__25_,s_r_7__24_,
  s_r_7__23_,s_r_7__22_,s_r_7__21_,s_r_7__20_,s_r_7__19_,s_r_7__18_,s_r_7__17_,
  s_r_7__16_,s_r_7__15_,s_r_7__14_,s_r_7__13_,s_r_7__12_,s_r_7__11_,s_r_7__10_,s_r_7__9_,
  s_r_7__8_,s_r_7__7_,s_r_7__6_,s_r_7__5_,s_r_7__4_,s_r_7__3_,s_r_7__2_,s_r_7__1_,
  s_r_7__0_,prod_accum_10__11_,prod_accum_10__10_,prod_accum_10__9_,
  prod_accum_10__8_,prod_accum_10__7_,prod_accum_10__6_,prod_accum_10__5_,prod_accum_10__4_,
  prod_accum_10__3_,prod_accum_10__2_,prod_accum_10__1_,prod_accum_10__0_,
  prod_accum_9__10_,prod_accum_9__9_,prod_accum_9__8_,prod_accum_9__7_,prod_accum_9__6_,
  prod_accum_9__5_,prod_accum_9__4_,prod_accum_9__3_,prod_accum_9__2_,prod_accum_9__1_,
  prod_accum_9__0_,prod_accum_8__9_,prod_accum_8__8_,prod_accum_8__7_,
  prod_accum_8__6_,prod_accum_8__5_,prod_accum_8__4_,prod_accum_8__3_,prod_accum_8__2_,
  prod_accum_8__1_,prod_accum_8__0_,prod_accum_7__8_,prod_accum_7__7_,prod_accum_7__6_,
  prod_accum_7__5_,prod_accum_7__4_,prod_accum_7__3_,prod_accum_7__2_,
  prod_accum_7__1_,prod_accum_7__0_,s_r_14__127_,s_r_14__126_,s_r_14__125_,s_r_14__124_,
  s_r_14__123_,s_r_14__122_,s_r_14__121_,s_r_14__120_,s_r_14__119_,s_r_14__118_,
  s_r_14__117_,s_r_14__116_,s_r_14__115_,s_r_14__114_,s_r_14__113_,s_r_14__112_,s_r_14__111_,
  s_r_14__110_,s_r_14__109_,s_r_14__108_,s_r_14__107_,s_r_14__106_,s_r_14__105_,
  s_r_14__104_,s_r_14__103_,s_r_14__102_,s_r_14__101_,s_r_14__100_,s_r_14__99_,
  s_r_14__98_,s_r_14__97_,s_r_14__96_,s_r_14__95_,s_r_14__94_,s_r_14__93_,s_r_14__92_,
  s_r_14__91_,s_r_14__90_,s_r_14__89_,s_r_14__88_,s_r_14__87_,s_r_14__86_,
  s_r_14__85_,s_r_14__84_,s_r_14__83_,s_r_14__82_,s_r_14__81_,s_r_14__80_,s_r_14__79_,
  s_r_14__78_,s_r_14__77_,s_r_14__76_,s_r_14__75_,s_r_14__74_,s_r_14__73_,s_r_14__72_,
  s_r_14__71_,s_r_14__70_,s_r_14__69_,s_r_14__68_,s_r_14__67_,s_r_14__66_,
  s_r_14__65_,s_r_14__64_,s_r_14__63_,s_r_14__62_,s_r_14__61_,s_r_14__60_,s_r_14__59_,
  s_r_14__58_,s_r_14__57_,s_r_14__56_,s_r_14__55_,s_r_14__54_,s_r_14__53_,s_r_14__52_,
  s_r_14__51_,s_r_14__50_,s_r_14__49_,s_r_14__48_,s_r_14__47_,s_r_14__46_,
  s_r_14__45_,s_r_14__44_,s_r_14__43_,s_r_14__42_,s_r_14__41_,s_r_14__40_,s_r_14__39_,
  s_r_14__38_,s_r_14__37_,s_r_14__36_,s_r_14__35_,s_r_14__34_,s_r_14__33_,s_r_14__32_,
  s_r_14__31_,s_r_14__30_,s_r_14__29_,s_r_14__28_,s_r_14__27_,s_r_14__26_,
  s_r_14__25_,s_r_14__24_,s_r_14__23_,s_r_14__22_,s_r_14__21_,s_r_14__20_,s_r_14__19_,
  s_r_14__18_,s_r_14__17_,s_r_14__16_,s_r_14__15_,s_r_14__14_,s_r_14__13_,s_r_14__12_,
  s_r_14__11_,s_r_14__10_,s_r_14__9_,s_r_14__8_,s_r_14__7_,s_r_14__6_,s_r_14__5_,
  s_r_14__4_,s_r_14__3_,s_r_14__2_,s_r_14__1_,s_r_14__0_,s_r_13__127_,s_r_13__126_,
  s_r_13__125_,s_r_13__124_,s_r_13__123_,s_r_13__122_,s_r_13__121_,s_r_13__120_,
  s_r_13__119_,s_r_13__118_,s_r_13__117_,s_r_13__116_,s_r_13__115_,s_r_13__114_,
  s_r_13__113_,s_r_13__112_,s_r_13__111_,s_r_13__110_,s_r_13__109_,s_r_13__108_,
  s_r_13__107_,s_r_13__106_,s_r_13__105_,s_r_13__104_,s_r_13__103_,s_r_13__102_,
  s_r_13__101_,s_r_13__100_,s_r_13__99_,s_r_13__98_,s_r_13__97_,s_r_13__96_,s_r_13__95_,
  s_r_13__94_,s_r_13__93_,s_r_13__92_,s_r_13__91_,s_r_13__90_,s_r_13__89_,s_r_13__88_,
  s_r_13__87_,s_r_13__86_,s_r_13__85_,s_r_13__84_,s_r_13__83_,s_r_13__82_,
  s_r_13__81_,s_r_13__80_,s_r_13__79_,s_r_13__78_,s_r_13__77_,s_r_13__76_,s_r_13__75_,
  s_r_13__74_,s_r_13__73_,s_r_13__72_,s_r_13__71_,s_r_13__70_,s_r_13__69_,s_r_13__68_,
  s_r_13__67_,s_r_13__66_,s_r_13__65_,s_r_13__64_,s_r_13__63_,s_r_13__62_,
  s_r_13__61_,s_r_13__60_,s_r_13__59_,s_r_13__58_,s_r_13__57_,s_r_13__56_,s_r_13__55_,
  s_r_13__54_,s_r_13__53_,s_r_13__52_,s_r_13__51_,s_r_13__50_,s_r_13__49_,s_r_13__48_,
  s_r_13__47_,s_r_13__46_,s_r_13__45_,s_r_13__44_,s_r_13__43_,s_r_13__42_,
  s_r_13__41_,s_r_13__40_,s_r_13__39_,s_r_13__38_,s_r_13__37_,s_r_13__36_,s_r_13__35_,
  s_r_13__34_,s_r_13__33_,s_r_13__32_,s_r_13__31_,s_r_13__30_,s_r_13__29_,s_r_13__28_,
  s_r_13__27_,s_r_13__26_,s_r_13__25_,s_r_13__24_,s_r_13__23_,s_r_13__22_,
  s_r_13__21_,s_r_13__20_,s_r_13__19_,s_r_13__18_,s_r_13__17_,s_r_13__16_,s_r_13__15_,
  s_r_13__14_,s_r_13__13_,s_r_13__12_,s_r_13__11_,s_r_13__10_,s_r_13__9_,s_r_13__8_,
  s_r_13__7_,s_r_13__6_,s_r_13__5_,s_r_13__4_,s_r_13__3_,s_r_13__2_,s_r_13__1_,
  s_r_13__0_,s_r_12__127_,s_r_12__126_,s_r_12__125_,s_r_12__124_,s_r_12__123_,
  s_r_12__122_,s_r_12__121_,s_r_12__120_,s_r_12__119_,s_r_12__118_,s_r_12__117_,
  s_r_12__116_,s_r_12__115_,s_r_12__114_,s_r_12__113_,s_r_12__112_,s_r_12__111_,s_r_12__110_,
  s_r_12__109_,s_r_12__108_,s_r_12__107_,s_r_12__106_,s_r_12__105_,s_r_12__104_,
  s_r_12__103_,s_r_12__102_,s_r_12__101_,s_r_12__100_,s_r_12__99_,s_r_12__98_,
  s_r_12__97_,s_r_12__96_,s_r_12__95_,s_r_12__94_,s_r_12__93_,s_r_12__92_,s_r_12__91_,
  s_r_12__90_,s_r_12__89_,s_r_12__88_,s_r_12__87_,s_r_12__86_,s_r_12__85_,
  s_r_12__84_,s_r_12__83_,s_r_12__82_,s_r_12__81_,s_r_12__80_,s_r_12__79_,s_r_12__78_,
  s_r_12__77_,s_r_12__76_,s_r_12__75_,s_r_12__74_,s_r_12__73_,s_r_12__72_,s_r_12__71_,
  s_r_12__70_,s_r_12__69_,s_r_12__68_,s_r_12__67_,s_r_12__66_,s_r_12__65_,
  s_r_12__64_,s_r_12__63_,s_r_12__62_,s_r_12__61_,s_r_12__60_,s_r_12__59_,s_r_12__58_,
  s_r_12__57_,s_r_12__56_,s_r_12__55_,s_r_12__54_,s_r_12__53_,s_r_12__52_,s_r_12__51_,
  s_r_12__50_,s_r_12__49_,s_r_12__48_,s_r_12__47_,s_r_12__46_,s_r_12__45_,
  s_r_12__44_,s_r_12__43_,s_r_12__42_,s_r_12__41_,s_r_12__40_,s_r_12__39_,s_r_12__38_,
  s_r_12__37_,s_r_12__36_,s_r_12__35_,s_r_12__34_,s_r_12__33_,s_r_12__32_,s_r_12__31_,
  s_r_12__30_,s_r_12__29_,s_r_12__28_,s_r_12__27_,s_r_12__26_,s_r_12__25_,
  s_r_12__24_,s_r_12__23_,s_r_12__22_,s_r_12__21_,s_r_12__20_,s_r_12__19_,s_r_12__18_,
  s_r_12__17_,s_r_12__16_,s_r_12__15_,s_r_12__14_,s_r_12__13_,s_r_12__12_,s_r_12__11_,
  s_r_12__10_,s_r_12__9_,s_r_12__8_,s_r_12__7_,s_r_12__6_,s_r_12__5_,s_r_12__4_,
  s_r_12__3_,s_r_12__2_,s_r_12__1_,s_r_12__0_,s_r_11__127_,s_r_11__126_,s_r_11__125_,
  s_r_11__124_,s_r_11__123_,s_r_11__122_,s_r_11__121_,s_r_11__120_,s_r_11__119_,
  s_r_11__118_,s_r_11__117_,s_r_11__116_,s_r_11__115_,s_r_11__114_,s_r_11__113_,
  s_r_11__112_,s_r_11__111_,s_r_11__110_,s_r_11__109_,s_r_11__108_,s_r_11__107_,
  s_r_11__106_,s_r_11__105_,s_r_11__104_,s_r_11__103_,s_r_11__102_,s_r_11__101_,
  s_r_11__100_,s_r_11__99_,s_r_11__98_,s_r_11__97_,s_r_11__96_,s_r_11__95_,s_r_11__94_,
  s_r_11__93_,s_r_11__92_,s_r_11__91_,s_r_11__90_,s_r_11__89_,s_r_11__88_,s_r_11__87_,
  s_r_11__86_,s_r_11__85_,s_r_11__84_,s_r_11__83_,s_r_11__82_,s_r_11__81_,
  s_r_11__80_,s_r_11__79_,s_r_11__78_,s_r_11__77_,s_r_11__76_,s_r_11__75_,s_r_11__74_,
  s_r_11__73_,s_r_11__72_,s_r_11__71_,s_r_11__70_,s_r_11__69_,s_r_11__68_,s_r_11__67_,
  s_r_11__66_,s_r_11__65_,s_r_11__64_,s_r_11__63_,s_r_11__62_,s_r_11__61_,
  s_r_11__60_,s_r_11__59_,s_r_11__58_,s_r_11__57_,s_r_11__56_,s_r_11__55_,s_r_11__54_,
  s_r_11__53_,s_r_11__52_,s_r_11__51_,s_r_11__50_,s_r_11__49_,s_r_11__48_,s_r_11__47_,
  s_r_11__46_,s_r_11__45_,s_r_11__44_,s_r_11__43_,s_r_11__42_,s_r_11__41_,
  s_r_11__40_,s_r_11__39_,s_r_11__38_,s_r_11__37_,s_r_11__36_,s_r_11__35_,s_r_11__34_,
  s_r_11__33_,s_r_11__32_,s_r_11__31_,s_r_11__30_,s_r_11__29_,s_r_11__28_,s_r_11__27_,
  s_r_11__26_,s_r_11__25_,s_r_11__24_,s_r_11__23_,s_r_11__22_,s_r_11__21_,
  s_r_11__20_,s_r_11__19_,s_r_11__18_,s_r_11__17_,s_r_11__16_,s_r_11__15_,s_r_11__14_,
  s_r_11__13_,s_r_11__12_,s_r_11__11_,s_r_11__10_,s_r_11__9_,s_r_11__8_,s_r_11__7_,
  s_r_11__6_,s_r_11__5_,s_r_11__4_,s_r_11__3_,s_r_11__2_,s_r_11__1_,s_r_11__0_,
  prod_accum_14__15_,prod_accum_14__14_,prod_accum_14__13_,prod_accum_14__12_,
  prod_accum_14__11_,prod_accum_14__10_,prod_accum_14__9_,prod_accum_14__8_,
  prod_accum_14__7_,prod_accum_14__6_,prod_accum_14__5_,prod_accum_14__4_,prod_accum_14__3_,
  prod_accum_14__2_,prod_accum_14__1_,prod_accum_14__0_,prod_accum_13__14_,
  prod_accum_13__13_,prod_accum_13__12_,prod_accum_13__11_,prod_accum_13__10_,
  prod_accum_13__9_,prod_accum_13__8_,prod_accum_13__7_,prod_accum_13__6_,prod_accum_13__5_,
  prod_accum_13__4_,prod_accum_13__3_,prod_accum_13__2_,prod_accum_13__1_,
  prod_accum_13__0_,prod_accum_12__13_,prod_accum_12__12_,prod_accum_12__11_,prod_accum_12__10_,
  prod_accum_12__9_,prod_accum_12__8_,prod_accum_12__7_,prod_accum_12__6_,
  prod_accum_12__5_,prod_accum_12__4_,prod_accum_12__3_,prod_accum_12__2_,
  prod_accum_12__1_,prod_accum_12__0_,prod_accum_11__12_,prod_accum_11__11_,prod_accum_11__10_,
  prod_accum_11__9_,prod_accum_11__8_,prod_accum_11__7_,prod_accum_11__6_,
  prod_accum_11__5_,prod_accum_11__4_,prod_accum_11__3_,prod_accum_11__2_,prod_accum_11__1_,
  prod_accum_11__0_,s_r_18__127_,s_r_18__126_,s_r_18__125_,s_r_18__124_,
  s_r_18__123_,s_r_18__122_,s_r_18__121_,s_r_18__120_,s_r_18__119_,s_r_18__118_,s_r_18__117_,
  s_r_18__116_,s_r_18__115_,s_r_18__114_,s_r_18__113_,s_r_18__112_,s_r_18__111_,
  s_r_18__110_,s_r_18__109_,s_r_18__108_,s_r_18__107_,s_r_18__106_,s_r_18__105_,
  s_r_18__104_,s_r_18__103_,s_r_18__102_,s_r_18__101_,s_r_18__100_,s_r_18__99_,
  s_r_18__98_,s_r_18__97_,s_r_18__96_,s_r_18__95_,s_r_18__94_,s_r_18__93_,s_r_18__92_,
  s_r_18__91_,s_r_18__90_,s_r_18__89_,s_r_18__88_,s_r_18__87_,s_r_18__86_,s_r_18__85_,
  s_r_18__84_,s_r_18__83_,s_r_18__82_,s_r_18__81_,s_r_18__80_,s_r_18__79_,
  s_r_18__78_,s_r_18__77_,s_r_18__76_,s_r_18__75_,s_r_18__74_,s_r_18__73_,s_r_18__72_,
  s_r_18__71_,s_r_18__70_,s_r_18__69_,s_r_18__68_,s_r_18__67_,s_r_18__66_,s_r_18__65_,
  s_r_18__64_,s_r_18__63_,s_r_18__62_,s_r_18__61_,s_r_18__60_,s_r_18__59_,
  s_r_18__58_,s_r_18__57_,s_r_18__56_,s_r_18__55_,s_r_18__54_,s_r_18__53_,s_r_18__52_,
  s_r_18__51_,s_r_18__50_,s_r_18__49_,s_r_18__48_,s_r_18__47_,s_r_18__46_,s_r_18__45_,
  s_r_18__44_,s_r_18__43_,s_r_18__42_,s_r_18__41_,s_r_18__40_,s_r_18__39_,
  s_r_18__38_,s_r_18__37_,s_r_18__36_,s_r_18__35_,s_r_18__34_,s_r_18__33_,s_r_18__32_,
  s_r_18__31_,s_r_18__30_,s_r_18__29_,s_r_18__28_,s_r_18__27_,s_r_18__26_,s_r_18__25_,
  s_r_18__24_,s_r_18__23_,s_r_18__22_,s_r_18__21_,s_r_18__20_,s_r_18__19_,
  s_r_18__18_,s_r_18__17_,s_r_18__16_,s_r_18__15_,s_r_18__14_,s_r_18__13_,s_r_18__12_,
  s_r_18__11_,s_r_18__10_,s_r_18__9_,s_r_18__8_,s_r_18__7_,s_r_18__6_,s_r_18__5_,
  s_r_18__4_,s_r_18__3_,s_r_18__2_,s_r_18__1_,s_r_18__0_,s_r_17__127_,s_r_17__126_,
  s_r_17__125_,s_r_17__124_,s_r_17__123_,s_r_17__122_,s_r_17__121_,s_r_17__120_,
  s_r_17__119_,s_r_17__118_,s_r_17__117_,s_r_17__116_,s_r_17__115_,s_r_17__114_,
  s_r_17__113_,s_r_17__112_,s_r_17__111_,s_r_17__110_,s_r_17__109_,s_r_17__108_,
  s_r_17__107_,s_r_17__106_,s_r_17__105_,s_r_17__104_,s_r_17__103_,s_r_17__102_,
  s_r_17__101_,s_r_17__100_,s_r_17__99_,s_r_17__98_,s_r_17__97_,s_r_17__96_,s_r_17__95_,
  s_r_17__94_,s_r_17__93_,s_r_17__92_,s_r_17__91_,s_r_17__90_,s_r_17__89_,s_r_17__88_,
  s_r_17__87_,s_r_17__86_,s_r_17__85_,s_r_17__84_,s_r_17__83_,s_r_17__82_,
  s_r_17__81_,s_r_17__80_,s_r_17__79_,s_r_17__78_,s_r_17__77_,s_r_17__76_,s_r_17__75_,
  s_r_17__74_,s_r_17__73_,s_r_17__72_,s_r_17__71_,s_r_17__70_,s_r_17__69_,s_r_17__68_,
  s_r_17__67_,s_r_17__66_,s_r_17__65_,s_r_17__64_,s_r_17__63_,s_r_17__62_,
  s_r_17__61_,s_r_17__60_,s_r_17__59_,s_r_17__58_,s_r_17__57_,s_r_17__56_,s_r_17__55_,
  s_r_17__54_,s_r_17__53_,s_r_17__52_,s_r_17__51_,s_r_17__50_,s_r_17__49_,s_r_17__48_,
  s_r_17__47_,s_r_17__46_,s_r_17__45_,s_r_17__44_,s_r_17__43_,s_r_17__42_,
  s_r_17__41_,s_r_17__40_,s_r_17__39_,s_r_17__38_,s_r_17__37_,s_r_17__36_,s_r_17__35_,
  s_r_17__34_,s_r_17__33_,s_r_17__32_,s_r_17__31_,s_r_17__30_,s_r_17__29_,s_r_17__28_,
  s_r_17__27_,s_r_17__26_,s_r_17__25_,s_r_17__24_,s_r_17__23_,s_r_17__22_,
  s_r_17__21_,s_r_17__20_,s_r_17__19_,s_r_17__18_,s_r_17__17_,s_r_17__16_,s_r_17__15_,
  s_r_17__14_,s_r_17__13_,s_r_17__12_,s_r_17__11_,s_r_17__10_,s_r_17__9_,s_r_17__8_,
  s_r_17__7_,s_r_17__6_,s_r_17__5_,s_r_17__4_,s_r_17__3_,s_r_17__2_,s_r_17__1_,
  s_r_17__0_,s_r_16__127_,s_r_16__126_,s_r_16__125_,s_r_16__124_,s_r_16__123_,
  s_r_16__122_,s_r_16__121_,s_r_16__120_,s_r_16__119_,s_r_16__118_,s_r_16__117_,s_r_16__116_,
  s_r_16__115_,s_r_16__114_,s_r_16__113_,s_r_16__112_,s_r_16__111_,s_r_16__110_,
  s_r_16__109_,s_r_16__108_,s_r_16__107_,s_r_16__106_,s_r_16__105_,s_r_16__104_,
  s_r_16__103_,s_r_16__102_,s_r_16__101_,s_r_16__100_,s_r_16__99_,s_r_16__98_,
  s_r_16__97_,s_r_16__96_,s_r_16__95_,s_r_16__94_,s_r_16__93_,s_r_16__92_,s_r_16__91_,
  s_r_16__90_,s_r_16__89_,s_r_16__88_,s_r_16__87_,s_r_16__86_,s_r_16__85_,s_r_16__84_,
  s_r_16__83_,s_r_16__82_,s_r_16__81_,s_r_16__80_,s_r_16__79_,s_r_16__78_,
  s_r_16__77_,s_r_16__76_,s_r_16__75_,s_r_16__74_,s_r_16__73_,s_r_16__72_,s_r_16__71_,
  s_r_16__70_,s_r_16__69_,s_r_16__68_,s_r_16__67_,s_r_16__66_,s_r_16__65_,s_r_16__64_,
  s_r_16__63_,s_r_16__62_,s_r_16__61_,s_r_16__60_,s_r_16__59_,s_r_16__58_,
  s_r_16__57_,s_r_16__56_,s_r_16__55_,s_r_16__54_,s_r_16__53_,s_r_16__52_,s_r_16__51_,
  s_r_16__50_,s_r_16__49_,s_r_16__48_,s_r_16__47_,s_r_16__46_,s_r_16__45_,s_r_16__44_,
  s_r_16__43_,s_r_16__42_,s_r_16__41_,s_r_16__40_,s_r_16__39_,s_r_16__38_,
  s_r_16__37_,s_r_16__36_,s_r_16__35_,s_r_16__34_,s_r_16__33_,s_r_16__32_,s_r_16__31_,
  s_r_16__30_,s_r_16__29_,s_r_16__28_,s_r_16__27_,s_r_16__26_,s_r_16__25_,s_r_16__24_,
  s_r_16__23_,s_r_16__22_,s_r_16__21_,s_r_16__20_,s_r_16__19_,s_r_16__18_,
  s_r_16__17_,s_r_16__16_,s_r_16__15_,s_r_16__14_,s_r_16__13_,s_r_16__12_,s_r_16__11_,
  s_r_16__10_,s_r_16__9_,s_r_16__8_,s_r_16__7_,s_r_16__6_,s_r_16__5_,s_r_16__4_,
  s_r_16__3_,s_r_16__2_,s_r_16__1_,s_r_16__0_,s_r_15__127_,s_r_15__126_,s_r_15__125_,
  s_r_15__124_,s_r_15__123_,s_r_15__122_,s_r_15__121_,s_r_15__120_,s_r_15__119_,
  s_r_15__118_,s_r_15__117_,s_r_15__116_,s_r_15__115_,s_r_15__114_,s_r_15__113_,
  s_r_15__112_,s_r_15__111_,s_r_15__110_,s_r_15__109_,s_r_15__108_,s_r_15__107_,
  s_r_15__106_,s_r_15__105_,s_r_15__104_,s_r_15__103_,s_r_15__102_,s_r_15__101_,
  s_r_15__100_,s_r_15__99_,s_r_15__98_,s_r_15__97_,s_r_15__96_,s_r_15__95_,s_r_15__94_,
  s_r_15__93_,s_r_15__92_,s_r_15__91_,s_r_15__90_,s_r_15__89_,s_r_15__88_,s_r_15__87_,
  s_r_15__86_,s_r_15__85_,s_r_15__84_,s_r_15__83_,s_r_15__82_,s_r_15__81_,
  s_r_15__80_,s_r_15__79_,s_r_15__78_,s_r_15__77_,s_r_15__76_,s_r_15__75_,s_r_15__74_,
  s_r_15__73_,s_r_15__72_,s_r_15__71_,s_r_15__70_,s_r_15__69_,s_r_15__68_,s_r_15__67_,
  s_r_15__66_,s_r_15__65_,s_r_15__64_,s_r_15__63_,s_r_15__62_,s_r_15__61_,
  s_r_15__60_,s_r_15__59_,s_r_15__58_,s_r_15__57_,s_r_15__56_,s_r_15__55_,s_r_15__54_,
  s_r_15__53_,s_r_15__52_,s_r_15__51_,s_r_15__50_,s_r_15__49_,s_r_15__48_,s_r_15__47_,
  s_r_15__46_,s_r_15__45_,s_r_15__44_,s_r_15__43_,s_r_15__42_,s_r_15__41_,
  s_r_15__40_,s_r_15__39_,s_r_15__38_,s_r_15__37_,s_r_15__36_,s_r_15__35_,s_r_15__34_,
  s_r_15__33_,s_r_15__32_,s_r_15__31_,s_r_15__30_,s_r_15__29_,s_r_15__28_,s_r_15__27_,
  s_r_15__26_,s_r_15__25_,s_r_15__24_,s_r_15__23_,s_r_15__22_,s_r_15__21_,
  s_r_15__20_,s_r_15__19_,s_r_15__18_,s_r_15__17_,s_r_15__16_,s_r_15__15_,s_r_15__14_,
  s_r_15__13_,s_r_15__12_,s_r_15__11_,s_r_15__10_,s_r_15__9_,s_r_15__8_,s_r_15__7_,
  s_r_15__6_,s_r_15__5_,s_r_15__4_,s_r_15__3_,s_r_15__2_,s_r_15__1_,s_r_15__0_,
  prod_accum_18__19_,prod_accum_18__18_,prod_accum_18__17_,prod_accum_18__16_,
  prod_accum_18__15_,prod_accum_18__14_,prod_accum_18__13_,prod_accum_18__12_,
  prod_accum_18__11_,prod_accum_18__10_,prod_accum_18__9_,prod_accum_18__8_,prod_accum_18__7_,
  prod_accum_18__6_,prod_accum_18__5_,prod_accum_18__4_,prod_accum_18__3_,
  prod_accum_18__2_,prod_accum_18__1_,prod_accum_18__0_,prod_accum_17__18_,prod_accum_17__17_,
  prod_accum_17__16_,prod_accum_17__15_,prod_accum_17__14_,prod_accum_17__13_,
  prod_accum_17__12_,prod_accum_17__11_,prod_accum_17__10_,prod_accum_17__9_,
  prod_accum_17__8_,prod_accum_17__7_,prod_accum_17__6_,prod_accum_17__5_,
  prod_accum_17__4_,prod_accum_17__3_,prod_accum_17__2_,prod_accum_17__1_,prod_accum_17__0_,
  prod_accum_16__17_,prod_accum_16__16_,prod_accum_16__15_,prod_accum_16__14_,
  prod_accum_16__13_,prod_accum_16__12_,prod_accum_16__11_,prod_accum_16__10_,
  prod_accum_16__9_,prod_accum_16__8_,prod_accum_16__7_,prod_accum_16__6_,prod_accum_16__5_,
  prod_accum_16__4_,prod_accum_16__3_,prod_accum_16__2_,prod_accum_16__1_,
  prod_accum_16__0_,prod_accum_15__16_,prod_accum_15__15_,prod_accum_15__14_,
  prod_accum_15__13_,prod_accum_15__12_,prod_accum_15__11_,prod_accum_15__10_,prod_accum_15__9_,
  prod_accum_15__8_,prod_accum_15__7_,prod_accum_15__6_,prod_accum_15__5_,
  prod_accum_15__4_,prod_accum_15__3_,prod_accum_15__2_,prod_accum_15__1_,prod_accum_15__0_,
  s_r_22__127_,s_r_22__126_,s_r_22__125_,s_r_22__124_,s_r_22__123_,s_r_22__122_,
  s_r_22__121_,s_r_22__120_,s_r_22__119_,s_r_22__118_,s_r_22__117_,s_r_22__116_,
  s_r_22__115_,s_r_22__114_,s_r_22__113_,s_r_22__112_,s_r_22__111_,s_r_22__110_,
  s_r_22__109_,s_r_22__108_,s_r_22__107_,s_r_22__106_,s_r_22__105_,s_r_22__104_,
  s_r_22__103_,s_r_22__102_,s_r_22__101_,s_r_22__100_,s_r_22__99_,s_r_22__98_,s_r_22__97_,
  s_r_22__96_,s_r_22__95_,s_r_22__94_,s_r_22__93_,s_r_22__92_,s_r_22__91_,
  s_r_22__90_,s_r_22__89_,s_r_22__88_,s_r_22__87_,s_r_22__86_,s_r_22__85_,s_r_22__84_,
  s_r_22__83_,s_r_22__82_,s_r_22__81_,s_r_22__80_,s_r_22__79_,s_r_22__78_,s_r_22__77_,
  s_r_22__76_,s_r_22__75_,s_r_22__74_,s_r_22__73_,s_r_22__72_,s_r_22__71_,
  s_r_22__70_,s_r_22__69_,s_r_22__68_,s_r_22__67_,s_r_22__66_,s_r_22__65_,s_r_22__64_,
  s_r_22__63_,s_r_22__62_,s_r_22__61_,s_r_22__60_,s_r_22__59_,s_r_22__58_,s_r_22__57_,
  s_r_22__56_,s_r_22__55_,s_r_22__54_,s_r_22__53_,s_r_22__52_,s_r_22__51_,
  s_r_22__50_,s_r_22__49_,s_r_22__48_,s_r_22__47_,s_r_22__46_,s_r_22__45_,s_r_22__44_,
  s_r_22__43_,s_r_22__42_,s_r_22__41_,s_r_22__40_,s_r_22__39_,s_r_22__38_,s_r_22__37_,
  s_r_22__36_,s_r_22__35_,s_r_22__34_,s_r_22__33_,s_r_22__32_,s_r_22__31_,
  s_r_22__30_,s_r_22__29_,s_r_22__28_,s_r_22__27_,s_r_22__26_,s_r_22__25_,s_r_22__24_,
  s_r_22__23_,s_r_22__22_,s_r_22__21_,s_r_22__20_,s_r_22__19_,s_r_22__18_,s_r_22__17_,
  s_r_22__16_,s_r_22__15_,s_r_22__14_,s_r_22__13_,s_r_22__12_,s_r_22__11_,
  s_r_22__10_,s_r_22__9_,s_r_22__8_,s_r_22__7_,s_r_22__6_,s_r_22__5_,s_r_22__4_,s_r_22__3_,
  s_r_22__2_,s_r_22__1_,s_r_22__0_,s_r_21__127_,s_r_21__126_,s_r_21__125_,
  s_r_21__124_,s_r_21__123_,s_r_21__122_,s_r_21__121_,s_r_21__120_,s_r_21__119_,
  s_r_21__118_,s_r_21__117_,s_r_21__116_,s_r_21__115_,s_r_21__114_,s_r_21__113_,s_r_21__112_,
  s_r_21__111_,s_r_21__110_,s_r_21__109_,s_r_21__108_,s_r_21__107_,s_r_21__106_,
  s_r_21__105_,s_r_21__104_,s_r_21__103_,s_r_21__102_,s_r_21__101_,s_r_21__100_,
  s_r_21__99_,s_r_21__98_,s_r_21__97_,s_r_21__96_,s_r_21__95_,s_r_21__94_,s_r_21__93_,
  s_r_21__92_,s_r_21__91_,s_r_21__90_,s_r_21__89_,s_r_21__88_,s_r_21__87_,
  s_r_21__86_,s_r_21__85_,s_r_21__84_,s_r_21__83_,s_r_21__82_,s_r_21__81_,s_r_21__80_,
  s_r_21__79_,s_r_21__78_,s_r_21__77_,s_r_21__76_,s_r_21__75_,s_r_21__74_,s_r_21__73_,
  s_r_21__72_,s_r_21__71_,s_r_21__70_,s_r_21__69_,s_r_21__68_,s_r_21__67_,
  s_r_21__66_,s_r_21__65_,s_r_21__64_,s_r_21__63_,s_r_21__62_,s_r_21__61_,s_r_21__60_,
  s_r_21__59_,s_r_21__58_,s_r_21__57_,s_r_21__56_,s_r_21__55_,s_r_21__54_,s_r_21__53_,
  s_r_21__52_,s_r_21__51_,s_r_21__50_,s_r_21__49_,s_r_21__48_,s_r_21__47_,
  s_r_21__46_,s_r_21__45_,s_r_21__44_,s_r_21__43_,s_r_21__42_,s_r_21__41_,s_r_21__40_,
  s_r_21__39_,s_r_21__38_,s_r_21__37_,s_r_21__36_,s_r_21__35_,s_r_21__34_,s_r_21__33_,
  s_r_21__32_,s_r_21__31_,s_r_21__30_,s_r_21__29_,s_r_21__28_,s_r_21__27_,
  s_r_21__26_,s_r_21__25_,s_r_21__24_,s_r_21__23_,s_r_21__22_,s_r_21__21_,s_r_21__20_,
  s_r_21__19_,s_r_21__18_,s_r_21__17_,s_r_21__16_,s_r_21__15_,s_r_21__14_,s_r_21__13_,
  s_r_21__12_,s_r_21__11_,s_r_21__10_,s_r_21__9_,s_r_21__8_,s_r_21__7_,s_r_21__6_,
  s_r_21__5_,s_r_21__4_,s_r_21__3_,s_r_21__2_,s_r_21__1_,s_r_21__0_,s_r_20__127_,
  s_r_20__126_,s_r_20__125_,s_r_20__124_,s_r_20__123_,s_r_20__122_,s_r_20__121_,
  s_r_20__120_,s_r_20__119_,s_r_20__118_,s_r_20__117_,s_r_20__116_,s_r_20__115_,
  s_r_20__114_,s_r_20__113_,s_r_20__112_,s_r_20__111_,s_r_20__110_,s_r_20__109_,
  s_r_20__108_,s_r_20__107_,s_r_20__106_,s_r_20__105_,s_r_20__104_,s_r_20__103_,
  s_r_20__102_,s_r_20__101_,s_r_20__100_,s_r_20__99_,s_r_20__98_,s_r_20__97_,s_r_20__96_,
  s_r_20__95_,s_r_20__94_,s_r_20__93_,s_r_20__92_,s_r_20__91_,s_r_20__90_,
  s_r_20__89_,s_r_20__88_,s_r_20__87_,s_r_20__86_,s_r_20__85_,s_r_20__84_,s_r_20__83_,
  s_r_20__82_,s_r_20__81_,s_r_20__80_,s_r_20__79_,s_r_20__78_,s_r_20__77_,s_r_20__76_,
  s_r_20__75_,s_r_20__74_,s_r_20__73_,s_r_20__72_,s_r_20__71_,s_r_20__70_,
  s_r_20__69_,s_r_20__68_,s_r_20__67_,s_r_20__66_,s_r_20__65_,s_r_20__64_,s_r_20__63_,
  s_r_20__62_,s_r_20__61_,s_r_20__60_,s_r_20__59_,s_r_20__58_,s_r_20__57_,s_r_20__56_,
  s_r_20__55_,s_r_20__54_,s_r_20__53_,s_r_20__52_,s_r_20__51_,s_r_20__50_,
  s_r_20__49_,s_r_20__48_,s_r_20__47_,s_r_20__46_,s_r_20__45_,s_r_20__44_,s_r_20__43_,
  s_r_20__42_,s_r_20__41_,s_r_20__40_,s_r_20__39_,s_r_20__38_,s_r_20__37_,s_r_20__36_,
  s_r_20__35_,s_r_20__34_,s_r_20__33_,s_r_20__32_,s_r_20__31_,s_r_20__30_,
  s_r_20__29_,s_r_20__28_,s_r_20__27_,s_r_20__26_,s_r_20__25_,s_r_20__24_,s_r_20__23_,
  s_r_20__22_,s_r_20__21_,s_r_20__20_,s_r_20__19_,s_r_20__18_,s_r_20__17_,s_r_20__16_,
  s_r_20__15_,s_r_20__14_,s_r_20__13_,s_r_20__12_,s_r_20__11_,s_r_20__10_,
  s_r_20__9_,s_r_20__8_,s_r_20__7_,s_r_20__6_,s_r_20__5_,s_r_20__4_,s_r_20__3_,s_r_20__2_,
  s_r_20__1_,s_r_20__0_,s_r_19__127_,s_r_19__126_,s_r_19__125_,s_r_19__124_,
  s_r_19__123_,s_r_19__122_,s_r_19__121_,s_r_19__120_,s_r_19__119_,s_r_19__118_,
  s_r_19__117_,s_r_19__116_,s_r_19__115_,s_r_19__114_,s_r_19__113_,s_r_19__112_,
  s_r_19__111_,s_r_19__110_,s_r_19__109_,s_r_19__108_,s_r_19__107_,s_r_19__106_,s_r_19__105_,
  s_r_19__104_,s_r_19__103_,s_r_19__102_,s_r_19__101_,s_r_19__100_,s_r_19__99_,
  s_r_19__98_,s_r_19__97_,s_r_19__96_,s_r_19__95_,s_r_19__94_,s_r_19__93_,s_r_19__92_,
  s_r_19__91_,s_r_19__90_,s_r_19__89_,s_r_19__88_,s_r_19__87_,s_r_19__86_,
  s_r_19__85_,s_r_19__84_,s_r_19__83_,s_r_19__82_,s_r_19__81_,s_r_19__80_,s_r_19__79_,
  s_r_19__78_,s_r_19__77_,s_r_19__76_,s_r_19__75_,s_r_19__74_,s_r_19__73_,s_r_19__72_,
  s_r_19__71_,s_r_19__70_,s_r_19__69_,s_r_19__68_,s_r_19__67_,s_r_19__66_,
  s_r_19__65_,s_r_19__64_,s_r_19__63_,s_r_19__62_,s_r_19__61_,s_r_19__60_,s_r_19__59_,
  s_r_19__58_,s_r_19__57_,s_r_19__56_,s_r_19__55_,s_r_19__54_,s_r_19__53_,s_r_19__52_,
  s_r_19__51_,s_r_19__50_,s_r_19__49_,s_r_19__48_,s_r_19__47_,s_r_19__46_,
  s_r_19__45_,s_r_19__44_,s_r_19__43_,s_r_19__42_,s_r_19__41_,s_r_19__40_,s_r_19__39_,
  s_r_19__38_,s_r_19__37_,s_r_19__36_,s_r_19__35_,s_r_19__34_,s_r_19__33_,s_r_19__32_,
  s_r_19__31_,s_r_19__30_,s_r_19__29_,s_r_19__28_,s_r_19__27_,s_r_19__26_,
  s_r_19__25_,s_r_19__24_,s_r_19__23_,s_r_19__22_,s_r_19__21_,s_r_19__20_,s_r_19__19_,
  s_r_19__18_,s_r_19__17_,s_r_19__16_,s_r_19__15_,s_r_19__14_,s_r_19__13_,s_r_19__12_,
  s_r_19__11_,s_r_19__10_,s_r_19__9_,s_r_19__8_,s_r_19__7_,s_r_19__6_,s_r_19__5_,
  s_r_19__4_,s_r_19__3_,s_r_19__2_,s_r_19__1_,s_r_19__0_,prod_accum_22__23_,
  prod_accum_22__22_,prod_accum_22__21_,prod_accum_22__20_,prod_accum_22__19_,
  prod_accum_22__18_,prod_accum_22__17_,prod_accum_22__16_,prod_accum_22__15_,
  prod_accum_22__14_,prod_accum_22__13_,prod_accum_22__12_,prod_accum_22__11_,prod_accum_22__10_,
  prod_accum_22__9_,prod_accum_22__8_,prod_accum_22__7_,prod_accum_22__6_,
  prod_accum_22__5_,prod_accum_22__4_,prod_accum_22__3_,prod_accum_22__2_,
  prod_accum_22__1_,prod_accum_22__0_,prod_accum_21__22_,prod_accum_21__21_,prod_accum_21__20_,
  prod_accum_21__19_,prod_accum_21__18_,prod_accum_21__17_,prod_accum_21__16_,
  prod_accum_21__15_,prod_accum_21__14_,prod_accum_21__13_,prod_accum_21__12_,
  prod_accum_21__11_,prod_accum_21__10_,prod_accum_21__9_,prod_accum_21__8_,
  prod_accum_21__7_,prod_accum_21__6_,prod_accum_21__5_,prod_accum_21__4_,prod_accum_21__3_,
  prod_accum_21__2_,prod_accum_21__1_,prod_accum_21__0_,prod_accum_20__21_,
  prod_accum_20__20_,prod_accum_20__19_,prod_accum_20__18_,prod_accum_20__17_,
  prod_accum_20__16_,prod_accum_20__15_,prod_accum_20__14_,prod_accum_20__13_,prod_accum_20__12_,
  prod_accum_20__11_,prod_accum_20__10_,prod_accum_20__9_,prod_accum_20__8_,
  prod_accum_20__7_,prod_accum_20__6_,prod_accum_20__5_,prod_accum_20__4_,
  prod_accum_20__3_,prod_accum_20__2_,prod_accum_20__1_,prod_accum_20__0_,prod_accum_19__20_,
  prod_accum_19__19_,prod_accum_19__18_,prod_accum_19__17_,prod_accum_19__16_,
  prod_accum_19__15_,prod_accum_19__14_,prod_accum_19__13_,prod_accum_19__12_,
  prod_accum_19__11_,prod_accum_19__10_,prod_accum_19__9_,prod_accum_19__8_,prod_accum_19__7_,
  prod_accum_19__6_,prod_accum_19__5_,prod_accum_19__4_,prod_accum_19__3_,
  prod_accum_19__2_,prod_accum_19__1_,prod_accum_19__0_,s_r_26__127_,s_r_26__126_,
  s_r_26__125_,s_r_26__124_,s_r_26__123_,s_r_26__122_,s_r_26__121_,s_r_26__120_,
  s_r_26__119_,s_r_26__118_,s_r_26__117_,s_r_26__116_,s_r_26__115_,s_r_26__114_,s_r_26__113_,
  s_r_26__112_,s_r_26__111_,s_r_26__110_,s_r_26__109_,s_r_26__108_,s_r_26__107_,
  s_r_26__106_,s_r_26__105_,s_r_26__104_,s_r_26__103_,s_r_26__102_,s_r_26__101_,
  s_r_26__100_,s_r_26__99_,s_r_26__98_,s_r_26__97_,s_r_26__96_,s_r_26__95_,s_r_26__94_,
  s_r_26__93_,s_r_26__92_,s_r_26__91_,s_r_26__90_,s_r_26__89_,s_r_26__88_,
  s_r_26__87_,s_r_26__86_,s_r_26__85_,s_r_26__84_,s_r_26__83_,s_r_26__82_,s_r_26__81_,
  s_r_26__80_,s_r_26__79_,s_r_26__78_,s_r_26__77_,s_r_26__76_,s_r_26__75_,s_r_26__74_,
  s_r_26__73_,s_r_26__72_,s_r_26__71_,s_r_26__70_,s_r_26__69_,s_r_26__68_,
  s_r_26__67_,s_r_26__66_,s_r_26__65_,s_r_26__64_,s_r_26__63_,s_r_26__62_,s_r_26__61_,
  s_r_26__60_,s_r_26__59_,s_r_26__58_,s_r_26__57_,s_r_26__56_,s_r_26__55_,s_r_26__54_,
  s_r_26__53_,s_r_26__52_,s_r_26__51_,s_r_26__50_,s_r_26__49_,s_r_26__48_,
  s_r_26__47_,s_r_26__46_,s_r_26__45_,s_r_26__44_,s_r_26__43_,s_r_26__42_,s_r_26__41_,
  s_r_26__40_,s_r_26__39_,s_r_26__38_,s_r_26__37_,s_r_26__36_,s_r_26__35_,s_r_26__34_,
  s_r_26__33_,s_r_26__32_,s_r_26__31_,s_r_26__30_,s_r_26__29_,s_r_26__28_,
  s_r_26__27_,s_r_26__26_,s_r_26__25_,s_r_26__24_,s_r_26__23_,s_r_26__22_,s_r_26__21_,
  s_r_26__20_,s_r_26__19_,s_r_26__18_,s_r_26__17_,s_r_26__16_,s_r_26__15_,s_r_26__14_,
  s_r_26__13_,s_r_26__12_,s_r_26__11_,s_r_26__10_,s_r_26__9_,s_r_26__8_,
  s_r_26__7_,s_r_26__6_,s_r_26__5_,s_r_26__4_,s_r_26__3_,s_r_26__2_,s_r_26__1_,s_r_26__0_,
  s_r_25__127_,s_r_25__126_,s_r_25__125_,s_r_25__124_,s_r_25__123_,s_r_25__122_,
  s_r_25__121_,s_r_25__120_,s_r_25__119_,s_r_25__118_,s_r_25__117_,s_r_25__116_,
  s_r_25__115_,s_r_25__114_,s_r_25__113_,s_r_25__112_,s_r_25__111_,s_r_25__110_,
  s_r_25__109_,s_r_25__108_,s_r_25__107_,s_r_25__106_,s_r_25__105_,s_r_25__104_,
  s_r_25__103_,s_r_25__102_,s_r_25__101_,s_r_25__100_,s_r_25__99_,s_r_25__98_,s_r_25__97_,
  s_r_25__96_,s_r_25__95_,s_r_25__94_,s_r_25__93_,s_r_25__92_,s_r_25__91_,
  s_r_25__90_,s_r_25__89_,s_r_25__88_,s_r_25__87_,s_r_25__86_,s_r_25__85_,s_r_25__84_,
  s_r_25__83_,s_r_25__82_,s_r_25__81_,s_r_25__80_,s_r_25__79_,s_r_25__78_,s_r_25__77_,
  s_r_25__76_,s_r_25__75_,s_r_25__74_,s_r_25__73_,s_r_25__72_,s_r_25__71_,
  s_r_25__70_,s_r_25__69_,s_r_25__68_,s_r_25__67_,s_r_25__66_,s_r_25__65_,s_r_25__64_,
  s_r_25__63_,s_r_25__62_,s_r_25__61_,s_r_25__60_,s_r_25__59_,s_r_25__58_,s_r_25__57_,
  s_r_25__56_,s_r_25__55_,s_r_25__54_,s_r_25__53_,s_r_25__52_,s_r_25__51_,
  s_r_25__50_,s_r_25__49_,s_r_25__48_,s_r_25__47_,s_r_25__46_,s_r_25__45_,s_r_25__44_,
  s_r_25__43_,s_r_25__42_,s_r_25__41_,s_r_25__40_,s_r_25__39_,s_r_25__38_,s_r_25__37_,
  s_r_25__36_,s_r_25__35_,s_r_25__34_,s_r_25__33_,s_r_25__32_,s_r_25__31_,
  s_r_25__30_,s_r_25__29_,s_r_25__28_,s_r_25__27_,s_r_25__26_,s_r_25__25_,s_r_25__24_,
  s_r_25__23_,s_r_25__22_,s_r_25__21_,s_r_25__20_,s_r_25__19_,s_r_25__18_,s_r_25__17_,
  s_r_25__16_,s_r_25__15_,s_r_25__14_,s_r_25__13_,s_r_25__12_,s_r_25__11_,
  s_r_25__10_,s_r_25__9_,s_r_25__8_,s_r_25__7_,s_r_25__6_,s_r_25__5_,s_r_25__4_,s_r_25__3_,
  s_r_25__2_,s_r_25__1_,s_r_25__0_,s_r_24__127_,s_r_24__126_,s_r_24__125_,
  s_r_24__124_,s_r_24__123_,s_r_24__122_,s_r_24__121_,s_r_24__120_,s_r_24__119_,
  s_r_24__118_,s_r_24__117_,s_r_24__116_,s_r_24__115_,s_r_24__114_,s_r_24__113_,s_r_24__112_,
  s_r_24__111_,s_r_24__110_,s_r_24__109_,s_r_24__108_,s_r_24__107_,s_r_24__106_,
  s_r_24__105_,s_r_24__104_,s_r_24__103_,s_r_24__102_,s_r_24__101_,s_r_24__100_,
  s_r_24__99_,s_r_24__98_,s_r_24__97_,s_r_24__96_,s_r_24__95_,s_r_24__94_,s_r_24__93_,
  s_r_24__92_,s_r_24__91_,s_r_24__90_,s_r_24__89_,s_r_24__88_,s_r_24__87_,
  s_r_24__86_,s_r_24__85_,s_r_24__84_,s_r_24__83_,s_r_24__82_,s_r_24__81_,s_r_24__80_,
  s_r_24__79_,s_r_24__78_,s_r_24__77_,s_r_24__76_,s_r_24__75_,s_r_24__74_,s_r_24__73_,
  s_r_24__72_,s_r_24__71_,s_r_24__70_,s_r_24__69_,s_r_24__68_,s_r_24__67_,
  s_r_24__66_,s_r_24__65_,s_r_24__64_,s_r_24__63_,s_r_24__62_,s_r_24__61_,s_r_24__60_,
  s_r_24__59_,s_r_24__58_,s_r_24__57_,s_r_24__56_,s_r_24__55_,s_r_24__54_,s_r_24__53_,
  s_r_24__52_,s_r_24__51_,s_r_24__50_,s_r_24__49_,s_r_24__48_,s_r_24__47_,
  s_r_24__46_,s_r_24__45_,s_r_24__44_,s_r_24__43_,s_r_24__42_,s_r_24__41_,s_r_24__40_,
  s_r_24__39_,s_r_24__38_,s_r_24__37_,s_r_24__36_,s_r_24__35_,s_r_24__34_,s_r_24__33_,
  s_r_24__32_,s_r_24__31_,s_r_24__30_,s_r_24__29_,s_r_24__28_,s_r_24__27_,
  s_r_24__26_,s_r_24__25_,s_r_24__24_,s_r_24__23_,s_r_24__22_,s_r_24__21_,s_r_24__20_,
  s_r_24__19_,s_r_24__18_,s_r_24__17_,s_r_24__16_,s_r_24__15_,s_r_24__14_,s_r_24__13_,
  s_r_24__12_,s_r_24__11_,s_r_24__10_,s_r_24__9_,s_r_24__8_,s_r_24__7_,s_r_24__6_,
  s_r_24__5_,s_r_24__4_,s_r_24__3_,s_r_24__2_,s_r_24__1_,s_r_24__0_,s_r_23__127_,
  s_r_23__126_,s_r_23__125_,s_r_23__124_,s_r_23__123_,s_r_23__122_,s_r_23__121_,
  s_r_23__120_,s_r_23__119_,s_r_23__118_,s_r_23__117_,s_r_23__116_,s_r_23__115_,
  s_r_23__114_,s_r_23__113_,s_r_23__112_,s_r_23__111_,s_r_23__110_,s_r_23__109_,
  s_r_23__108_,s_r_23__107_,s_r_23__106_,s_r_23__105_,s_r_23__104_,s_r_23__103_,
  s_r_23__102_,s_r_23__101_,s_r_23__100_,s_r_23__99_,s_r_23__98_,s_r_23__97_,s_r_23__96_,
  s_r_23__95_,s_r_23__94_,s_r_23__93_,s_r_23__92_,s_r_23__91_,s_r_23__90_,
  s_r_23__89_,s_r_23__88_,s_r_23__87_,s_r_23__86_,s_r_23__85_,s_r_23__84_,s_r_23__83_,
  s_r_23__82_,s_r_23__81_,s_r_23__80_,s_r_23__79_,s_r_23__78_,s_r_23__77_,s_r_23__76_,
  s_r_23__75_,s_r_23__74_,s_r_23__73_,s_r_23__72_,s_r_23__71_,s_r_23__70_,
  s_r_23__69_,s_r_23__68_,s_r_23__67_,s_r_23__66_,s_r_23__65_,s_r_23__64_,s_r_23__63_,
  s_r_23__62_,s_r_23__61_,s_r_23__60_,s_r_23__59_,s_r_23__58_,s_r_23__57_,s_r_23__56_,
  s_r_23__55_,s_r_23__54_,s_r_23__53_,s_r_23__52_,s_r_23__51_,s_r_23__50_,
  s_r_23__49_,s_r_23__48_,s_r_23__47_,s_r_23__46_,s_r_23__45_,s_r_23__44_,s_r_23__43_,
  s_r_23__42_,s_r_23__41_,s_r_23__40_,s_r_23__39_,s_r_23__38_,s_r_23__37_,s_r_23__36_,
  s_r_23__35_,s_r_23__34_,s_r_23__33_,s_r_23__32_,s_r_23__31_,s_r_23__30_,
  s_r_23__29_,s_r_23__28_,s_r_23__27_,s_r_23__26_,s_r_23__25_,s_r_23__24_,s_r_23__23_,
  s_r_23__22_,s_r_23__21_,s_r_23__20_,s_r_23__19_,s_r_23__18_,s_r_23__17_,s_r_23__16_,
  s_r_23__15_,s_r_23__14_,s_r_23__13_,s_r_23__12_,s_r_23__11_,s_r_23__10_,
  s_r_23__9_,s_r_23__8_,s_r_23__7_,s_r_23__6_,s_r_23__5_,s_r_23__4_,s_r_23__3_,s_r_23__2_,
  s_r_23__1_,s_r_23__0_,prod_accum_26__27_,prod_accum_26__26_,prod_accum_26__25_,
  prod_accum_26__24_,prod_accum_26__23_,prod_accum_26__22_,prod_accum_26__21_,
  prod_accum_26__20_,prod_accum_26__19_,prod_accum_26__18_,prod_accum_26__17_,
  prod_accum_26__16_,prod_accum_26__15_,prod_accum_26__14_,prod_accum_26__13_,
  prod_accum_26__12_,prod_accum_26__11_,prod_accum_26__10_,prod_accum_26__9_,prod_accum_26__8_,
  prod_accum_26__7_,prod_accum_26__6_,prod_accum_26__5_,prod_accum_26__4_,
  prod_accum_26__3_,prod_accum_26__2_,prod_accum_26__1_,prod_accum_26__0_,
  prod_accum_25__26_,prod_accum_25__25_,prod_accum_25__24_,prod_accum_25__23_,prod_accum_25__22_,
  prod_accum_25__21_,prod_accum_25__20_,prod_accum_25__19_,prod_accum_25__18_,
  prod_accum_25__17_,prod_accum_25__16_,prod_accum_25__15_,prod_accum_25__14_,
  prod_accum_25__13_,prod_accum_25__12_,prod_accum_25__11_,prod_accum_25__10_,
  prod_accum_25__9_,prod_accum_25__8_,prod_accum_25__7_,prod_accum_25__6_,prod_accum_25__5_,
  prod_accum_25__4_,prod_accum_25__3_,prod_accum_25__2_,prod_accum_25__1_,
  prod_accum_25__0_,prod_accum_24__25_,prod_accum_24__24_,prod_accum_24__23_,
  prod_accum_24__22_,prod_accum_24__21_,prod_accum_24__20_,prod_accum_24__19_,prod_accum_24__18_,
  prod_accum_24__17_,prod_accum_24__16_,prod_accum_24__15_,prod_accum_24__14_,
  prod_accum_24__13_,prod_accum_24__12_,prod_accum_24__11_,prod_accum_24__10_,
  prod_accum_24__9_,prod_accum_24__8_,prod_accum_24__7_,prod_accum_24__6_,prod_accum_24__5_,
  prod_accum_24__4_,prod_accum_24__3_,prod_accum_24__2_,prod_accum_24__1_,
  prod_accum_24__0_,prod_accum_23__24_,prod_accum_23__23_,prod_accum_23__22_,
  prod_accum_23__21_,prod_accum_23__20_,prod_accum_23__19_,prod_accum_23__18_,
  prod_accum_23__17_,prod_accum_23__16_,prod_accum_23__15_,prod_accum_23__14_,prod_accum_23__13_,
  prod_accum_23__12_,prod_accum_23__11_,prod_accum_23__10_,prod_accum_23__9_,
  prod_accum_23__8_,prod_accum_23__7_,prod_accum_23__6_,prod_accum_23__5_,
  prod_accum_23__4_,prod_accum_23__3_,prod_accum_23__2_,prod_accum_23__1_,prod_accum_23__0_,
  s_r_30__127_,s_r_30__126_,s_r_30__125_,s_r_30__124_,s_r_30__123_,s_r_30__122_,
  s_r_30__121_,s_r_30__120_,s_r_30__119_,s_r_30__118_,s_r_30__117_,s_r_30__116_,
  s_r_30__115_,s_r_30__114_,s_r_30__113_,s_r_30__112_,s_r_30__111_,s_r_30__110_,
  s_r_30__109_,s_r_30__108_,s_r_30__107_,s_r_30__106_,s_r_30__105_,s_r_30__104_,s_r_30__103_,
  s_r_30__102_,s_r_30__101_,s_r_30__100_,s_r_30__99_,s_r_30__98_,s_r_30__97_,
  s_r_30__96_,s_r_30__95_,s_r_30__94_,s_r_30__93_,s_r_30__92_,s_r_30__91_,s_r_30__90_,
  s_r_30__89_,s_r_30__88_,s_r_30__87_,s_r_30__86_,s_r_30__85_,s_r_30__84_,
  s_r_30__83_,s_r_30__82_,s_r_30__81_,s_r_30__80_,s_r_30__79_,s_r_30__78_,s_r_30__77_,
  s_r_30__76_,s_r_30__75_,s_r_30__74_,s_r_30__73_,s_r_30__72_,s_r_30__71_,s_r_30__70_,
  s_r_30__69_,s_r_30__68_,s_r_30__67_,s_r_30__66_,s_r_30__65_,s_r_30__64_,
  s_r_30__63_,s_r_30__62_,s_r_30__61_,s_r_30__60_,s_r_30__59_,s_r_30__58_,s_r_30__57_,
  s_r_30__56_,s_r_30__55_,s_r_30__54_,s_r_30__53_,s_r_30__52_,s_r_30__51_,s_r_30__50_,
  s_r_30__49_,s_r_30__48_,s_r_30__47_,s_r_30__46_,s_r_30__45_,s_r_30__44_,
  s_r_30__43_,s_r_30__42_,s_r_30__41_,s_r_30__40_,s_r_30__39_,s_r_30__38_,s_r_30__37_,
  s_r_30__36_,s_r_30__35_,s_r_30__34_,s_r_30__33_,s_r_30__32_,s_r_30__31_,s_r_30__30_,
  s_r_30__29_,s_r_30__28_,s_r_30__27_,s_r_30__26_,s_r_30__25_,s_r_30__24_,
  s_r_30__23_,s_r_30__22_,s_r_30__21_,s_r_30__20_,s_r_30__19_,s_r_30__18_,s_r_30__17_,
  s_r_30__16_,s_r_30__15_,s_r_30__14_,s_r_30__13_,s_r_30__12_,s_r_30__11_,s_r_30__10_,
  s_r_30__9_,s_r_30__8_,s_r_30__7_,s_r_30__6_,s_r_30__5_,s_r_30__4_,s_r_30__3_,
  s_r_30__2_,s_r_30__1_,s_r_30__0_,s_r_29__127_,s_r_29__126_,s_r_29__125_,s_r_29__124_,
  s_r_29__123_,s_r_29__122_,s_r_29__121_,s_r_29__120_,s_r_29__119_,s_r_29__118_,
  s_r_29__117_,s_r_29__116_,s_r_29__115_,s_r_29__114_,s_r_29__113_,s_r_29__112_,
  s_r_29__111_,s_r_29__110_,s_r_29__109_,s_r_29__108_,s_r_29__107_,s_r_29__106_,
  s_r_29__105_,s_r_29__104_,s_r_29__103_,s_r_29__102_,s_r_29__101_,s_r_29__100_,
  s_r_29__99_,s_r_29__98_,s_r_29__97_,s_r_29__96_,s_r_29__95_,s_r_29__94_,s_r_29__93_,
  s_r_29__92_,s_r_29__91_,s_r_29__90_,s_r_29__89_,s_r_29__88_,s_r_29__87_,s_r_29__86_,
  s_r_29__85_,s_r_29__84_,s_r_29__83_,s_r_29__82_,s_r_29__81_,s_r_29__80_,
  s_r_29__79_,s_r_29__78_,s_r_29__77_,s_r_29__76_,s_r_29__75_,s_r_29__74_,s_r_29__73_,
  s_r_29__72_,s_r_29__71_,s_r_29__70_,s_r_29__69_,s_r_29__68_,s_r_29__67_,s_r_29__66_,
  s_r_29__65_,s_r_29__64_,s_r_29__63_,s_r_29__62_,s_r_29__61_,s_r_29__60_,
  s_r_29__59_,s_r_29__58_,s_r_29__57_,s_r_29__56_,s_r_29__55_,s_r_29__54_,s_r_29__53_,
  s_r_29__52_,s_r_29__51_,s_r_29__50_,s_r_29__49_,s_r_29__48_,s_r_29__47_,s_r_29__46_,
  s_r_29__45_,s_r_29__44_,s_r_29__43_,s_r_29__42_,s_r_29__41_,s_r_29__40_,
  s_r_29__39_,s_r_29__38_,s_r_29__37_,s_r_29__36_,s_r_29__35_,s_r_29__34_,s_r_29__33_,
  s_r_29__32_,s_r_29__31_,s_r_29__30_,s_r_29__29_,s_r_29__28_,s_r_29__27_,s_r_29__26_,
  s_r_29__25_,s_r_29__24_,s_r_29__23_,s_r_29__22_,s_r_29__21_,s_r_29__20_,
  s_r_29__19_,s_r_29__18_,s_r_29__17_,s_r_29__16_,s_r_29__15_,s_r_29__14_,s_r_29__13_,
  s_r_29__12_,s_r_29__11_,s_r_29__10_,s_r_29__9_,s_r_29__8_,s_r_29__7_,s_r_29__6_,
  s_r_29__5_,s_r_29__4_,s_r_29__3_,s_r_29__2_,s_r_29__1_,s_r_29__0_,s_r_28__127_,
  s_r_28__126_,s_r_28__125_,s_r_28__124_,s_r_28__123_,s_r_28__122_,s_r_28__121_,
  s_r_28__120_,s_r_28__119_,s_r_28__118_,s_r_28__117_,s_r_28__116_,s_r_28__115_,
  s_r_28__114_,s_r_28__113_,s_r_28__112_,s_r_28__111_,s_r_28__110_,s_r_28__109_,
  s_r_28__108_,s_r_28__107_,s_r_28__106_,s_r_28__105_,s_r_28__104_,s_r_28__103_,s_r_28__102_,
  s_r_28__101_,s_r_28__100_,s_r_28__99_,s_r_28__98_,s_r_28__97_,s_r_28__96_,
  s_r_28__95_,s_r_28__94_,s_r_28__93_,s_r_28__92_,s_r_28__91_,s_r_28__90_,s_r_28__89_,
  s_r_28__88_,s_r_28__87_,s_r_28__86_,s_r_28__85_,s_r_28__84_,s_r_28__83_,
  s_r_28__82_,s_r_28__81_,s_r_28__80_,s_r_28__79_,s_r_28__78_,s_r_28__77_,s_r_28__76_,
  s_r_28__75_,s_r_28__74_,s_r_28__73_,s_r_28__72_,s_r_28__71_,s_r_28__70_,s_r_28__69_,
  s_r_28__68_,s_r_28__67_,s_r_28__66_,s_r_28__65_,s_r_28__64_,s_r_28__63_,
  s_r_28__62_,s_r_28__61_,s_r_28__60_,s_r_28__59_,s_r_28__58_,s_r_28__57_,s_r_28__56_,
  s_r_28__55_,s_r_28__54_,s_r_28__53_,s_r_28__52_,s_r_28__51_,s_r_28__50_,s_r_28__49_,
  s_r_28__48_,s_r_28__47_,s_r_28__46_,s_r_28__45_,s_r_28__44_,s_r_28__43_,
  s_r_28__42_,s_r_28__41_,s_r_28__40_,s_r_28__39_,s_r_28__38_,s_r_28__37_,s_r_28__36_,
  s_r_28__35_,s_r_28__34_,s_r_28__33_,s_r_28__32_,s_r_28__31_,s_r_28__30_,s_r_28__29_,
  s_r_28__28_,s_r_28__27_,s_r_28__26_,s_r_28__25_,s_r_28__24_,s_r_28__23_,
  s_r_28__22_,s_r_28__21_,s_r_28__20_,s_r_28__19_,s_r_28__18_,s_r_28__17_,s_r_28__16_,
  s_r_28__15_,s_r_28__14_,s_r_28__13_,s_r_28__12_,s_r_28__11_,s_r_28__10_,s_r_28__9_,
  s_r_28__8_,s_r_28__7_,s_r_28__6_,s_r_28__5_,s_r_28__4_,s_r_28__3_,s_r_28__2_,
  s_r_28__1_,s_r_28__0_,s_r_27__127_,s_r_27__126_,s_r_27__125_,s_r_27__124_,
  s_r_27__123_,s_r_27__122_,s_r_27__121_,s_r_27__120_,s_r_27__119_,s_r_27__118_,s_r_27__117_,
  s_r_27__116_,s_r_27__115_,s_r_27__114_,s_r_27__113_,s_r_27__112_,s_r_27__111_,
  s_r_27__110_,s_r_27__109_,s_r_27__108_,s_r_27__107_,s_r_27__106_,s_r_27__105_,
  s_r_27__104_,s_r_27__103_,s_r_27__102_,s_r_27__101_,s_r_27__100_,s_r_27__99_,
  s_r_27__98_,s_r_27__97_,s_r_27__96_,s_r_27__95_,s_r_27__94_,s_r_27__93_,s_r_27__92_,
  s_r_27__91_,s_r_27__90_,s_r_27__89_,s_r_27__88_,s_r_27__87_,s_r_27__86_,s_r_27__85_,
  s_r_27__84_,s_r_27__83_,s_r_27__82_,s_r_27__81_,s_r_27__80_,s_r_27__79_,
  s_r_27__78_,s_r_27__77_,s_r_27__76_,s_r_27__75_,s_r_27__74_,s_r_27__73_,s_r_27__72_,
  s_r_27__71_,s_r_27__70_,s_r_27__69_,s_r_27__68_,s_r_27__67_,s_r_27__66_,s_r_27__65_,
  s_r_27__64_,s_r_27__63_,s_r_27__62_,s_r_27__61_,s_r_27__60_,s_r_27__59_,
  s_r_27__58_,s_r_27__57_,s_r_27__56_,s_r_27__55_,s_r_27__54_,s_r_27__53_,s_r_27__52_,
  s_r_27__51_,s_r_27__50_,s_r_27__49_,s_r_27__48_,s_r_27__47_,s_r_27__46_,s_r_27__45_,
  s_r_27__44_,s_r_27__43_,s_r_27__42_,s_r_27__41_,s_r_27__40_,s_r_27__39_,
  s_r_27__38_,s_r_27__37_,s_r_27__36_,s_r_27__35_,s_r_27__34_,s_r_27__33_,s_r_27__32_,
  s_r_27__31_,s_r_27__30_,s_r_27__29_,s_r_27__28_,s_r_27__27_,s_r_27__26_,s_r_27__25_,
  s_r_27__24_,s_r_27__23_,s_r_27__22_,s_r_27__21_,s_r_27__20_,s_r_27__19_,
  s_r_27__18_,s_r_27__17_,s_r_27__16_,s_r_27__15_,s_r_27__14_,s_r_27__13_,s_r_27__12_,
  s_r_27__11_,s_r_27__10_,s_r_27__9_,s_r_27__8_,s_r_27__7_,s_r_27__6_,s_r_27__5_,
  s_r_27__4_,s_r_27__3_,s_r_27__2_,s_r_27__1_,s_r_27__0_,prod_accum_30__31_,
  prod_accum_30__30_,prod_accum_30__29_,prod_accum_30__28_,prod_accum_30__27_,
  prod_accum_30__26_,prod_accum_30__25_,prod_accum_30__24_,prod_accum_30__23_,prod_accum_30__22_,
  prod_accum_30__21_,prod_accum_30__20_,prod_accum_30__19_,prod_accum_30__18_,
  prod_accum_30__17_,prod_accum_30__16_,prod_accum_30__15_,prod_accum_30__14_,
  prod_accum_30__13_,prod_accum_30__12_,prod_accum_30__11_,prod_accum_30__10_,
  prod_accum_30__9_,prod_accum_30__8_,prod_accum_30__7_,prod_accum_30__6_,prod_accum_30__5_,
  prod_accum_30__4_,prod_accum_30__3_,prod_accum_30__2_,prod_accum_30__1_,
  prod_accum_30__0_,prod_accum_29__30_,prod_accum_29__29_,prod_accum_29__28_,
  prod_accum_29__27_,prod_accum_29__26_,prod_accum_29__25_,prod_accum_29__24_,prod_accum_29__23_,
  prod_accum_29__22_,prod_accum_29__21_,prod_accum_29__20_,prod_accum_29__19_,
  prod_accum_29__18_,prod_accum_29__17_,prod_accum_29__16_,prod_accum_29__15_,
  prod_accum_29__14_,prod_accum_29__13_,prod_accum_29__12_,prod_accum_29__11_,
  prod_accum_29__10_,prod_accum_29__9_,prod_accum_29__8_,prod_accum_29__7_,prod_accum_29__6_,
  prod_accum_29__5_,prod_accum_29__4_,prod_accum_29__3_,prod_accum_29__2_,
  prod_accum_29__1_,prod_accum_29__0_,prod_accum_28__29_,prod_accum_28__28_,
  prod_accum_28__27_,prod_accum_28__26_,prod_accum_28__25_,prod_accum_28__24_,prod_accum_28__23_,
  prod_accum_28__22_,prod_accum_28__21_,prod_accum_28__20_,prod_accum_28__19_,
  prod_accum_28__18_,prod_accum_28__17_,prod_accum_28__16_,prod_accum_28__15_,
  prod_accum_28__14_,prod_accum_28__13_,prod_accum_28__12_,prod_accum_28__11_,
  prod_accum_28__10_,prod_accum_28__9_,prod_accum_28__8_,prod_accum_28__7_,prod_accum_28__6_,
  prod_accum_28__5_,prod_accum_28__4_,prod_accum_28__3_,prod_accum_28__2_,
  prod_accum_28__1_,prod_accum_28__0_,prod_accum_27__28_,prod_accum_27__27_,
  prod_accum_27__26_,prod_accum_27__25_,prod_accum_27__24_,prod_accum_27__23_,prod_accum_27__22_,
  prod_accum_27__21_,prod_accum_27__20_,prod_accum_27__19_,prod_accum_27__18_,
  prod_accum_27__17_,prod_accum_27__16_,prod_accum_27__15_,prod_accum_27__14_,
  prod_accum_27__13_,prod_accum_27__12_,prod_accum_27__11_,prod_accum_27__10_,
  prod_accum_27__9_,prod_accum_27__8_,prod_accum_27__7_,prod_accum_27__6_,prod_accum_27__5_,
  prod_accum_27__4_,prod_accum_27__3_,prod_accum_27__2_,prod_accum_27__1_,
  prod_accum_27__0_,s_r_34__127_,s_r_34__126_,s_r_34__125_,s_r_34__124_,s_r_34__123_,
  s_r_34__122_,s_r_34__121_,s_r_34__120_,s_r_34__119_,s_r_34__118_,s_r_34__117_,
  s_r_34__116_,s_r_34__115_,s_r_34__114_,s_r_34__113_,s_r_34__112_,s_r_34__111_,
  s_r_34__110_,s_r_34__109_,s_r_34__108_,s_r_34__107_,s_r_34__106_,s_r_34__105_,s_r_34__104_,
  s_r_34__103_,s_r_34__102_,s_r_34__101_,s_r_34__100_,s_r_34__99_,s_r_34__98_,
  s_r_34__97_,s_r_34__96_,s_r_34__95_,s_r_34__94_,s_r_34__93_,s_r_34__92_,s_r_34__91_,
  s_r_34__90_,s_r_34__89_,s_r_34__88_,s_r_34__87_,s_r_34__86_,s_r_34__85_,
  s_r_34__84_,s_r_34__83_,s_r_34__82_,s_r_34__81_,s_r_34__80_,s_r_34__79_,s_r_34__78_,
  s_r_34__77_,s_r_34__76_,s_r_34__75_,s_r_34__74_,s_r_34__73_,s_r_34__72_,s_r_34__71_,
  s_r_34__70_,s_r_34__69_,s_r_34__68_,s_r_34__67_,s_r_34__66_,s_r_34__65_,
  s_r_34__64_,s_r_34__63_,s_r_34__62_,s_r_34__61_,s_r_34__60_,s_r_34__59_,s_r_34__58_,
  s_r_34__57_,s_r_34__56_,s_r_34__55_,s_r_34__54_,s_r_34__53_,s_r_34__52_,s_r_34__51_,
  s_r_34__50_,s_r_34__49_,s_r_34__48_,s_r_34__47_,s_r_34__46_,s_r_34__45_,
  s_r_34__44_,s_r_34__43_,s_r_34__42_,s_r_34__41_,s_r_34__40_,s_r_34__39_,s_r_34__38_,
  s_r_34__37_,s_r_34__36_,s_r_34__35_,s_r_34__34_,s_r_34__33_,s_r_34__32_,s_r_34__31_,
  s_r_34__30_,s_r_34__29_,s_r_34__28_,s_r_34__27_,s_r_34__26_,s_r_34__25_,
  s_r_34__24_,s_r_34__23_,s_r_34__22_,s_r_34__21_,s_r_34__20_,s_r_34__19_,s_r_34__18_,
  s_r_34__17_,s_r_34__16_,s_r_34__15_,s_r_34__14_,s_r_34__13_,s_r_34__12_,s_r_34__11_,
  s_r_34__10_,s_r_34__9_,s_r_34__8_,s_r_34__7_,s_r_34__6_,s_r_34__5_,s_r_34__4_,
  s_r_34__3_,s_r_34__2_,s_r_34__1_,s_r_34__0_,s_r_33__127_,s_r_33__126_,
  s_r_33__125_,s_r_33__124_,s_r_33__123_,s_r_33__122_,s_r_33__121_,s_r_33__120_,s_r_33__119_,
  s_r_33__118_,s_r_33__117_,s_r_33__116_,s_r_33__115_,s_r_33__114_,s_r_33__113_,
  s_r_33__112_,s_r_33__111_,s_r_33__110_,s_r_33__109_,s_r_33__108_,s_r_33__107_,
  s_r_33__106_,s_r_33__105_,s_r_33__104_,s_r_33__103_,s_r_33__102_,s_r_33__101_,
  s_r_33__100_,s_r_33__99_,s_r_33__98_,s_r_33__97_,s_r_33__96_,s_r_33__95_,s_r_33__94_,
  s_r_33__93_,s_r_33__92_,s_r_33__91_,s_r_33__90_,s_r_33__89_,s_r_33__88_,
  s_r_33__87_,s_r_33__86_,s_r_33__85_,s_r_33__84_,s_r_33__83_,s_r_33__82_,s_r_33__81_,
  s_r_33__80_,s_r_33__79_,s_r_33__78_,s_r_33__77_,s_r_33__76_,s_r_33__75_,s_r_33__74_,
  s_r_33__73_,s_r_33__72_,s_r_33__71_,s_r_33__70_,s_r_33__69_,s_r_33__68_,
  s_r_33__67_,s_r_33__66_,s_r_33__65_,s_r_33__64_,s_r_33__63_,s_r_33__62_,s_r_33__61_,
  s_r_33__60_,s_r_33__59_,s_r_33__58_,s_r_33__57_,s_r_33__56_,s_r_33__55_,s_r_33__54_,
  s_r_33__53_,s_r_33__52_,s_r_33__51_,s_r_33__50_,s_r_33__49_,s_r_33__48_,
  s_r_33__47_,s_r_33__46_,s_r_33__45_,s_r_33__44_,s_r_33__43_,s_r_33__42_,s_r_33__41_,
  s_r_33__40_,s_r_33__39_,s_r_33__38_,s_r_33__37_,s_r_33__36_,s_r_33__35_,s_r_33__34_,
  s_r_33__33_,s_r_33__32_,s_r_33__31_,s_r_33__30_,s_r_33__29_,s_r_33__28_,
  s_r_33__27_,s_r_33__26_,s_r_33__25_,s_r_33__24_,s_r_33__23_,s_r_33__22_,s_r_33__21_,
  s_r_33__20_,s_r_33__19_,s_r_33__18_,s_r_33__17_,s_r_33__16_,s_r_33__15_,s_r_33__14_,
  s_r_33__13_,s_r_33__12_,s_r_33__11_,s_r_33__10_,s_r_33__9_,s_r_33__8_,s_r_33__7_,
  s_r_33__6_,s_r_33__5_,s_r_33__4_,s_r_33__3_,s_r_33__2_,s_r_33__1_,s_r_33__0_,
  s_r_32__127_,s_r_32__126_,s_r_32__125_,s_r_32__124_,s_r_32__123_,s_r_32__122_,
  s_r_32__121_,s_r_32__120_,s_r_32__119_,s_r_32__118_,s_r_32__117_,s_r_32__116_,
  s_r_32__115_,s_r_32__114_,s_r_32__113_,s_r_32__112_,s_r_32__111_,s_r_32__110_,
  s_r_32__109_,s_r_32__108_,s_r_32__107_,s_r_32__106_,s_r_32__105_,s_r_32__104_,
  s_r_32__103_,s_r_32__102_,s_r_32__101_,s_r_32__100_,s_r_32__99_,s_r_32__98_,s_r_32__97_,
  s_r_32__96_,s_r_32__95_,s_r_32__94_,s_r_32__93_,s_r_32__92_,s_r_32__91_,s_r_32__90_,
  s_r_32__89_,s_r_32__88_,s_r_32__87_,s_r_32__86_,s_r_32__85_,s_r_32__84_,
  s_r_32__83_,s_r_32__82_,s_r_32__81_,s_r_32__80_,s_r_32__79_,s_r_32__78_,s_r_32__77_,
  s_r_32__76_,s_r_32__75_,s_r_32__74_,s_r_32__73_,s_r_32__72_,s_r_32__71_,s_r_32__70_,
  s_r_32__69_,s_r_32__68_,s_r_32__67_,s_r_32__66_,s_r_32__65_,s_r_32__64_,
  s_r_32__63_,s_r_32__62_,s_r_32__61_,s_r_32__60_,s_r_32__59_,s_r_32__58_,s_r_32__57_,
  s_r_32__56_,s_r_32__55_,s_r_32__54_,s_r_32__53_,s_r_32__52_,s_r_32__51_,s_r_32__50_,
  s_r_32__49_,s_r_32__48_,s_r_32__47_,s_r_32__46_,s_r_32__45_,s_r_32__44_,
  s_r_32__43_,s_r_32__42_,s_r_32__41_,s_r_32__40_,s_r_32__39_,s_r_32__38_,s_r_32__37_,
  s_r_32__36_,s_r_32__35_,s_r_32__34_,s_r_32__33_,s_r_32__32_,s_r_32__31_,s_r_32__30_,
  s_r_32__29_,s_r_32__28_,s_r_32__27_,s_r_32__26_,s_r_32__25_,s_r_32__24_,
  s_r_32__23_,s_r_32__22_,s_r_32__21_,s_r_32__20_,s_r_32__19_,s_r_32__18_,s_r_32__17_,
  s_r_32__16_,s_r_32__15_,s_r_32__14_,s_r_32__13_,s_r_32__12_,s_r_32__11_,s_r_32__10_,
  s_r_32__9_,s_r_32__8_,s_r_32__7_,s_r_32__6_,s_r_32__5_,s_r_32__4_,s_r_32__3_,
  s_r_32__2_,s_r_32__1_,s_r_32__0_,s_r_31__127_,s_r_31__126_,s_r_31__125_,
  s_r_31__124_,s_r_31__123_,s_r_31__122_,s_r_31__121_,s_r_31__120_,s_r_31__119_,s_r_31__118_,
  s_r_31__117_,s_r_31__116_,s_r_31__115_,s_r_31__114_,s_r_31__113_,s_r_31__112_,
  s_r_31__111_,s_r_31__110_,s_r_31__109_,s_r_31__108_,s_r_31__107_,s_r_31__106_,
  s_r_31__105_,s_r_31__104_,s_r_31__103_,s_r_31__102_,s_r_31__101_,s_r_31__100_,
  s_r_31__99_,s_r_31__98_,s_r_31__97_,s_r_31__96_,s_r_31__95_,s_r_31__94_,s_r_31__93_,
  s_r_31__92_,s_r_31__91_,s_r_31__90_,s_r_31__89_,s_r_31__88_,s_r_31__87_,
  s_r_31__86_,s_r_31__85_,s_r_31__84_,s_r_31__83_,s_r_31__82_,s_r_31__81_,s_r_31__80_,
  s_r_31__79_,s_r_31__78_,s_r_31__77_,s_r_31__76_,s_r_31__75_,s_r_31__74_,s_r_31__73_,
  s_r_31__72_,s_r_31__71_,s_r_31__70_,s_r_31__69_,s_r_31__68_,s_r_31__67_,
  s_r_31__66_,s_r_31__65_,s_r_31__64_,s_r_31__63_,s_r_31__62_,s_r_31__61_,s_r_31__60_,
  s_r_31__59_,s_r_31__58_,s_r_31__57_,s_r_31__56_,s_r_31__55_,s_r_31__54_,s_r_31__53_,
  s_r_31__52_,s_r_31__51_,s_r_31__50_,s_r_31__49_,s_r_31__48_,s_r_31__47_,
  s_r_31__46_,s_r_31__45_,s_r_31__44_,s_r_31__43_,s_r_31__42_,s_r_31__41_,s_r_31__40_,
  s_r_31__39_,s_r_31__38_,s_r_31__37_,s_r_31__36_,s_r_31__35_,s_r_31__34_,s_r_31__33_,
  s_r_31__32_,s_r_31__31_,s_r_31__30_,s_r_31__29_,s_r_31__28_,s_r_31__27_,
  s_r_31__26_,s_r_31__25_,s_r_31__24_,s_r_31__23_,s_r_31__22_,s_r_31__21_,s_r_31__20_,
  s_r_31__19_,s_r_31__18_,s_r_31__17_,s_r_31__16_,s_r_31__15_,s_r_31__14_,s_r_31__13_,
  s_r_31__12_,s_r_31__11_,s_r_31__10_,s_r_31__9_,s_r_31__8_,s_r_31__7_,s_r_31__6_,
  s_r_31__5_,s_r_31__4_,s_r_31__3_,s_r_31__2_,s_r_31__1_,s_r_31__0_,
  prod_accum_34__35_,prod_accum_34__34_,prod_accum_34__33_,prod_accum_34__32_,prod_accum_34__31_,
  prod_accum_34__30_,prod_accum_34__29_,prod_accum_34__28_,prod_accum_34__27_,
  prod_accum_34__26_,prod_accum_34__25_,prod_accum_34__24_,prod_accum_34__23_,
  prod_accum_34__22_,prod_accum_34__21_,prod_accum_34__20_,prod_accum_34__19_,
  prod_accum_34__18_,prod_accum_34__17_,prod_accum_34__16_,prod_accum_34__15_,
  prod_accum_34__14_,prod_accum_34__13_,prod_accum_34__12_,prod_accum_34__11_,prod_accum_34__10_,
  prod_accum_34__9_,prod_accum_34__8_,prod_accum_34__7_,prod_accum_34__6_,
  prod_accum_34__5_,prod_accum_34__4_,prod_accum_34__3_,prod_accum_34__2_,prod_accum_34__1_,
  prod_accum_34__0_,prod_accum_33__34_,prod_accum_33__33_,prod_accum_33__32_,
  prod_accum_33__31_,prod_accum_33__30_,prod_accum_33__29_,prod_accum_33__28_,
  prod_accum_33__27_,prod_accum_33__26_,prod_accum_33__25_,prod_accum_33__24_,
  prod_accum_33__23_,prod_accum_33__22_,prod_accum_33__21_,prod_accum_33__20_,
  prod_accum_33__19_,prod_accum_33__18_,prod_accum_33__17_,prod_accum_33__16_,prod_accum_33__15_,
  prod_accum_33__14_,prod_accum_33__13_,prod_accum_33__12_,prod_accum_33__11_,
  prod_accum_33__10_,prod_accum_33__9_,prod_accum_33__8_,prod_accum_33__7_,
  prod_accum_33__6_,prod_accum_33__5_,prod_accum_33__4_,prod_accum_33__3_,prod_accum_33__2_,
  prod_accum_33__1_,prod_accum_33__0_,prod_accum_32__33_,prod_accum_32__32_,
  prod_accum_32__31_,prod_accum_32__30_,prod_accum_32__29_,prod_accum_32__28_,
  prod_accum_32__27_,prod_accum_32__26_,prod_accum_32__25_,prod_accum_32__24_,
  prod_accum_32__23_,prod_accum_32__22_,prod_accum_32__21_,prod_accum_32__20_,prod_accum_32__19_,
  prod_accum_32__18_,prod_accum_32__17_,prod_accum_32__16_,prod_accum_32__15_,
  prod_accum_32__14_,prod_accum_32__13_,prod_accum_32__12_,prod_accum_32__11_,
  prod_accum_32__10_,prod_accum_32__9_,prod_accum_32__8_,prod_accum_32__7_,
  prod_accum_32__6_,prod_accum_32__5_,prod_accum_32__4_,prod_accum_32__3_,prod_accum_32__2_,
  prod_accum_32__1_,prod_accum_32__0_,prod_accum_31__32_,prod_accum_31__31_,
  prod_accum_31__30_,prod_accum_31__29_,prod_accum_31__28_,prod_accum_31__27_,
  prod_accum_31__26_,prod_accum_31__25_,prod_accum_31__24_,prod_accum_31__23_,prod_accum_31__22_,
  prod_accum_31__21_,prod_accum_31__20_,prod_accum_31__19_,prod_accum_31__18_,
  prod_accum_31__17_,prod_accum_31__16_,prod_accum_31__15_,prod_accum_31__14_,
  prod_accum_31__13_,prod_accum_31__12_,prod_accum_31__11_,prod_accum_31__10_,
  prod_accum_31__9_,prod_accum_31__8_,prod_accum_31__7_,prod_accum_31__6_,prod_accum_31__5_,
  prod_accum_31__4_,prod_accum_31__3_,prod_accum_31__2_,prod_accum_31__1_,
  prod_accum_31__0_,s_r_38__127_,s_r_38__126_,s_r_38__125_,s_r_38__124_,s_r_38__123_,
  s_r_38__122_,s_r_38__121_,s_r_38__120_,s_r_38__119_,s_r_38__118_,s_r_38__117_,
  s_r_38__116_,s_r_38__115_,s_r_38__114_,s_r_38__113_,s_r_38__112_,s_r_38__111_,s_r_38__110_,
  s_r_38__109_,s_r_38__108_,s_r_38__107_,s_r_38__106_,s_r_38__105_,s_r_38__104_,
  s_r_38__103_,s_r_38__102_,s_r_38__101_,s_r_38__100_,s_r_38__99_,s_r_38__98_,
  s_r_38__97_,s_r_38__96_,s_r_38__95_,s_r_38__94_,s_r_38__93_,s_r_38__92_,s_r_38__91_,
  s_r_38__90_,s_r_38__89_,s_r_38__88_,s_r_38__87_,s_r_38__86_,s_r_38__85_,
  s_r_38__84_,s_r_38__83_,s_r_38__82_,s_r_38__81_,s_r_38__80_,s_r_38__79_,s_r_38__78_,
  s_r_38__77_,s_r_38__76_,s_r_38__75_,s_r_38__74_,s_r_38__73_,s_r_38__72_,s_r_38__71_,
  s_r_38__70_,s_r_38__69_,s_r_38__68_,s_r_38__67_,s_r_38__66_,s_r_38__65_,
  s_r_38__64_,s_r_38__63_,s_r_38__62_,s_r_38__61_,s_r_38__60_,s_r_38__59_,s_r_38__58_,
  s_r_38__57_,s_r_38__56_,s_r_38__55_,s_r_38__54_,s_r_38__53_,s_r_38__52_,s_r_38__51_,
  s_r_38__50_,s_r_38__49_,s_r_38__48_,s_r_38__47_,s_r_38__46_,s_r_38__45_,
  s_r_38__44_,s_r_38__43_,s_r_38__42_,s_r_38__41_,s_r_38__40_,s_r_38__39_,s_r_38__38_,
  s_r_38__37_,s_r_38__36_,s_r_38__35_,s_r_38__34_,s_r_38__33_,s_r_38__32_,s_r_38__31_,
  s_r_38__30_,s_r_38__29_,s_r_38__28_,s_r_38__27_,s_r_38__26_,s_r_38__25_,
  s_r_38__24_,s_r_38__23_,s_r_38__22_,s_r_38__21_,s_r_38__20_,s_r_38__19_,s_r_38__18_,
  s_r_38__17_,s_r_38__16_,s_r_38__15_,s_r_38__14_,s_r_38__13_,s_r_38__12_,s_r_38__11_,
  s_r_38__10_,s_r_38__9_,s_r_38__8_,s_r_38__7_,s_r_38__6_,s_r_38__5_,s_r_38__4_,
  s_r_38__3_,s_r_38__2_,s_r_38__1_,s_r_38__0_,s_r_37__127_,s_r_37__126_,s_r_37__125_,
  s_r_37__124_,s_r_37__123_,s_r_37__122_,s_r_37__121_,s_r_37__120_,s_r_37__119_,
  s_r_37__118_,s_r_37__117_,s_r_37__116_,s_r_37__115_,s_r_37__114_,s_r_37__113_,
  s_r_37__112_,s_r_37__111_,s_r_37__110_,s_r_37__109_,s_r_37__108_,s_r_37__107_,
  s_r_37__106_,s_r_37__105_,s_r_37__104_,s_r_37__103_,s_r_37__102_,s_r_37__101_,
  s_r_37__100_,s_r_37__99_,s_r_37__98_,s_r_37__97_,s_r_37__96_,s_r_37__95_,s_r_37__94_,
  s_r_37__93_,s_r_37__92_,s_r_37__91_,s_r_37__90_,s_r_37__89_,s_r_37__88_,s_r_37__87_,
  s_r_37__86_,s_r_37__85_,s_r_37__84_,s_r_37__83_,s_r_37__82_,s_r_37__81_,
  s_r_37__80_,s_r_37__79_,s_r_37__78_,s_r_37__77_,s_r_37__76_,s_r_37__75_,s_r_37__74_,
  s_r_37__73_,s_r_37__72_,s_r_37__71_,s_r_37__70_,s_r_37__69_,s_r_37__68_,s_r_37__67_,
  s_r_37__66_,s_r_37__65_,s_r_37__64_,s_r_37__63_,s_r_37__62_,s_r_37__61_,
  s_r_37__60_,s_r_37__59_,s_r_37__58_,s_r_37__57_,s_r_37__56_,s_r_37__55_,s_r_37__54_,
  s_r_37__53_,s_r_37__52_,s_r_37__51_,s_r_37__50_,s_r_37__49_,s_r_37__48_,s_r_37__47_,
  s_r_37__46_,s_r_37__45_,s_r_37__44_,s_r_37__43_,s_r_37__42_,s_r_37__41_,
  s_r_37__40_,s_r_37__39_,s_r_37__38_,s_r_37__37_,s_r_37__36_,s_r_37__35_,s_r_37__34_,
  s_r_37__33_,s_r_37__32_,s_r_37__31_,s_r_37__30_,s_r_37__29_,s_r_37__28_,s_r_37__27_,
  s_r_37__26_,s_r_37__25_,s_r_37__24_,s_r_37__23_,s_r_37__22_,s_r_37__21_,
  s_r_37__20_,s_r_37__19_,s_r_37__18_,s_r_37__17_,s_r_37__16_,s_r_37__15_,s_r_37__14_,
  s_r_37__13_,s_r_37__12_,s_r_37__11_,s_r_37__10_,s_r_37__9_,s_r_37__8_,s_r_37__7_,
  s_r_37__6_,s_r_37__5_,s_r_37__4_,s_r_37__3_,s_r_37__2_,s_r_37__1_,s_r_37__0_,
  s_r_36__127_,s_r_36__126_,s_r_36__125_,s_r_36__124_,s_r_36__123_,s_r_36__122_,
  s_r_36__121_,s_r_36__120_,s_r_36__119_,s_r_36__118_,s_r_36__117_,s_r_36__116_,
  s_r_36__115_,s_r_36__114_,s_r_36__113_,s_r_36__112_,s_r_36__111_,s_r_36__110_,
  s_r_36__109_,s_r_36__108_,s_r_36__107_,s_r_36__106_,s_r_36__105_,s_r_36__104_,s_r_36__103_,
  s_r_36__102_,s_r_36__101_,s_r_36__100_,s_r_36__99_,s_r_36__98_,s_r_36__97_,
  s_r_36__96_,s_r_36__95_,s_r_36__94_,s_r_36__93_,s_r_36__92_,s_r_36__91_,s_r_36__90_,
  s_r_36__89_,s_r_36__88_,s_r_36__87_,s_r_36__86_,s_r_36__85_,s_r_36__84_,
  s_r_36__83_,s_r_36__82_,s_r_36__81_,s_r_36__80_,s_r_36__79_,s_r_36__78_,s_r_36__77_,
  s_r_36__76_,s_r_36__75_,s_r_36__74_,s_r_36__73_,s_r_36__72_,s_r_36__71_,s_r_36__70_,
  s_r_36__69_,s_r_36__68_,s_r_36__67_,s_r_36__66_,s_r_36__65_,s_r_36__64_,
  s_r_36__63_,s_r_36__62_,s_r_36__61_,s_r_36__60_,s_r_36__59_,s_r_36__58_,s_r_36__57_,
  s_r_36__56_,s_r_36__55_,s_r_36__54_,s_r_36__53_,s_r_36__52_,s_r_36__51_,s_r_36__50_,
  s_r_36__49_,s_r_36__48_,s_r_36__47_,s_r_36__46_,s_r_36__45_,s_r_36__44_,
  s_r_36__43_,s_r_36__42_,s_r_36__41_,s_r_36__40_,s_r_36__39_,s_r_36__38_,s_r_36__37_,
  s_r_36__36_,s_r_36__35_,s_r_36__34_,s_r_36__33_,s_r_36__32_,s_r_36__31_,s_r_36__30_,
  s_r_36__29_,s_r_36__28_,s_r_36__27_,s_r_36__26_,s_r_36__25_,s_r_36__24_,
  s_r_36__23_,s_r_36__22_,s_r_36__21_,s_r_36__20_,s_r_36__19_,s_r_36__18_,s_r_36__17_,
  s_r_36__16_,s_r_36__15_,s_r_36__14_,s_r_36__13_,s_r_36__12_,s_r_36__11_,s_r_36__10_,
  s_r_36__9_,s_r_36__8_,s_r_36__7_,s_r_36__6_,s_r_36__5_,s_r_36__4_,s_r_36__3_,
  s_r_36__2_,s_r_36__1_,s_r_36__0_,s_r_35__127_,s_r_35__126_,s_r_35__125_,s_r_35__124_,
  s_r_35__123_,s_r_35__122_,s_r_35__121_,s_r_35__120_,s_r_35__119_,s_r_35__118_,
  s_r_35__117_,s_r_35__116_,s_r_35__115_,s_r_35__114_,s_r_35__113_,s_r_35__112_,
  s_r_35__111_,s_r_35__110_,s_r_35__109_,s_r_35__108_,s_r_35__107_,s_r_35__106_,
  s_r_35__105_,s_r_35__104_,s_r_35__103_,s_r_35__102_,s_r_35__101_,s_r_35__100_,
  s_r_35__99_,s_r_35__98_,s_r_35__97_,s_r_35__96_,s_r_35__95_,s_r_35__94_,s_r_35__93_,
  s_r_35__92_,s_r_35__91_,s_r_35__90_,s_r_35__89_,s_r_35__88_,s_r_35__87_,s_r_35__86_,
  s_r_35__85_,s_r_35__84_,s_r_35__83_,s_r_35__82_,s_r_35__81_,s_r_35__80_,
  s_r_35__79_,s_r_35__78_,s_r_35__77_,s_r_35__76_,s_r_35__75_,s_r_35__74_,s_r_35__73_,
  s_r_35__72_,s_r_35__71_,s_r_35__70_,s_r_35__69_,s_r_35__68_,s_r_35__67_,s_r_35__66_,
  s_r_35__65_,s_r_35__64_,s_r_35__63_,s_r_35__62_,s_r_35__61_,s_r_35__60_,
  s_r_35__59_,s_r_35__58_,s_r_35__57_,s_r_35__56_,s_r_35__55_,s_r_35__54_,s_r_35__53_,
  s_r_35__52_,s_r_35__51_,s_r_35__50_,s_r_35__49_,s_r_35__48_,s_r_35__47_,s_r_35__46_,
  s_r_35__45_,s_r_35__44_,s_r_35__43_,s_r_35__42_,s_r_35__41_,s_r_35__40_,
  s_r_35__39_,s_r_35__38_,s_r_35__37_,s_r_35__36_,s_r_35__35_,s_r_35__34_,s_r_35__33_,
  s_r_35__32_,s_r_35__31_,s_r_35__30_,s_r_35__29_,s_r_35__28_,s_r_35__27_,s_r_35__26_,
  s_r_35__25_,s_r_35__24_,s_r_35__23_,s_r_35__22_,s_r_35__21_,s_r_35__20_,
  s_r_35__19_,s_r_35__18_,s_r_35__17_,s_r_35__16_,s_r_35__15_,s_r_35__14_,s_r_35__13_,
  s_r_35__12_,s_r_35__11_,s_r_35__10_,s_r_35__9_,s_r_35__8_,s_r_35__7_,s_r_35__6_,
  s_r_35__5_,s_r_35__4_,s_r_35__3_,s_r_35__2_,s_r_35__1_,s_r_35__0_,
  prod_accum_38__39_,prod_accum_38__38_,prod_accum_38__37_,prod_accum_38__36_,prod_accum_38__35_,
  prod_accum_38__34_,prod_accum_38__33_,prod_accum_38__32_,prod_accum_38__31_,
  prod_accum_38__30_,prod_accum_38__29_,prod_accum_38__28_,prod_accum_38__27_,
  prod_accum_38__26_,prod_accum_38__25_,prod_accum_38__24_,prod_accum_38__23_,
  prod_accum_38__22_,prod_accum_38__21_,prod_accum_38__20_,prod_accum_38__19_,prod_accum_38__18_,
  prod_accum_38__17_,prod_accum_38__16_,prod_accum_38__15_,prod_accum_38__14_,
  prod_accum_38__13_,prod_accum_38__12_,prod_accum_38__11_,prod_accum_38__10_,
  prod_accum_38__9_,prod_accum_38__8_,prod_accum_38__7_,prod_accum_38__6_,
  prod_accum_38__5_,prod_accum_38__4_,prod_accum_38__3_,prod_accum_38__2_,prod_accum_38__1_,
  prod_accum_38__0_,prod_accum_37__38_,prod_accum_37__37_,prod_accum_37__36_,
  prod_accum_37__35_,prod_accum_37__34_,prod_accum_37__33_,prod_accum_37__32_,
  prod_accum_37__31_,prod_accum_37__30_,prod_accum_37__29_,prod_accum_37__28_,prod_accum_37__27_,
  prod_accum_37__26_,prod_accum_37__25_,prod_accum_37__24_,prod_accum_37__23_,
  prod_accum_37__22_,prod_accum_37__21_,prod_accum_37__20_,prod_accum_37__19_,
  prod_accum_37__18_,prod_accum_37__17_,prod_accum_37__16_,prod_accum_37__15_,
  prod_accum_37__14_,prod_accum_37__13_,prod_accum_37__12_,prod_accum_37__11_,
  prod_accum_37__10_,prod_accum_37__9_,prod_accum_37__8_,prod_accum_37__7_,prod_accum_37__6_,
  prod_accum_37__5_,prod_accum_37__4_,prod_accum_37__3_,prod_accum_37__2_,
  prod_accum_37__1_,prod_accum_37__0_,prod_accum_36__37_,prod_accum_36__36_,prod_accum_36__35_,
  prod_accum_36__34_,prod_accum_36__33_,prod_accum_36__32_,prod_accum_36__31_,
  prod_accum_36__30_,prod_accum_36__29_,prod_accum_36__28_,prod_accum_36__27_,
  prod_accum_36__26_,prod_accum_36__25_,prod_accum_36__24_,prod_accum_36__23_,
  prod_accum_36__22_,prod_accum_36__21_,prod_accum_36__20_,prod_accum_36__19_,
  prod_accum_36__18_,prod_accum_36__17_,prod_accum_36__16_,prod_accum_36__15_,prod_accum_36__14_,
  prod_accum_36__13_,prod_accum_36__12_,prod_accum_36__11_,prod_accum_36__10_,
  prod_accum_36__9_,prod_accum_36__8_,prod_accum_36__7_,prod_accum_36__6_,
  prod_accum_36__5_,prod_accum_36__4_,prod_accum_36__3_,prod_accum_36__2_,prod_accum_36__1_,
  prod_accum_36__0_,prod_accum_35__36_,prod_accum_35__35_,prod_accum_35__34_,
  prod_accum_35__33_,prod_accum_35__32_,prod_accum_35__31_,prod_accum_35__30_,
  prod_accum_35__29_,prod_accum_35__28_,prod_accum_35__27_,prod_accum_35__26_,
  prod_accum_35__25_,prod_accum_35__24_,prod_accum_35__23_,prod_accum_35__22_,prod_accum_35__21_,
  prod_accum_35__20_,prod_accum_35__19_,prod_accum_35__18_,prod_accum_35__17_,
  prod_accum_35__16_,prod_accum_35__15_,prod_accum_35__14_,prod_accum_35__13_,
  prod_accum_35__12_,prod_accum_35__11_,prod_accum_35__10_,prod_accum_35__9_,
  prod_accum_35__8_,prod_accum_35__7_,prod_accum_35__6_,prod_accum_35__5_,prod_accum_35__4_,
  prod_accum_35__3_,prod_accum_35__2_,prod_accum_35__1_,prod_accum_35__0_,
  s_r_42__127_,s_r_42__126_,s_r_42__125_,s_r_42__124_,s_r_42__123_,s_r_42__122_,s_r_42__121_,
  s_r_42__120_,s_r_42__119_,s_r_42__118_,s_r_42__117_,s_r_42__116_,s_r_42__115_,
  s_r_42__114_,s_r_42__113_,s_r_42__112_,s_r_42__111_,s_r_42__110_,s_r_42__109_,
  s_r_42__108_,s_r_42__107_,s_r_42__106_,s_r_42__105_,s_r_42__104_,s_r_42__103_,
  s_r_42__102_,s_r_42__101_,s_r_42__100_,s_r_42__99_,s_r_42__98_,s_r_42__97_,s_r_42__96_,
  s_r_42__95_,s_r_42__94_,s_r_42__93_,s_r_42__92_,s_r_42__91_,s_r_42__90_,
  s_r_42__89_,s_r_42__88_,s_r_42__87_,s_r_42__86_,s_r_42__85_,s_r_42__84_,s_r_42__83_,
  s_r_42__82_,s_r_42__81_,s_r_42__80_,s_r_42__79_,s_r_42__78_,s_r_42__77_,s_r_42__76_,
  s_r_42__75_,s_r_42__74_,s_r_42__73_,s_r_42__72_,s_r_42__71_,s_r_42__70_,
  s_r_42__69_,s_r_42__68_,s_r_42__67_,s_r_42__66_,s_r_42__65_,s_r_42__64_,s_r_42__63_,
  s_r_42__62_,s_r_42__61_,s_r_42__60_,s_r_42__59_,s_r_42__58_,s_r_42__57_,s_r_42__56_,
  s_r_42__55_,s_r_42__54_,s_r_42__53_,s_r_42__52_,s_r_42__51_,s_r_42__50_,
  s_r_42__49_,s_r_42__48_,s_r_42__47_,s_r_42__46_,s_r_42__45_,s_r_42__44_,s_r_42__43_,
  s_r_42__42_,s_r_42__41_,s_r_42__40_,s_r_42__39_,s_r_42__38_,s_r_42__37_,s_r_42__36_,
  s_r_42__35_,s_r_42__34_,s_r_42__33_,s_r_42__32_,s_r_42__31_,s_r_42__30_,
  s_r_42__29_,s_r_42__28_,s_r_42__27_,s_r_42__26_,s_r_42__25_,s_r_42__24_,s_r_42__23_,
  s_r_42__22_,s_r_42__21_,s_r_42__20_,s_r_42__19_,s_r_42__18_,s_r_42__17_,s_r_42__16_,
  s_r_42__15_,s_r_42__14_,s_r_42__13_,s_r_42__12_,s_r_42__11_,s_r_42__10_,
  s_r_42__9_,s_r_42__8_,s_r_42__7_,s_r_42__6_,s_r_42__5_,s_r_42__4_,s_r_42__3_,s_r_42__2_,
  s_r_42__1_,s_r_42__0_,s_r_41__127_,s_r_41__126_,s_r_41__125_,s_r_41__124_,
  s_r_41__123_,s_r_41__122_,s_r_41__121_,s_r_41__120_,s_r_41__119_,s_r_41__118_,
  s_r_41__117_,s_r_41__116_,s_r_41__115_,s_r_41__114_,s_r_41__113_,s_r_41__112_,
  s_r_41__111_,s_r_41__110_,s_r_41__109_,s_r_41__108_,s_r_41__107_,s_r_41__106_,
  s_r_41__105_,s_r_41__104_,s_r_41__103_,s_r_41__102_,s_r_41__101_,s_r_41__100_,s_r_41__99_,
  s_r_41__98_,s_r_41__97_,s_r_41__96_,s_r_41__95_,s_r_41__94_,s_r_41__93_,
  s_r_41__92_,s_r_41__91_,s_r_41__90_,s_r_41__89_,s_r_41__88_,s_r_41__87_,s_r_41__86_,
  s_r_41__85_,s_r_41__84_,s_r_41__83_,s_r_41__82_,s_r_41__81_,s_r_41__80_,s_r_41__79_,
  s_r_41__78_,s_r_41__77_,s_r_41__76_,s_r_41__75_,s_r_41__74_,s_r_41__73_,
  s_r_41__72_,s_r_41__71_,s_r_41__70_,s_r_41__69_,s_r_41__68_,s_r_41__67_,s_r_41__66_,
  s_r_41__65_,s_r_41__64_,s_r_41__63_,s_r_41__62_,s_r_41__61_,s_r_41__60_,s_r_41__59_,
  s_r_41__58_,s_r_41__57_,s_r_41__56_,s_r_41__55_,s_r_41__54_,s_r_41__53_,
  s_r_41__52_,s_r_41__51_,s_r_41__50_,s_r_41__49_,s_r_41__48_,s_r_41__47_,s_r_41__46_,
  s_r_41__45_,s_r_41__44_,s_r_41__43_,s_r_41__42_,s_r_41__41_,s_r_41__40_,s_r_41__39_,
  s_r_41__38_,s_r_41__37_,s_r_41__36_,s_r_41__35_,s_r_41__34_,s_r_41__33_,
  s_r_41__32_,s_r_41__31_,s_r_41__30_,s_r_41__29_,s_r_41__28_,s_r_41__27_,s_r_41__26_,
  s_r_41__25_,s_r_41__24_,s_r_41__23_,s_r_41__22_,s_r_41__21_,s_r_41__20_,s_r_41__19_,
  s_r_41__18_,s_r_41__17_,s_r_41__16_,s_r_41__15_,s_r_41__14_,s_r_41__13_,
  s_r_41__12_,s_r_41__11_,s_r_41__10_,s_r_41__9_,s_r_41__8_,s_r_41__7_,s_r_41__6_,
  s_r_41__5_,s_r_41__4_,s_r_41__3_,s_r_41__2_,s_r_41__1_,s_r_41__0_,s_r_40__127_,
  s_r_40__126_,s_r_40__125_,s_r_40__124_,s_r_40__123_,s_r_40__122_,s_r_40__121_,s_r_40__120_,
  s_r_40__119_,s_r_40__118_,s_r_40__117_,s_r_40__116_,s_r_40__115_,s_r_40__114_,
  s_r_40__113_,s_r_40__112_,s_r_40__111_,s_r_40__110_,s_r_40__109_,s_r_40__108_,
  s_r_40__107_,s_r_40__106_,s_r_40__105_,s_r_40__104_,s_r_40__103_,s_r_40__102_,
  s_r_40__101_,s_r_40__100_,s_r_40__99_,s_r_40__98_,s_r_40__97_,s_r_40__96_,s_r_40__95_,
  s_r_40__94_,s_r_40__93_,s_r_40__92_,s_r_40__91_,s_r_40__90_,s_r_40__89_,
  s_r_40__88_,s_r_40__87_,s_r_40__86_,s_r_40__85_,s_r_40__84_,s_r_40__83_,s_r_40__82_,
  s_r_40__81_,s_r_40__80_,s_r_40__79_,s_r_40__78_,s_r_40__77_,s_r_40__76_,s_r_40__75_,
  s_r_40__74_,s_r_40__73_,s_r_40__72_,s_r_40__71_,s_r_40__70_,s_r_40__69_,
  s_r_40__68_,s_r_40__67_,s_r_40__66_,s_r_40__65_,s_r_40__64_,s_r_40__63_,s_r_40__62_,
  s_r_40__61_,s_r_40__60_,s_r_40__59_,s_r_40__58_,s_r_40__57_,s_r_40__56_,s_r_40__55_,
  s_r_40__54_,s_r_40__53_,s_r_40__52_,s_r_40__51_,s_r_40__50_,s_r_40__49_,
  s_r_40__48_,s_r_40__47_,s_r_40__46_,s_r_40__45_,s_r_40__44_,s_r_40__43_,s_r_40__42_,
  s_r_40__41_,s_r_40__40_,s_r_40__39_,s_r_40__38_,s_r_40__37_,s_r_40__36_,s_r_40__35_,
  s_r_40__34_,s_r_40__33_,s_r_40__32_,s_r_40__31_,s_r_40__30_,s_r_40__29_,
  s_r_40__28_,s_r_40__27_,s_r_40__26_,s_r_40__25_,s_r_40__24_,s_r_40__23_,s_r_40__22_,
  s_r_40__21_,s_r_40__20_,s_r_40__19_,s_r_40__18_,s_r_40__17_,s_r_40__16_,s_r_40__15_,
  s_r_40__14_,s_r_40__13_,s_r_40__12_,s_r_40__11_,s_r_40__10_,s_r_40__9_,
  s_r_40__8_,s_r_40__7_,s_r_40__6_,s_r_40__5_,s_r_40__4_,s_r_40__3_,s_r_40__2_,s_r_40__1_,
  s_r_40__0_,s_r_39__127_,s_r_39__126_,s_r_39__125_,s_r_39__124_,s_r_39__123_,
  s_r_39__122_,s_r_39__121_,s_r_39__120_,s_r_39__119_,s_r_39__118_,s_r_39__117_,
  s_r_39__116_,s_r_39__115_,s_r_39__114_,s_r_39__113_,s_r_39__112_,s_r_39__111_,
  s_r_39__110_,s_r_39__109_,s_r_39__108_,s_r_39__107_,s_r_39__106_,s_r_39__105_,
  s_r_39__104_,s_r_39__103_,s_r_39__102_,s_r_39__101_,s_r_39__100_,s_r_39__99_,s_r_39__98_,
  s_r_39__97_,s_r_39__96_,s_r_39__95_,s_r_39__94_,s_r_39__93_,s_r_39__92_,
  s_r_39__91_,s_r_39__90_,s_r_39__89_,s_r_39__88_,s_r_39__87_,s_r_39__86_,s_r_39__85_,
  s_r_39__84_,s_r_39__83_,s_r_39__82_,s_r_39__81_,s_r_39__80_,s_r_39__79_,s_r_39__78_,
  s_r_39__77_,s_r_39__76_,s_r_39__75_,s_r_39__74_,s_r_39__73_,s_r_39__72_,
  s_r_39__71_,s_r_39__70_,s_r_39__69_,s_r_39__68_,s_r_39__67_,s_r_39__66_,s_r_39__65_,
  s_r_39__64_,s_r_39__63_,s_r_39__62_,s_r_39__61_,s_r_39__60_,s_r_39__59_,s_r_39__58_,
  s_r_39__57_,s_r_39__56_,s_r_39__55_,s_r_39__54_,s_r_39__53_,s_r_39__52_,
  s_r_39__51_,s_r_39__50_,s_r_39__49_,s_r_39__48_,s_r_39__47_,s_r_39__46_,s_r_39__45_,
  s_r_39__44_,s_r_39__43_,s_r_39__42_,s_r_39__41_,s_r_39__40_,s_r_39__39_,s_r_39__38_,
  s_r_39__37_,s_r_39__36_,s_r_39__35_,s_r_39__34_,s_r_39__33_,s_r_39__32_,
  s_r_39__31_,s_r_39__30_,s_r_39__29_,s_r_39__28_,s_r_39__27_,s_r_39__26_,s_r_39__25_,
  s_r_39__24_,s_r_39__23_,s_r_39__22_,s_r_39__21_,s_r_39__20_,s_r_39__19_,s_r_39__18_,
  s_r_39__17_,s_r_39__16_,s_r_39__15_,s_r_39__14_,s_r_39__13_,s_r_39__12_,
  s_r_39__11_,s_r_39__10_,s_r_39__9_,s_r_39__8_,s_r_39__7_,s_r_39__6_,s_r_39__5_,s_r_39__4_,
  s_r_39__3_,s_r_39__2_,s_r_39__1_,s_r_39__0_,prod_accum_42__43_,
  prod_accum_42__42_,prod_accum_42__41_,prod_accum_42__40_,prod_accum_42__39_,prod_accum_42__38_,
  prod_accum_42__37_,prod_accum_42__36_,prod_accum_42__35_,prod_accum_42__34_,
  prod_accum_42__33_,prod_accum_42__32_,prod_accum_42__31_,prod_accum_42__30_,
  prod_accum_42__29_,prod_accum_42__28_,prod_accum_42__27_,prod_accum_42__26_,
  prod_accum_42__25_,prod_accum_42__24_,prod_accum_42__23_,prod_accum_42__22_,
  prod_accum_42__21_,prod_accum_42__20_,prod_accum_42__19_,prod_accum_42__18_,prod_accum_42__17_,
  prod_accum_42__16_,prod_accum_42__15_,prod_accum_42__14_,prod_accum_42__13_,
  prod_accum_42__12_,prod_accum_42__11_,prod_accum_42__10_,prod_accum_42__9_,
  prod_accum_42__8_,prod_accum_42__7_,prod_accum_42__6_,prod_accum_42__5_,prod_accum_42__4_,
  prod_accum_42__3_,prod_accum_42__2_,prod_accum_42__1_,prod_accum_42__0_,
  prod_accum_41__42_,prod_accum_41__41_,prod_accum_41__40_,prod_accum_41__39_,
  prod_accum_41__38_,prod_accum_41__37_,prod_accum_41__36_,prod_accum_41__35_,
  prod_accum_41__34_,prod_accum_41__33_,prod_accum_41__32_,prod_accum_41__31_,prod_accum_41__30_,
  prod_accum_41__29_,prod_accum_41__28_,prod_accum_41__27_,prod_accum_41__26_,
  prod_accum_41__25_,prod_accum_41__24_,prod_accum_41__23_,prod_accum_41__22_,
  prod_accum_41__21_,prod_accum_41__20_,prod_accum_41__19_,prod_accum_41__18_,
  prod_accum_41__17_,prod_accum_41__16_,prod_accum_41__15_,prod_accum_41__14_,prod_accum_41__13_,
  prod_accum_41__12_,prod_accum_41__11_,prod_accum_41__10_,prod_accum_41__9_,
  prod_accum_41__8_,prod_accum_41__7_,prod_accum_41__6_,prod_accum_41__5_,
  prod_accum_41__4_,prod_accum_41__3_,prod_accum_41__2_,prod_accum_41__1_,prod_accum_41__0_,
  prod_accum_40__41_,prod_accum_40__40_,prod_accum_40__39_,prod_accum_40__38_,
  prod_accum_40__37_,prod_accum_40__36_,prod_accum_40__35_,prod_accum_40__34_,
  prod_accum_40__33_,prod_accum_40__32_,prod_accum_40__31_,prod_accum_40__30_,
  prod_accum_40__29_,prod_accum_40__28_,prod_accum_40__27_,prod_accum_40__26_,prod_accum_40__25_,
  prod_accum_40__24_,prod_accum_40__23_,prod_accum_40__22_,prod_accum_40__21_,
  prod_accum_40__20_,prod_accum_40__19_,prod_accum_40__18_,prod_accum_40__17_,
  prod_accum_40__16_,prod_accum_40__15_,prod_accum_40__14_,prod_accum_40__13_,
  prod_accum_40__12_,prod_accum_40__11_,prod_accum_40__10_,prod_accum_40__9_,
  prod_accum_40__8_,prod_accum_40__7_,prod_accum_40__6_,prod_accum_40__5_,prod_accum_40__4_,
  prod_accum_40__3_,prod_accum_40__2_,prod_accum_40__1_,prod_accum_40__0_,
  prod_accum_39__40_,prod_accum_39__39_,prod_accum_39__38_,prod_accum_39__37_,prod_accum_39__36_,
  prod_accum_39__35_,prod_accum_39__34_,prod_accum_39__33_,prod_accum_39__32_,
  prod_accum_39__31_,prod_accum_39__30_,prod_accum_39__29_,prod_accum_39__28_,
  prod_accum_39__27_,prod_accum_39__26_,prod_accum_39__25_,prod_accum_39__24_,
  prod_accum_39__23_,prod_accum_39__22_,prod_accum_39__21_,prod_accum_39__20_,
  prod_accum_39__19_,prod_accum_39__18_,prod_accum_39__17_,prod_accum_39__16_,prod_accum_39__15_,
  prod_accum_39__14_,prod_accum_39__13_,prod_accum_39__12_,prod_accum_39__11_,
  prod_accum_39__10_,prod_accum_39__9_,prod_accum_39__8_,prod_accum_39__7_,
  prod_accum_39__6_,prod_accum_39__5_,prod_accum_39__4_,prod_accum_39__3_,prod_accum_39__2_,
  prod_accum_39__1_,prod_accum_39__0_,s_r_46__127_,s_r_46__126_,s_r_46__125_,
  s_r_46__124_,s_r_46__123_,s_r_46__122_,s_r_46__121_,s_r_46__120_,s_r_46__119_,
  s_r_46__118_,s_r_46__117_,s_r_46__116_,s_r_46__115_,s_r_46__114_,s_r_46__113_,
  s_r_46__112_,s_r_46__111_,s_r_46__110_,s_r_46__109_,s_r_46__108_,s_r_46__107_,s_r_46__106_,
  s_r_46__105_,s_r_46__104_,s_r_46__103_,s_r_46__102_,s_r_46__101_,s_r_46__100_,
  s_r_46__99_,s_r_46__98_,s_r_46__97_,s_r_46__96_,s_r_46__95_,s_r_46__94_,
  s_r_46__93_,s_r_46__92_,s_r_46__91_,s_r_46__90_,s_r_46__89_,s_r_46__88_,s_r_46__87_,
  s_r_46__86_,s_r_46__85_,s_r_46__84_,s_r_46__83_,s_r_46__82_,s_r_46__81_,s_r_46__80_,
  s_r_46__79_,s_r_46__78_,s_r_46__77_,s_r_46__76_,s_r_46__75_,s_r_46__74_,
  s_r_46__73_,s_r_46__72_,s_r_46__71_,s_r_46__70_,s_r_46__69_,s_r_46__68_,s_r_46__67_,
  s_r_46__66_,s_r_46__65_,s_r_46__64_,s_r_46__63_,s_r_46__62_,s_r_46__61_,s_r_46__60_,
  s_r_46__59_,s_r_46__58_,s_r_46__57_,s_r_46__56_,s_r_46__55_,s_r_46__54_,
  s_r_46__53_,s_r_46__52_,s_r_46__51_,s_r_46__50_,s_r_46__49_,s_r_46__48_,s_r_46__47_,
  s_r_46__46_,s_r_46__45_,s_r_46__44_,s_r_46__43_,s_r_46__42_,s_r_46__41_,s_r_46__40_,
  s_r_46__39_,s_r_46__38_,s_r_46__37_,s_r_46__36_,s_r_46__35_,s_r_46__34_,
  s_r_46__33_,s_r_46__32_,s_r_46__31_,s_r_46__30_,s_r_46__29_,s_r_46__28_,s_r_46__27_,
  s_r_46__26_,s_r_46__25_,s_r_46__24_,s_r_46__23_,s_r_46__22_,s_r_46__21_,s_r_46__20_,
  s_r_46__19_,s_r_46__18_,s_r_46__17_,s_r_46__16_,s_r_46__15_,s_r_46__14_,
  s_r_46__13_,s_r_46__12_,s_r_46__11_,s_r_46__10_,s_r_46__9_,s_r_46__8_,s_r_46__7_,
  s_r_46__6_,s_r_46__5_,s_r_46__4_,s_r_46__3_,s_r_46__2_,s_r_46__1_,s_r_46__0_,
  s_r_45__127_,s_r_45__126_,s_r_45__125_,s_r_45__124_,s_r_45__123_,s_r_45__122_,s_r_45__121_,
  s_r_45__120_,s_r_45__119_,s_r_45__118_,s_r_45__117_,s_r_45__116_,s_r_45__115_,
  s_r_45__114_,s_r_45__113_,s_r_45__112_,s_r_45__111_,s_r_45__110_,s_r_45__109_,
  s_r_45__108_,s_r_45__107_,s_r_45__106_,s_r_45__105_,s_r_45__104_,s_r_45__103_,
  s_r_45__102_,s_r_45__101_,s_r_45__100_,s_r_45__99_,s_r_45__98_,s_r_45__97_,s_r_45__96_,
  s_r_45__95_,s_r_45__94_,s_r_45__93_,s_r_45__92_,s_r_45__91_,s_r_45__90_,
  s_r_45__89_,s_r_45__88_,s_r_45__87_,s_r_45__86_,s_r_45__85_,s_r_45__84_,s_r_45__83_,
  s_r_45__82_,s_r_45__81_,s_r_45__80_,s_r_45__79_,s_r_45__78_,s_r_45__77_,s_r_45__76_,
  s_r_45__75_,s_r_45__74_,s_r_45__73_,s_r_45__72_,s_r_45__71_,s_r_45__70_,
  s_r_45__69_,s_r_45__68_,s_r_45__67_,s_r_45__66_,s_r_45__65_,s_r_45__64_,s_r_45__63_,
  s_r_45__62_,s_r_45__61_,s_r_45__60_,s_r_45__59_,s_r_45__58_,s_r_45__57_,s_r_45__56_,
  s_r_45__55_,s_r_45__54_,s_r_45__53_,s_r_45__52_,s_r_45__51_,s_r_45__50_,
  s_r_45__49_,s_r_45__48_,s_r_45__47_,s_r_45__46_,s_r_45__45_,s_r_45__44_,s_r_45__43_,
  s_r_45__42_,s_r_45__41_,s_r_45__40_,s_r_45__39_,s_r_45__38_,s_r_45__37_,s_r_45__36_,
  s_r_45__35_,s_r_45__34_,s_r_45__33_,s_r_45__32_,s_r_45__31_,s_r_45__30_,
  s_r_45__29_,s_r_45__28_,s_r_45__27_,s_r_45__26_,s_r_45__25_,s_r_45__24_,s_r_45__23_,
  s_r_45__22_,s_r_45__21_,s_r_45__20_,s_r_45__19_,s_r_45__18_,s_r_45__17_,s_r_45__16_,
  s_r_45__15_,s_r_45__14_,s_r_45__13_,s_r_45__12_,s_r_45__11_,s_r_45__10_,
  s_r_45__9_,s_r_45__8_,s_r_45__7_,s_r_45__6_,s_r_45__5_,s_r_45__4_,s_r_45__3_,s_r_45__2_,
  s_r_45__1_,s_r_45__0_,s_r_44__127_,s_r_44__126_,s_r_44__125_,s_r_44__124_,
  s_r_44__123_,s_r_44__122_,s_r_44__121_,s_r_44__120_,s_r_44__119_,s_r_44__118_,
  s_r_44__117_,s_r_44__116_,s_r_44__115_,s_r_44__114_,s_r_44__113_,s_r_44__112_,
  s_r_44__111_,s_r_44__110_,s_r_44__109_,s_r_44__108_,s_r_44__107_,s_r_44__106_,
  s_r_44__105_,s_r_44__104_,s_r_44__103_,s_r_44__102_,s_r_44__101_,s_r_44__100_,s_r_44__99_,
  s_r_44__98_,s_r_44__97_,s_r_44__96_,s_r_44__95_,s_r_44__94_,s_r_44__93_,
  s_r_44__92_,s_r_44__91_,s_r_44__90_,s_r_44__89_,s_r_44__88_,s_r_44__87_,s_r_44__86_,
  s_r_44__85_,s_r_44__84_,s_r_44__83_,s_r_44__82_,s_r_44__81_,s_r_44__80_,s_r_44__79_,
  s_r_44__78_,s_r_44__77_,s_r_44__76_,s_r_44__75_,s_r_44__74_,s_r_44__73_,
  s_r_44__72_,s_r_44__71_,s_r_44__70_,s_r_44__69_,s_r_44__68_,s_r_44__67_,s_r_44__66_,
  s_r_44__65_,s_r_44__64_,s_r_44__63_,s_r_44__62_,s_r_44__61_,s_r_44__60_,s_r_44__59_,
  s_r_44__58_,s_r_44__57_,s_r_44__56_,s_r_44__55_,s_r_44__54_,s_r_44__53_,
  s_r_44__52_,s_r_44__51_,s_r_44__50_,s_r_44__49_,s_r_44__48_,s_r_44__47_,s_r_44__46_,
  s_r_44__45_,s_r_44__44_,s_r_44__43_,s_r_44__42_,s_r_44__41_,s_r_44__40_,s_r_44__39_,
  s_r_44__38_,s_r_44__37_,s_r_44__36_,s_r_44__35_,s_r_44__34_,s_r_44__33_,
  s_r_44__32_,s_r_44__31_,s_r_44__30_,s_r_44__29_,s_r_44__28_,s_r_44__27_,s_r_44__26_,
  s_r_44__25_,s_r_44__24_,s_r_44__23_,s_r_44__22_,s_r_44__21_,s_r_44__20_,s_r_44__19_,
  s_r_44__18_,s_r_44__17_,s_r_44__16_,s_r_44__15_,s_r_44__14_,s_r_44__13_,
  s_r_44__12_,s_r_44__11_,s_r_44__10_,s_r_44__9_,s_r_44__8_,s_r_44__7_,s_r_44__6_,
  s_r_44__5_,s_r_44__4_,s_r_44__3_,s_r_44__2_,s_r_44__1_,s_r_44__0_,s_r_43__127_,
  s_r_43__126_,s_r_43__125_,s_r_43__124_,s_r_43__123_,s_r_43__122_,s_r_43__121_,s_r_43__120_,
  s_r_43__119_,s_r_43__118_,s_r_43__117_,s_r_43__116_,s_r_43__115_,s_r_43__114_,
  s_r_43__113_,s_r_43__112_,s_r_43__111_,s_r_43__110_,s_r_43__109_,s_r_43__108_,
  s_r_43__107_,s_r_43__106_,s_r_43__105_,s_r_43__104_,s_r_43__103_,s_r_43__102_,
  s_r_43__101_,s_r_43__100_,s_r_43__99_,s_r_43__98_,s_r_43__97_,s_r_43__96_,s_r_43__95_,
  s_r_43__94_,s_r_43__93_,s_r_43__92_,s_r_43__91_,s_r_43__90_,s_r_43__89_,
  s_r_43__88_,s_r_43__87_,s_r_43__86_,s_r_43__85_,s_r_43__84_,s_r_43__83_,s_r_43__82_,
  s_r_43__81_,s_r_43__80_,s_r_43__79_,s_r_43__78_,s_r_43__77_,s_r_43__76_,s_r_43__75_,
  s_r_43__74_,s_r_43__73_,s_r_43__72_,s_r_43__71_,s_r_43__70_,s_r_43__69_,
  s_r_43__68_,s_r_43__67_,s_r_43__66_,s_r_43__65_,s_r_43__64_,s_r_43__63_,s_r_43__62_,
  s_r_43__61_,s_r_43__60_,s_r_43__59_,s_r_43__58_,s_r_43__57_,s_r_43__56_,s_r_43__55_,
  s_r_43__54_,s_r_43__53_,s_r_43__52_,s_r_43__51_,s_r_43__50_,s_r_43__49_,
  s_r_43__48_,s_r_43__47_,s_r_43__46_,s_r_43__45_,s_r_43__44_,s_r_43__43_,s_r_43__42_,
  s_r_43__41_,s_r_43__40_,s_r_43__39_,s_r_43__38_,s_r_43__37_,s_r_43__36_,s_r_43__35_,
  s_r_43__34_,s_r_43__33_,s_r_43__32_,s_r_43__31_,s_r_43__30_,s_r_43__29_,
  s_r_43__28_,s_r_43__27_,s_r_43__26_,s_r_43__25_,s_r_43__24_,s_r_43__23_,s_r_43__22_,
  s_r_43__21_,s_r_43__20_,s_r_43__19_,s_r_43__18_,s_r_43__17_,s_r_43__16_,s_r_43__15_,
  s_r_43__14_,s_r_43__13_,s_r_43__12_,s_r_43__11_,s_r_43__10_,s_r_43__9_,
  s_r_43__8_,s_r_43__7_,s_r_43__6_,s_r_43__5_,s_r_43__4_,s_r_43__3_,s_r_43__2_,s_r_43__1_,
  s_r_43__0_,prod_accum_46__47_,prod_accum_46__46_,prod_accum_46__45_,
  prod_accum_46__44_,prod_accum_46__43_,prod_accum_46__42_,prod_accum_46__41_,
  prod_accum_46__40_,prod_accum_46__39_,prod_accum_46__38_,prod_accum_46__37_,prod_accum_46__36_,
  prod_accum_46__35_,prod_accum_46__34_,prod_accum_46__33_,prod_accum_46__32_,
  prod_accum_46__31_,prod_accum_46__30_,prod_accum_46__29_,prod_accum_46__28_,
  prod_accum_46__27_,prod_accum_46__26_,prod_accum_46__25_,prod_accum_46__24_,
  prod_accum_46__23_,prod_accum_46__22_,prod_accum_46__21_,prod_accum_46__20_,
  prod_accum_46__19_,prod_accum_46__18_,prod_accum_46__17_,prod_accum_46__16_,prod_accum_46__15_,
  prod_accum_46__14_,prod_accum_46__13_,prod_accum_46__12_,prod_accum_46__11_,
  prod_accum_46__10_,prod_accum_46__9_,prod_accum_46__8_,prod_accum_46__7_,
  prod_accum_46__6_,prod_accum_46__5_,prod_accum_46__4_,prod_accum_46__3_,prod_accum_46__2_,
  prod_accum_46__1_,prod_accum_46__0_,prod_accum_45__46_,prod_accum_45__45_,
  prod_accum_45__44_,prod_accum_45__43_,prod_accum_45__42_,prod_accum_45__41_,
  prod_accum_45__40_,prod_accum_45__39_,prod_accum_45__38_,prod_accum_45__37_,
  prod_accum_45__36_,prod_accum_45__35_,prod_accum_45__34_,prod_accum_45__33_,prod_accum_45__32_,
  prod_accum_45__31_,prod_accum_45__30_,prod_accum_45__29_,prod_accum_45__28_,
  prod_accum_45__27_,prod_accum_45__26_,prod_accum_45__25_,prod_accum_45__24_,
  prod_accum_45__23_,prod_accum_45__22_,prod_accum_45__21_,prod_accum_45__20_,
  prod_accum_45__19_,prod_accum_45__18_,prod_accum_45__17_,prod_accum_45__16_,prod_accum_45__15_,
  prod_accum_45__14_,prod_accum_45__13_,prod_accum_45__12_,prod_accum_45__11_,
  prod_accum_45__10_,prod_accum_45__9_,prod_accum_45__8_,prod_accum_45__7_,
  prod_accum_45__6_,prod_accum_45__5_,prod_accum_45__4_,prod_accum_45__3_,prod_accum_45__2_,
  prod_accum_45__1_,prod_accum_45__0_,prod_accum_44__45_,prod_accum_44__44_,
  prod_accum_44__43_,prod_accum_44__42_,prod_accum_44__41_,prod_accum_44__40_,
  prod_accum_44__39_,prod_accum_44__38_,prod_accum_44__37_,prod_accum_44__36_,
  prod_accum_44__35_,prod_accum_44__34_,prod_accum_44__33_,prod_accum_44__32_,prod_accum_44__31_,
  prod_accum_44__30_,prod_accum_44__29_,prod_accum_44__28_,prod_accum_44__27_,
  prod_accum_44__26_,prod_accum_44__25_,prod_accum_44__24_,prod_accum_44__23_,
  prod_accum_44__22_,prod_accum_44__21_,prod_accum_44__20_,prod_accum_44__19_,
  prod_accum_44__18_,prod_accum_44__17_,prod_accum_44__16_,prod_accum_44__15_,
  prod_accum_44__14_,prod_accum_44__13_,prod_accum_44__12_,prod_accum_44__11_,prod_accum_44__10_,
  prod_accum_44__9_,prod_accum_44__8_,prod_accum_44__7_,prod_accum_44__6_,
  prod_accum_44__5_,prod_accum_44__4_,prod_accum_44__3_,prod_accum_44__2_,
  prod_accum_44__1_,prod_accum_44__0_,prod_accum_43__44_,prod_accum_43__43_,prod_accum_43__42_,
  prod_accum_43__41_,prod_accum_43__40_,prod_accum_43__39_,prod_accum_43__38_,
  prod_accum_43__37_,prod_accum_43__36_,prod_accum_43__35_,prod_accum_43__34_,
  prod_accum_43__33_,prod_accum_43__32_,prod_accum_43__31_,prod_accum_43__30_,
  prod_accum_43__29_,prod_accum_43__28_,prod_accum_43__27_,prod_accum_43__26_,prod_accum_43__25_,
  prod_accum_43__24_,prod_accum_43__23_,prod_accum_43__22_,prod_accum_43__21_,
  prod_accum_43__20_,prod_accum_43__19_,prod_accum_43__18_,prod_accum_43__17_,
  prod_accum_43__16_,prod_accum_43__15_,prod_accum_43__14_,prod_accum_43__13_,
  prod_accum_43__12_,prod_accum_43__11_,prod_accum_43__10_,prod_accum_43__9_,prod_accum_43__8_,
  prod_accum_43__7_,prod_accum_43__6_,prod_accum_43__5_,prod_accum_43__4_,
  prod_accum_43__3_,prod_accum_43__2_,prod_accum_43__1_,prod_accum_43__0_,s_r_50__127_,
  s_r_50__126_,s_r_50__125_,s_r_50__124_,s_r_50__123_,s_r_50__122_,s_r_50__121_,
  s_r_50__120_,s_r_50__119_,s_r_50__118_,s_r_50__117_,s_r_50__116_,s_r_50__115_,
  s_r_50__114_,s_r_50__113_,s_r_50__112_,s_r_50__111_,s_r_50__110_,s_r_50__109_,
  s_r_50__108_,s_r_50__107_,s_r_50__106_,s_r_50__105_,s_r_50__104_,s_r_50__103_,
  s_r_50__102_,s_r_50__101_,s_r_50__100_,s_r_50__99_,s_r_50__98_,s_r_50__97_,s_r_50__96_,
  s_r_50__95_,s_r_50__94_,s_r_50__93_,s_r_50__92_,s_r_50__91_,s_r_50__90_,s_r_50__89_,
  s_r_50__88_,s_r_50__87_,s_r_50__86_,s_r_50__85_,s_r_50__84_,s_r_50__83_,
  s_r_50__82_,s_r_50__81_,s_r_50__80_,s_r_50__79_,s_r_50__78_,s_r_50__77_,s_r_50__76_,
  s_r_50__75_,s_r_50__74_,s_r_50__73_,s_r_50__72_,s_r_50__71_,s_r_50__70_,s_r_50__69_,
  s_r_50__68_,s_r_50__67_,s_r_50__66_,s_r_50__65_,s_r_50__64_,s_r_50__63_,
  s_r_50__62_,s_r_50__61_,s_r_50__60_,s_r_50__59_,s_r_50__58_,s_r_50__57_,s_r_50__56_,
  s_r_50__55_,s_r_50__54_,s_r_50__53_,s_r_50__52_,s_r_50__51_,s_r_50__50_,s_r_50__49_,
  s_r_50__48_,s_r_50__47_,s_r_50__46_,s_r_50__45_,s_r_50__44_,s_r_50__43_,
  s_r_50__42_,s_r_50__41_,s_r_50__40_,s_r_50__39_,s_r_50__38_,s_r_50__37_,s_r_50__36_,
  s_r_50__35_,s_r_50__34_,s_r_50__33_,s_r_50__32_,s_r_50__31_,s_r_50__30_,s_r_50__29_,
  s_r_50__28_,s_r_50__27_,s_r_50__26_,s_r_50__25_,s_r_50__24_,s_r_50__23_,
  s_r_50__22_,s_r_50__21_,s_r_50__20_,s_r_50__19_,s_r_50__18_,s_r_50__17_,s_r_50__16_,
  s_r_50__15_,s_r_50__14_,s_r_50__13_,s_r_50__12_,s_r_50__11_,s_r_50__10_,s_r_50__9_,
  s_r_50__8_,s_r_50__7_,s_r_50__6_,s_r_50__5_,s_r_50__4_,s_r_50__3_,s_r_50__2_,
  s_r_50__1_,s_r_50__0_,s_r_49__127_,s_r_49__126_,s_r_49__125_,s_r_49__124_,
  s_r_49__123_,s_r_49__122_,s_r_49__121_,s_r_49__120_,s_r_49__119_,s_r_49__118_,
  s_r_49__117_,s_r_49__116_,s_r_49__115_,s_r_49__114_,s_r_49__113_,s_r_49__112_,s_r_49__111_,
  s_r_49__110_,s_r_49__109_,s_r_49__108_,s_r_49__107_,s_r_49__106_,s_r_49__105_,
  s_r_49__104_,s_r_49__103_,s_r_49__102_,s_r_49__101_,s_r_49__100_,s_r_49__99_,
  s_r_49__98_,s_r_49__97_,s_r_49__96_,s_r_49__95_,s_r_49__94_,s_r_49__93_,s_r_49__92_,
  s_r_49__91_,s_r_49__90_,s_r_49__89_,s_r_49__88_,s_r_49__87_,s_r_49__86_,
  s_r_49__85_,s_r_49__84_,s_r_49__83_,s_r_49__82_,s_r_49__81_,s_r_49__80_,s_r_49__79_,
  s_r_49__78_,s_r_49__77_,s_r_49__76_,s_r_49__75_,s_r_49__74_,s_r_49__73_,s_r_49__72_,
  s_r_49__71_,s_r_49__70_,s_r_49__69_,s_r_49__68_,s_r_49__67_,s_r_49__66_,
  s_r_49__65_,s_r_49__64_,s_r_49__63_,s_r_49__62_,s_r_49__61_,s_r_49__60_,s_r_49__59_,
  s_r_49__58_,s_r_49__57_,s_r_49__56_,s_r_49__55_,s_r_49__54_,s_r_49__53_,s_r_49__52_,
  s_r_49__51_,s_r_49__50_,s_r_49__49_,s_r_49__48_,s_r_49__47_,s_r_49__46_,
  s_r_49__45_,s_r_49__44_,s_r_49__43_,s_r_49__42_,s_r_49__41_,s_r_49__40_,s_r_49__39_,
  s_r_49__38_,s_r_49__37_,s_r_49__36_,s_r_49__35_,s_r_49__34_,s_r_49__33_,s_r_49__32_,
  s_r_49__31_,s_r_49__30_,s_r_49__29_,s_r_49__28_,s_r_49__27_,s_r_49__26_,
  s_r_49__25_,s_r_49__24_,s_r_49__23_,s_r_49__22_,s_r_49__21_,s_r_49__20_,s_r_49__19_,
  s_r_49__18_,s_r_49__17_,s_r_49__16_,s_r_49__15_,s_r_49__14_,s_r_49__13_,s_r_49__12_,
  s_r_49__11_,s_r_49__10_,s_r_49__9_,s_r_49__8_,s_r_49__7_,s_r_49__6_,s_r_49__5_,
  s_r_49__4_,s_r_49__3_,s_r_49__2_,s_r_49__1_,s_r_49__0_,s_r_48__127_,s_r_48__126_,
  s_r_48__125_,s_r_48__124_,s_r_48__123_,s_r_48__122_,s_r_48__121_,s_r_48__120_,
  s_r_48__119_,s_r_48__118_,s_r_48__117_,s_r_48__116_,s_r_48__115_,s_r_48__114_,
  s_r_48__113_,s_r_48__112_,s_r_48__111_,s_r_48__110_,s_r_48__109_,s_r_48__108_,
  s_r_48__107_,s_r_48__106_,s_r_48__105_,s_r_48__104_,s_r_48__103_,s_r_48__102_,
  s_r_48__101_,s_r_48__100_,s_r_48__99_,s_r_48__98_,s_r_48__97_,s_r_48__96_,s_r_48__95_,
  s_r_48__94_,s_r_48__93_,s_r_48__92_,s_r_48__91_,s_r_48__90_,s_r_48__89_,s_r_48__88_,
  s_r_48__87_,s_r_48__86_,s_r_48__85_,s_r_48__84_,s_r_48__83_,s_r_48__82_,
  s_r_48__81_,s_r_48__80_,s_r_48__79_,s_r_48__78_,s_r_48__77_,s_r_48__76_,s_r_48__75_,
  s_r_48__74_,s_r_48__73_,s_r_48__72_,s_r_48__71_,s_r_48__70_,s_r_48__69_,s_r_48__68_,
  s_r_48__67_,s_r_48__66_,s_r_48__65_,s_r_48__64_,s_r_48__63_,s_r_48__62_,
  s_r_48__61_,s_r_48__60_,s_r_48__59_,s_r_48__58_,s_r_48__57_,s_r_48__56_,s_r_48__55_,
  s_r_48__54_,s_r_48__53_,s_r_48__52_,s_r_48__51_,s_r_48__50_,s_r_48__49_,s_r_48__48_,
  s_r_48__47_,s_r_48__46_,s_r_48__45_,s_r_48__44_,s_r_48__43_,s_r_48__42_,
  s_r_48__41_,s_r_48__40_,s_r_48__39_,s_r_48__38_,s_r_48__37_,s_r_48__36_,s_r_48__35_,
  s_r_48__34_,s_r_48__33_,s_r_48__32_,s_r_48__31_,s_r_48__30_,s_r_48__29_,s_r_48__28_,
  s_r_48__27_,s_r_48__26_,s_r_48__25_,s_r_48__24_,s_r_48__23_,s_r_48__22_,
  s_r_48__21_,s_r_48__20_,s_r_48__19_,s_r_48__18_,s_r_48__17_,s_r_48__16_,s_r_48__15_,
  s_r_48__14_,s_r_48__13_,s_r_48__12_,s_r_48__11_,s_r_48__10_,s_r_48__9_,s_r_48__8_,
  s_r_48__7_,s_r_48__6_,s_r_48__5_,s_r_48__4_,s_r_48__3_,s_r_48__2_,s_r_48__1_,
  s_r_48__0_,s_r_47__127_,s_r_47__126_,s_r_47__125_,s_r_47__124_,s_r_47__123_,
  s_r_47__122_,s_r_47__121_,s_r_47__120_,s_r_47__119_,s_r_47__118_,s_r_47__117_,
  s_r_47__116_,s_r_47__115_,s_r_47__114_,s_r_47__113_,s_r_47__112_,s_r_47__111_,s_r_47__110_,
  s_r_47__109_,s_r_47__108_,s_r_47__107_,s_r_47__106_,s_r_47__105_,s_r_47__104_,
  s_r_47__103_,s_r_47__102_,s_r_47__101_,s_r_47__100_,s_r_47__99_,s_r_47__98_,
  s_r_47__97_,s_r_47__96_,s_r_47__95_,s_r_47__94_,s_r_47__93_,s_r_47__92_,s_r_47__91_,
  s_r_47__90_,s_r_47__89_,s_r_47__88_,s_r_47__87_,s_r_47__86_,s_r_47__85_,
  s_r_47__84_,s_r_47__83_,s_r_47__82_,s_r_47__81_,s_r_47__80_,s_r_47__79_,s_r_47__78_,
  s_r_47__77_,s_r_47__76_,s_r_47__75_,s_r_47__74_,s_r_47__73_,s_r_47__72_,s_r_47__71_,
  s_r_47__70_,s_r_47__69_,s_r_47__68_,s_r_47__67_,s_r_47__66_,s_r_47__65_,
  s_r_47__64_,s_r_47__63_,s_r_47__62_,s_r_47__61_,s_r_47__60_,s_r_47__59_,s_r_47__58_,
  s_r_47__57_,s_r_47__56_,s_r_47__55_,s_r_47__54_,s_r_47__53_,s_r_47__52_,s_r_47__51_,
  s_r_47__50_,s_r_47__49_,s_r_47__48_,s_r_47__47_,s_r_47__46_,s_r_47__45_,
  s_r_47__44_,s_r_47__43_,s_r_47__42_,s_r_47__41_,s_r_47__40_,s_r_47__39_,s_r_47__38_,
  s_r_47__37_,s_r_47__36_,s_r_47__35_,s_r_47__34_,s_r_47__33_,s_r_47__32_,s_r_47__31_,
  s_r_47__30_,s_r_47__29_,s_r_47__28_,s_r_47__27_,s_r_47__26_,s_r_47__25_,
  s_r_47__24_,s_r_47__23_,s_r_47__22_,s_r_47__21_,s_r_47__20_,s_r_47__19_,s_r_47__18_,
  s_r_47__17_,s_r_47__16_,s_r_47__15_,s_r_47__14_,s_r_47__13_,s_r_47__12_,s_r_47__11_,
  s_r_47__10_,s_r_47__9_,s_r_47__8_,s_r_47__7_,s_r_47__6_,s_r_47__5_,s_r_47__4_,
  s_r_47__3_,s_r_47__2_,s_r_47__1_,s_r_47__0_,prod_accum_50__51_,prod_accum_50__50_,
  prod_accum_50__49_,prod_accum_50__48_,prod_accum_50__47_,prod_accum_50__46_,
  prod_accum_50__45_,prod_accum_50__44_,prod_accum_50__43_,prod_accum_50__42_,
  prod_accum_50__41_,prod_accum_50__40_,prod_accum_50__39_,prod_accum_50__38_,
  prod_accum_50__37_,prod_accum_50__36_,prod_accum_50__35_,prod_accum_50__34_,
  prod_accum_50__33_,prod_accum_50__32_,prod_accum_50__31_,prod_accum_50__30_,prod_accum_50__29_,
  prod_accum_50__28_,prod_accum_50__27_,prod_accum_50__26_,prod_accum_50__25_,
  prod_accum_50__24_,prod_accum_50__23_,prod_accum_50__22_,prod_accum_50__21_,
  prod_accum_50__20_,prod_accum_50__19_,prod_accum_50__18_,prod_accum_50__17_,
  prod_accum_50__16_,prod_accum_50__15_,prod_accum_50__14_,prod_accum_50__13_,prod_accum_50__12_,
  prod_accum_50__11_,prod_accum_50__10_,prod_accum_50__9_,prod_accum_50__8_,
  prod_accum_50__7_,prod_accum_50__6_,prod_accum_50__5_,prod_accum_50__4_,
  prod_accum_50__3_,prod_accum_50__2_,prod_accum_50__1_,prod_accum_50__0_,prod_accum_49__50_,
  prod_accum_49__49_,prod_accum_49__48_,prod_accum_49__47_,prod_accum_49__46_,
  prod_accum_49__45_,prod_accum_49__44_,prod_accum_49__43_,prod_accum_49__42_,
  prod_accum_49__41_,prod_accum_49__40_,prod_accum_49__39_,prod_accum_49__38_,
  prod_accum_49__37_,prod_accum_49__36_,prod_accum_49__35_,prod_accum_49__34_,prod_accum_49__33_,
  prod_accum_49__32_,prod_accum_49__31_,prod_accum_49__30_,prod_accum_49__29_,
  prod_accum_49__28_,prod_accum_49__27_,prod_accum_49__26_,prod_accum_49__25_,
  prod_accum_49__24_,prod_accum_49__23_,prod_accum_49__22_,prod_accum_49__21_,
  prod_accum_49__20_,prod_accum_49__19_,prod_accum_49__18_,prod_accum_49__17_,
  prod_accum_49__16_,prod_accum_49__15_,prod_accum_49__14_,prod_accum_49__13_,prod_accum_49__12_,
  prod_accum_49__11_,prod_accum_49__10_,prod_accum_49__9_,prod_accum_49__8_,
  prod_accum_49__7_,prod_accum_49__6_,prod_accum_49__5_,prod_accum_49__4_,
  prod_accum_49__3_,prod_accum_49__2_,prod_accum_49__1_,prod_accum_49__0_,prod_accum_48__49_,
  prod_accum_48__48_,prod_accum_48__47_,prod_accum_48__46_,prod_accum_48__45_,
  prod_accum_48__44_,prod_accum_48__43_,prod_accum_48__42_,prod_accum_48__41_,
  prod_accum_48__40_,prod_accum_48__39_,prod_accum_48__38_,prod_accum_48__37_,
  prod_accum_48__36_,prod_accum_48__35_,prod_accum_48__34_,prod_accum_48__33_,prod_accum_48__32_,
  prod_accum_48__31_,prod_accum_48__30_,prod_accum_48__29_,prod_accum_48__28_,
  prod_accum_48__27_,prod_accum_48__26_,prod_accum_48__25_,prod_accum_48__24_,
  prod_accum_48__23_,prod_accum_48__22_,prod_accum_48__21_,prod_accum_48__20_,
  prod_accum_48__19_,prod_accum_48__18_,prod_accum_48__17_,prod_accum_48__16_,
  prod_accum_48__15_,prod_accum_48__14_,prod_accum_48__13_,prod_accum_48__12_,prod_accum_48__11_,
  prod_accum_48__10_,prod_accum_48__9_,prod_accum_48__8_,prod_accum_48__7_,
  prod_accum_48__6_,prod_accum_48__5_,prod_accum_48__4_,prod_accum_48__3_,
  prod_accum_48__2_,prod_accum_48__1_,prod_accum_48__0_,prod_accum_47__48_,prod_accum_47__47_,
  prod_accum_47__46_,prod_accum_47__45_,prod_accum_47__44_,prod_accum_47__43_,
  prod_accum_47__42_,prod_accum_47__41_,prod_accum_47__40_,prod_accum_47__39_,
  prod_accum_47__38_,prod_accum_47__37_,prod_accum_47__36_,prod_accum_47__35_,
  prod_accum_47__34_,prod_accum_47__33_,prod_accum_47__32_,prod_accum_47__31_,prod_accum_47__30_,
  prod_accum_47__29_,prod_accum_47__28_,prod_accum_47__27_,prod_accum_47__26_,
  prod_accum_47__25_,prod_accum_47__24_,prod_accum_47__23_,prod_accum_47__22_,
  prod_accum_47__21_,prod_accum_47__20_,prod_accum_47__19_,prod_accum_47__18_,
  prod_accum_47__17_,prod_accum_47__16_,prod_accum_47__15_,prod_accum_47__14_,
  prod_accum_47__13_,prod_accum_47__12_,prod_accum_47__11_,prod_accum_47__10_,prod_accum_47__9_,
  prod_accum_47__8_,prod_accum_47__7_,prod_accum_47__6_,prod_accum_47__5_,
  prod_accum_47__4_,prod_accum_47__3_,prod_accum_47__2_,prod_accum_47__1_,prod_accum_47__0_,
  s_r_54__127_,s_r_54__126_,s_r_54__125_,s_r_54__124_,s_r_54__123_,s_r_54__122_,
  s_r_54__121_,s_r_54__120_,s_r_54__119_,s_r_54__118_,s_r_54__117_,s_r_54__116_,
  s_r_54__115_,s_r_54__114_,s_r_54__113_,s_r_54__112_,s_r_54__111_,s_r_54__110_,
  s_r_54__109_,s_r_54__108_,s_r_54__107_,s_r_54__106_,s_r_54__105_,s_r_54__104_,
  s_r_54__103_,s_r_54__102_,s_r_54__101_,s_r_54__100_,s_r_54__99_,s_r_54__98_,s_r_54__97_,
  s_r_54__96_,s_r_54__95_,s_r_54__94_,s_r_54__93_,s_r_54__92_,s_r_54__91_,
  s_r_54__90_,s_r_54__89_,s_r_54__88_,s_r_54__87_,s_r_54__86_,s_r_54__85_,s_r_54__84_,
  s_r_54__83_,s_r_54__82_,s_r_54__81_,s_r_54__80_,s_r_54__79_,s_r_54__78_,s_r_54__77_,
  s_r_54__76_,s_r_54__75_,s_r_54__74_,s_r_54__73_,s_r_54__72_,s_r_54__71_,
  s_r_54__70_,s_r_54__69_,s_r_54__68_,s_r_54__67_,s_r_54__66_,s_r_54__65_,s_r_54__64_,
  s_r_54__63_,s_r_54__62_,s_r_54__61_,s_r_54__60_,s_r_54__59_,s_r_54__58_,s_r_54__57_,
  s_r_54__56_,s_r_54__55_,s_r_54__54_,s_r_54__53_,s_r_54__52_,s_r_54__51_,
  s_r_54__50_,s_r_54__49_,s_r_54__48_,s_r_54__47_,s_r_54__46_,s_r_54__45_,s_r_54__44_,
  s_r_54__43_,s_r_54__42_,s_r_54__41_,s_r_54__40_,s_r_54__39_,s_r_54__38_,s_r_54__37_,
  s_r_54__36_,s_r_54__35_,s_r_54__34_,s_r_54__33_,s_r_54__32_,s_r_54__31_,
  s_r_54__30_,s_r_54__29_,s_r_54__28_,s_r_54__27_,s_r_54__26_,s_r_54__25_,s_r_54__24_,
  s_r_54__23_,s_r_54__22_,s_r_54__21_,s_r_54__20_,s_r_54__19_,s_r_54__18_,s_r_54__17_,
  s_r_54__16_,s_r_54__15_,s_r_54__14_,s_r_54__13_,s_r_54__12_,s_r_54__11_,
  s_r_54__10_,s_r_54__9_,s_r_54__8_,s_r_54__7_,s_r_54__6_,s_r_54__5_,s_r_54__4_,s_r_54__3_,
  s_r_54__2_,s_r_54__1_,s_r_54__0_,s_r_53__127_,s_r_53__126_,s_r_53__125_,
  s_r_53__124_,s_r_53__123_,s_r_53__122_,s_r_53__121_,s_r_53__120_,s_r_53__119_,
  s_r_53__118_,s_r_53__117_,s_r_53__116_,s_r_53__115_,s_r_53__114_,s_r_53__113_,s_r_53__112_,
  s_r_53__111_,s_r_53__110_,s_r_53__109_,s_r_53__108_,s_r_53__107_,s_r_53__106_,
  s_r_53__105_,s_r_53__104_,s_r_53__103_,s_r_53__102_,s_r_53__101_,s_r_53__100_,
  s_r_53__99_,s_r_53__98_,s_r_53__97_,s_r_53__96_,s_r_53__95_,s_r_53__94_,s_r_53__93_,
  s_r_53__92_,s_r_53__91_,s_r_53__90_,s_r_53__89_,s_r_53__88_,s_r_53__87_,
  s_r_53__86_,s_r_53__85_,s_r_53__84_,s_r_53__83_,s_r_53__82_,s_r_53__81_,s_r_53__80_,
  s_r_53__79_,s_r_53__78_,s_r_53__77_,s_r_53__76_,s_r_53__75_,s_r_53__74_,s_r_53__73_,
  s_r_53__72_,s_r_53__71_,s_r_53__70_,s_r_53__69_,s_r_53__68_,s_r_53__67_,
  s_r_53__66_,s_r_53__65_,s_r_53__64_,s_r_53__63_,s_r_53__62_,s_r_53__61_,s_r_53__60_,
  s_r_53__59_,s_r_53__58_,s_r_53__57_,s_r_53__56_,s_r_53__55_,s_r_53__54_,s_r_53__53_,
  s_r_53__52_,s_r_53__51_,s_r_53__50_,s_r_53__49_,s_r_53__48_,s_r_53__47_,
  s_r_53__46_,s_r_53__45_,s_r_53__44_,s_r_53__43_,s_r_53__42_,s_r_53__41_,s_r_53__40_,
  s_r_53__39_,s_r_53__38_,s_r_53__37_,s_r_53__36_,s_r_53__35_,s_r_53__34_,s_r_53__33_,
  s_r_53__32_,s_r_53__31_,s_r_53__30_,s_r_53__29_,s_r_53__28_,s_r_53__27_,
  s_r_53__26_,s_r_53__25_,s_r_53__24_,s_r_53__23_,s_r_53__22_,s_r_53__21_,s_r_53__20_,
  s_r_53__19_,s_r_53__18_,s_r_53__17_,s_r_53__16_,s_r_53__15_,s_r_53__14_,s_r_53__13_,
  s_r_53__12_,s_r_53__11_,s_r_53__10_,s_r_53__9_,s_r_53__8_,s_r_53__7_,s_r_53__6_,
  s_r_53__5_,s_r_53__4_,s_r_53__3_,s_r_53__2_,s_r_53__1_,s_r_53__0_,s_r_52__127_,
  s_r_52__126_,s_r_52__125_,s_r_52__124_,s_r_52__123_,s_r_52__122_,s_r_52__121_,
  s_r_52__120_,s_r_52__119_,s_r_52__118_,s_r_52__117_,s_r_52__116_,s_r_52__115_,
  s_r_52__114_,s_r_52__113_,s_r_52__112_,s_r_52__111_,s_r_52__110_,s_r_52__109_,
  s_r_52__108_,s_r_52__107_,s_r_52__106_,s_r_52__105_,s_r_52__104_,s_r_52__103_,
  s_r_52__102_,s_r_52__101_,s_r_52__100_,s_r_52__99_,s_r_52__98_,s_r_52__97_,s_r_52__96_,
  s_r_52__95_,s_r_52__94_,s_r_52__93_,s_r_52__92_,s_r_52__91_,s_r_52__90_,
  s_r_52__89_,s_r_52__88_,s_r_52__87_,s_r_52__86_,s_r_52__85_,s_r_52__84_,s_r_52__83_,
  s_r_52__82_,s_r_52__81_,s_r_52__80_,s_r_52__79_,s_r_52__78_,s_r_52__77_,s_r_52__76_,
  s_r_52__75_,s_r_52__74_,s_r_52__73_,s_r_52__72_,s_r_52__71_,s_r_52__70_,
  s_r_52__69_,s_r_52__68_,s_r_52__67_,s_r_52__66_,s_r_52__65_,s_r_52__64_,s_r_52__63_,
  s_r_52__62_,s_r_52__61_,s_r_52__60_,s_r_52__59_,s_r_52__58_,s_r_52__57_,s_r_52__56_,
  s_r_52__55_,s_r_52__54_,s_r_52__53_,s_r_52__52_,s_r_52__51_,s_r_52__50_,
  s_r_52__49_,s_r_52__48_,s_r_52__47_,s_r_52__46_,s_r_52__45_,s_r_52__44_,s_r_52__43_,
  s_r_52__42_,s_r_52__41_,s_r_52__40_,s_r_52__39_,s_r_52__38_,s_r_52__37_,s_r_52__36_,
  s_r_52__35_,s_r_52__34_,s_r_52__33_,s_r_52__32_,s_r_52__31_,s_r_52__30_,
  s_r_52__29_,s_r_52__28_,s_r_52__27_,s_r_52__26_,s_r_52__25_,s_r_52__24_,s_r_52__23_,
  s_r_52__22_,s_r_52__21_,s_r_52__20_,s_r_52__19_,s_r_52__18_,s_r_52__17_,s_r_52__16_,
  s_r_52__15_,s_r_52__14_,s_r_52__13_,s_r_52__12_,s_r_52__11_,s_r_52__10_,
  s_r_52__9_,s_r_52__8_,s_r_52__7_,s_r_52__6_,s_r_52__5_,s_r_52__4_,s_r_52__3_,s_r_52__2_,
  s_r_52__1_,s_r_52__0_,s_r_51__127_,s_r_51__126_,s_r_51__125_,s_r_51__124_,
  s_r_51__123_,s_r_51__122_,s_r_51__121_,s_r_51__120_,s_r_51__119_,s_r_51__118_,
  s_r_51__117_,s_r_51__116_,s_r_51__115_,s_r_51__114_,s_r_51__113_,s_r_51__112_,
  s_r_51__111_,s_r_51__110_,s_r_51__109_,s_r_51__108_,s_r_51__107_,s_r_51__106_,s_r_51__105_,
  s_r_51__104_,s_r_51__103_,s_r_51__102_,s_r_51__101_,s_r_51__100_,s_r_51__99_,
  s_r_51__98_,s_r_51__97_,s_r_51__96_,s_r_51__95_,s_r_51__94_,s_r_51__93_,s_r_51__92_,
  s_r_51__91_,s_r_51__90_,s_r_51__89_,s_r_51__88_,s_r_51__87_,s_r_51__86_,
  s_r_51__85_,s_r_51__84_,s_r_51__83_,s_r_51__82_,s_r_51__81_,s_r_51__80_,s_r_51__79_,
  s_r_51__78_,s_r_51__77_,s_r_51__76_,s_r_51__75_,s_r_51__74_,s_r_51__73_,s_r_51__72_,
  s_r_51__71_,s_r_51__70_,s_r_51__69_,s_r_51__68_,s_r_51__67_,s_r_51__66_,
  s_r_51__65_,s_r_51__64_,s_r_51__63_,s_r_51__62_,s_r_51__61_,s_r_51__60_,s_r_51__59_,
  s_r_51__58_,s_r_51__57_,s_r_51__56_,s_r_51__55_,s_r_51__54_,s_r_51__53_,s_r_51__52_,
  s_r_51__51_,s_r_51__50_,s_r_51__49_,s_r_51__48_,s_r_51__47_,s_r_51__46_,
  s_r_51__45_,s_r_51__44_,s_r_51__43_,s_r_51__42_,s_r_51__41_,s_r_51__40_,s_r_51__39_,
  s_r_51__38_,s_r_51__37_,s_r_51__36_,s_r_51__35_,s_r_51__34_,s_r_51__33_,s_r_51__32_,
  s_r_51__31_,s_r_51__30_,s_r_51__29_,s_r_51__28_,s_r_51__27_,s_r_51__26_,
  s_r_51__25_,s_r_51__24_,s_r_51__23_,s_r_51__22_,s_r_51__21_,s_r_51__20_,s_r_51__19_,
  s_r_51__18_,s_r_51__17_,s_r_51__16_,s_r_51__15_,s_r_51__14_,s_r_51__13_,s_r_51__12_,
  s_r_51__11_,s_r_51__10_,s_r_51__9_,s_r_51__8_,s_r_51__7_,s_r_51__6_,s_r_51__5_,
  s_r_51__4_,s_r_51__3_,s_r_51__2_,s_r_51__1_,s_r_51__0_,prod_accum_54__55_,
  prod_accum_54__54_,prod_accum_54__53_,prod_accum_54__52_,prod_accum_54__51_,
  prod_accum_54__50_,prod_accum_54__49_,prod_accum_54__48_,prod_accum_54__47_,
  prod_accum_54__46_,prod_accum_54__45_,prod_accum_54__44_,prod_accum_54__43_,prod_accum_54__42_,
  prod_accum_54__41_,prod_accum_54__40_,prod_accum_54__39_,prod_accum_54__38_,
  prod_accum_54__37_,prod_accum_54__36_,prod_accum_54__35_,prod_accum_54__34_,
  prod_accum_54__33_,prod_accum_54__32_,prod_accum_54__31_,prod_accum_54__30_,
  prod_accum_54__29_,prod_accum_54__28_,prod_accum_54__27_,prod_accum_54__26_,
  prod_accum_54__25_,prod_accum_54__24_,prod_accum_54__23_,prod_accum_54__22_,prod_accum_54__21_,
  prod_accum_54__20_,prod_accum_54__19_,prod_accum_54__18_,prod_accum_54__17_,
  prod_accum_54__16_,prod_accum_54__15_,prod_accum_54__14_,prod_accum_54__13_,
  prod_accum_54__12_,prod_accum_54__11_,prod_accum_54__10_,prod_accum_54__9_,
  prod_accum_54__8_,prod_accum_54__7_,prod_accum_54__6_,prod_accum_54__5_,prod_accum_54__4_,
  prod_accum_54__3_,prod_accum_54__2_,prod_accum_54__1_,prod_accum_54__0_,
  prod_accum_53__54_,prod_accum_53__53_,prod_accum_53__52_,prod_accum_53__51_,
  prod_accum_53__50_,prod_accum_53__49_,prod_accum_53__48_,prod_accum_53__47_,prod_accum_53__46_,
  prod_accum_53__45_,prod_accum_53__44_,prod_accum_53__43_,prod_accum_53__42_,
  prod_accum_53__41_,prod_accum_53__40_,prod_accum_53__39_,prod_accum_53__38_,
  prod_accum_53__37_,prod_accum_53__36_,prod_accum_53__35_,prod_accum_53__34_,
  prod_accum_53__33_,prod_accum_53__32_,prod_accum_53__31_,prod_accum_53__30_,
  prod_accum_53__29_,prod_accum_53__28_,prod_accum_53__27_,prod_accum_53__26_,prod_accum_53__25_,
  prod_accum_53__24_,prod_accum_53__23_,prod_accum_53__22_,prod_accum_53__21_,
  prod_accum_53__20_,prod_accum_53__19_,prod_accum_53__18_,prod_accum_53__17_,
  prod_accum_53__16_,prod_accum_53__15_,prod_accum_53__14_,prod_accum_53__13_,
  prod_accum_53__12_,prod_accum_53__11_,prod_accum_53__10_,prod_accum_53__9_,prod_accum_53__8_,
  prod_accum_53__7_,prod_accum_53__6_,prod_accum_53__5_,prod_accum_53__4_,
  prod_accum_53__3_,prod_accum_53__2_,prod_accum_53__1_,prod_accum_53__0_,
  prod_accum_52__53_,prod_accum_52__52_,prod_accum_52__51_,prod_accum_52__50_,prod_accum_52__49_,
  prod_accum_52__48_,prod_accum_52__47_,prod_accum_52__46_,prod_accum_52__45_,
  prod_accum_52__44_,prod_accum_52__43_,prod_accum_52__42_,prod_accum_52__41_,
  prod_accum_52__40_,prod_accum_52__39_,prod_accum_52__38_,prod_accum_52__37_,
  prod_accum_52__36_,prod_accum_52__35_,prod_accum_52__34_,prod_accum_52__33_,
  prod_accum_52__32_,prod_accum_52__31_,prod_accum_52__30_,prod_accum_52__29_,prod_accum_52__28_,
  prod_accum_52__27_,prod_accum_52__26_,prod_accum_52__25_,prod_accum_52__24_,
  prod_accum_52__23_,prod_accum_52__22_,prod_accum_52__21_,prod_accum_52__20_,
  prod_accum_52__19_,prod_accum_52__18_,prod_accum_52__17_,prod_accum_52__16_,
  prod_accum_52__15_,prod_accum_52__14_,prod_accum_52__13_,prod_accum_52__12_,prod_accum_52__11_,
  prod_accum_52__10_,prod_accum_52__9_,prod_accum_52__8_,prod_accum_52__7_,
  prod_accum_52__6_,prod_accum_52__5_,prod_accum_52__4_,prod_accum_52__3_,
  prod_accum_52__2_,prod_accum_52__1_,prod_accum_52__0_,prod_accum_51__52_,prod_accum_51__51_,
  prod_accum_51__50_,prod_accum_51__49_,prod_accum_51__48_,prod_accum_51__47_,
  prod_accum_51__46_,prod_accum_51__45_,prod_accum_51__44_,prod_accum_51__43_,
  prod_accum_51__42_,prod_accum_51__41_,prod_accum_51__40_,prod_accum_51__39_,
  prod_accum_51__38_,prod_accum_51__37_,prod_accum_51__36_,prod_accum_51__35_,prod_accum_51__34_,
  prod_accum_51__33_,prod_accum_51__32_,prod_accum_51__31_,prod_accum_51__30_,
  prod_accum_51__29_,prod_accum_51__28_,prod_accum_51__27_,prod_accum_51__26_,
  prod_accum_51__25_,prod_accum_51__24_,prod_accum_51__23_,prod_accum_51__22_,
  prod_accum_51__21_,prod_accum_51__20_,prod_accum_51__19_,prod_accum_51__18_,
  prod_accum_51__17_,prod_accum_51__16_,prod_accum_51__15_,prod_accum_51__14_,prod_accum_51__13_,
  prod_accum_51__12_,prod_accum_51__11_,prod_accum_51__10_,prod_accum_51__9_,
  prod_accum_51__8_,prod_accum_51__7_,prod_accum_51__6_,prod_accum_51__5_,
  prod_accum_51__4_,prod_accum_51__3_,prod_accum_51__2_,prod_accum_51__1_,prod_accum_51__0_,
  s_r_58__127_,s_r_58__126_,s_r_58__125_,s_r_58__124_,s_r_58__123_,s_r_58__122_,
  s_r_58__121_,s_r_58__120_,s_r_58__119_,s_r_58__118_,s_r_58__117_,s_r_58__116_,
  s_r_58__115_,s_r_58__114_,s_r_58__113_,s_r_58__112_,s_r_58__111_,s_r_58__110_,
  s_r_58__109_,s_r_58__108_,s_r_58__107_,s_r_58__106_,s_r_58__105_,s_r_58__104_,
  s_r_58__103_,s_r_58__102_,s_r_58__101_,s_r_58__100_,s_r_58__99_,s_r_58__98_,s_r_58__97_,
  s_r_58__96_,s_r_58__95_,s_r_58__94_,s_r_58__93_,s_r_58__92_,s_r_58__91_,s_r_58__90_,
  s_r_58__89_,s_r_58__88_,s_r_58__87_,s_r_58__86_,s_r_58__85_,s_r_58__84_,
  s_r_58__83_,s_r_58__82_,s_r_58__81_,s_r_58__80_,s_r_58__79_,s_r_58__78_,s_r_58__77_,
  s_r_58__76_,s_r_58__75_,s_r_58__74_,s_r_58__73_,s_r_58__72_,s_r_58__71_,s_r_58__70_,
  s_r_58__69_,s_r_58__68_,s_r_58__67_,s_r_58__66_,s_r_58__65_,s_r_58__64_,
  s_r_58__63_,s_r_58__62_,s_r_58__61_,s_r_58__60_,s_r_58__59_,s_r_58__58_,s_r_58__57_,
  s_r_58__56_,s_r_58__55_,s_r_58__54_,s_r_58__53_,s_r_58__52_,s_r_58__51_,s_r_58__50_,
  s_r_58__49_,s_r_58__48_,s_r_58__47_,s_r_58__46_,s_r_58__45_,s_r_58__44_,
  s_r_58__43_,s_r_58__42_,s_r_58__41_,s_r_58__40_,s_r_58__39_,s_r_58__38_,s_r_58__37_,
  s_r_58__36_,s_r_58__35_,s_r_58__34_,s_r_58__33_,s_r_58__32_,s_r_58__31_,s_r_58__30_,
  s_r_58__29_,s_r_58__28_,s_r_58__27_,s_r_58__26_,s_r_58__25_,s_r_58__24_,
  s_r_58__23_,s_r_58__22_,s_r_58__21_,s_r_58__20_,s_r_58__19_,s_r_58__18_,s_r_58__17_,
  s_r_58__16_,s_r_58__15_,s_r_58__14_,s_r_58__13_,s_r_58__12_,s_r_58__11_,s_r_58__10_,
  s_r_58__9_,s_r_58__8_,s_r_58__7_,s_r_58__6_,s_r_58__5_,s_r_58__4_,s_r_58__3_,
  s_r_58__2_,s_r_58__1_,s_r_58__0_,s_r_57__127_,s_r_57__126_,s_r_57__125_,
  s_r_57__124_,s_r_57__123_,s_r_57__122_,s_r_57__121_,s_r_57__120_,s_r_57__119_,s_r_57__118_,
  s_r_57__117_,s_r_57__116_,s_r_57__115_,s_r_57__114_,s_r_57__113_,s_r_57__112_,
  s_r_57__111_,s_r_57__110_,s_r_57__109_,s_r_57__108_,s_r_57__107_,s_r_57__106_,
  s_r_57__105_,s_r_57__104_,s_r_57__103_,s_r_57__102_,s_r_57__101_,s_r_57__100_,
  s_r_57__99_,s_r_57__98_,s_r_57__97_,s_r_57__96_,s_r_57__95_,s_r_57__94_,s_r_57__93_,
  s_r_57__92_,s_r_57__91_,s_r_57__90_,s_r_57__89_,s_r_57__88_,s_r_57__87_,
  s_r_57__86_,s_r_57__85_,s_r_57__84_,s_r_57__83_,s_r_57__82_,s_r_57__81_,s_r_57__80_,
  s_r_57__79_,s_r_57__78_,s_r_57__77_,s_r_57__76_,s_r_57__75_,s_r_57__74_,s_r_57__73_,
  s_r_57__72_,s_r_57__71_,s_r_57__70_,s_r_57__69_,s_r_57__68_,s_r_57__67_,
  s_r_57__66_,s_r_57__65_,s_r_57__64_,s_r_57__63_,s_r_57__62_,s_r_57__61_,s_r_57__60_,
  s_r_57__59_,s_r_57__58_,s_r_57__57_,s_r_57__56_,s_r_57__55_,s_r_57__54_,s_r_57__53_,
  s_r_57__52_,s_r_57__51_,s_r_57__50_,s_r_57__49_,s_r_57__48_,s_r_57__47_,
  s_r_57__46_,s_r_57__45_,s_r_57__44_,s_r_57__43_,s_r_57__42_,s_r_57__41_,s_r_57__40_,
  s_r_57__39_,s_r_57__38_,s_r_57__37_,s_r_57__36_,s_r_57__35_,s_r_57__34_,s_r_57__33_,
  s_r_57__32_,s_r_57__31_,s_r_57__30_,s_r_57__29_,s_r_57__28_,s_r_57__27_,
  s_r_57__26_,s_r_57__25_,s_r_57__24_,s_r_57__23_,s_r_57__22_,s_r_57__21_,s_r_57__20_,
  s_r_57__19_,s_r_57__18_,s_r_57__17_,s_r_57__16_,s_r_57__15_,s_r_57__14_,s_r_57__13_,
  s_r_57__12_,s_r_57__11_,s_r_57__10_,s_r_57__9_,s_r_57__8_,s_r_57__7_,s_r_57__6_,
  s_r_57__5_,s_r_57__4_,s_r_57__3_,s_r_57__2_,s_r_57__1_,s_r_57__0_,s_r_56__127_,
  s_r_56__126_,s_r_56__125_,s_r_56__124_,s_r_56__123_,s_r_56__122_,s_r_56__121_,
  s_r_56__120_,s_r_56__119_,s_r_56__118_,s_r_56__117_,s_r_56__116_,s_r_56__115_,
  s_r_56__114_,s_r_56__113_,s_r_56__112_,s_r_56__111_,s_r_56__110_,s_r_56__109_,
  s_r_56__108_,s_r_56__107_,s_r_56__106_,s_r_56__105_,s_r_56__104_,s_r_56__103_,
  s_r_56__102_,s_r_56__101_,s_r_56__100_,s_r_56__99_,s_r_56__98_,s_r_56__97_,s_r_56__96_,
  s_r_56__95_,s_r_56__94_,s_r_56__93_,s_r_56__92_,s_r_56__91_,s_r_56__90_,s_r_56__89_,
  s_r_56__88_,s_r_56__87_,s_r_56__86_,s_r_56__85_,s_r_56__84_,s_r_56__83_,
  s_r_56__82_,s_r_56__81_,s_r_56__80_,s_r_56__79_,s_r_56__78_,s_r_56__77_,s_r_56__76_,
  s_r_56__75_,s_r_56__74_,s_r_56__73_,s_r_56__72_,s_r_56__71_,s_r_56__70_,s_r_56__69_,
  s_r_56__68_,s_r_56__67_,s_r_56__66_,s_r_56__65_,s_r_56__64_,s_r_56__63_,
  s_r_56__62_,s_r_56__61_,s_r_56__60_,s_r_56__59_,s_r_56__58_,s_r_56__57_,s_r_56__56_,
  s_r_56__55_,s_r_56__54_,s_r_56__53_,s_r_56__52_,s_r_56__51_,s_r_56__50_,s_r_56__49_,
  s_r_56__48_,s_r_56__47_,s_r_56__46_,s_r_56__45_,s_r_56__44_,s_r_56__43_,
  s_r_56__42_,s_r_56__41_,s_r_56__40_,s_r_56__39_,s_r_56__38_,s_r_56__37_,s_r_56__36_,
  s_r_56__35_,s_r_56__34_,s_r_56__33_,s_r_56__32_,s_r_56__31_,s_r_56__30_,s_r_56__29_,
  s_r_56__28_,s_r_56__27_,s_r_56__26_,s_r_56__25_,s_r_56__24_,s_r_56__23_,
  s_r_56__22_,s_r_56__21_,s_r_56__20_,s_r_56__19_,s_r_56__18_,s_r_56__17_,s_r_56__16_,
  s_r_56__15_,s_r_56__14_,s_r_56__13_,s_r_56__12_,s_r_56__11_,s_r_56__10_,s_r_56__9_,
  s_r_56__8_,s_r_56__7_,s_r_56__6_,s_r_56__5_,s_r_56__4_,s_r_56__3_,s_r_56__2_,
  s_r_56__1_,s_r_56__0_,s_r_55__127_,s_r_55__126_,s_r_55__125_,s_r_55__124_,
  s_r_55__123_,s_r_55__122_,s_r_55__121_,s_r_55__120_,s_r_55__119_,s_r_55__118_,
  s_r_55__117_,s_r_55__116_,s_r_55__115_,s_r_55__114_,s_r_55__113_,s_r_55__112_,s_r_55__111_,
  s_r_55__110_,s_r_55__109_,s_r_55__108_,s_r_55__107_,s_r_55__106_,s_r_55__105_,
  s_r_55__104_,s_r_55__103_,s_r_55__102_,s_r_55__101_,s_r_55__100_,s_r_55__99_,
  s_r_55__98_,s_r_55__97_,s_r_55__96_,s_r_55__95_,s_r_55__94_,s_r_55__93_,s_r_55__92_,
  s_r_55__91_,s_r_55__90_,s_r_55__89_,s_r_55__88_,s_r_55__87_,s_r_55__86_,
  s_r_55__85_,s_r_55__84_,s_r_55__83_,s_r_55__82_,s_r_55__81_,s_r_55__80_,s_r_55__79_,
  s_r_55__78_,s_r_55__77_,s_r_55__76_,s_r_55__75_,s_r_55__74_,s_r_55__73_,s_r_55__72_,
  s_r_55__71_,s_r_55__70_,s_r_55__69_,s_r_55__68_,s_r_55__67_,s_r_55__66_,
  s_r_55__65_,s_r_55__64_,s_r_55__63_,s_r_55__62_,s_r_55__61_,s_r_55__60_,s_r_55__59_,
  s_r_55__58_,s_r_55__57_,s_r_55__56_,s_r_55__55_,s_r_55__54_,s_r_55__53_,s_r_55__52_,
  s_r_55__51_,s_r_55__50_,s_r_55__49_,s_r_55__48_,s_r_55__47_,s_r_55__46_,
  s_r_55__45_,s_r_55__44_,s_r_55__43_,s_r_55__42_,s_r_55__41_,s_r_55__40_,s_r_55__39_,
  s_r_55__38_,s_r_55__37_,s_r_55__36_,s_r_55__35_,s_r_55__34_,s_r_55__33_,s_r_55__32_,
  s_r_55__31_,s_r_55__30_,s_r_55__29_,s_r_55__28_,s_r_55__27_,s_r_55__26_,
  s_r_55__25_,s_r_55__24_,s_r_55__23_,s_r_55__22_,s_r_55__21_,s_r_55__20_,s_r_55__19_,
  s_r_55__18_,s_r_55__17_,s_r_55__16_,s_r_55__15_,s_r_55__14_,s_r_55__13_,s_r_55__12_,
  s_r_55__11_,s_r_55__10_,s_r_55__9_,s_r_55__8_,s_r_55__7_,s_r_55__6_,s_r_55__5_,
  s_r_55__4_,s_r_55__3_,s_r_55__2_,s_r_55__1_,s_r_55__0_,prod_accum_58__59_,
  prod_accum_58__58_,prod_accum_58__57_,prod_accum_58__56_,prod_accum_58__55_,
  prod_accum_58__54_,prod_accum_58__53_,prod_accum_58__52_,prod_accum_58__51_,
  prod_accum_58__50_,prod_accum_58__49_,prod_accum_58__48_,prod_accum_58__47_,prod_accum_58__46_,
  prod_accum_58__45_,prod_accum_58__44_,prod_accum_58__43_,prod_accum_58__42_,
  prod_accum_58__41_,prod_accum_58__40_,prod_accum_58__39_,prod_accum_58__38_,
  prod_accum_58__37_,prod_accum_58__36_,prod_accum_58__35_,prod_accum_58__34_,
  prod_accum_58__33_,prod_accum_58__32_,prod_accum_58__31_,prod_accum_58__30_,
  prod_accum_58__29_,prod_accum_58__28_,prod_accum_58__27_,prod_accum_58__26_,prod_accum_58__25_,
  prod_accum_58__24_,prod_accum_58__23_,prod_accum_58__22_,prod_accum_58__21_,
  prod_accum_58__20_,prod_accum_58__19_,prod_accum_58__18_,prod_accum_58__17_,
  prod_accum_58__16_,prod_accum_58__15_,prod_accum_58__14_,prod_accum_58__13_,
  prod_accum_58__12_,prod_accum_58__11_,prod_accum_58__10_,prod_accum_58__9_,prod_accum_58__8_,
  prod_accum_58__7_,prod_accum_58__6_,prod_accum_58__5_,prod_accum_58__4_,
  prod_accum_58__3_,prod_accum_58__2_,prod_accum_58__1_,prod_accum_58__0_,
  prod_accum_57__58_,prod_accum_57__57_,prod_accum_57__56_,prod_accum_57__55_,prod_accum_57__54_,
  prod_accum_57__53_,prod_accum_57__52_,prod_accum_57__51_,prod_accum_57__50_,
  prod_accum_57__49_,prod_accum_57__48_,prod_accum_57__47_,prod_accum_57__46_,
  prod_accum_57__45_,prod_accum_57__44_,prod_accum_57__43_,prod_accum_57__42_,
  prod_accum_57__41_,prod_accum_57__40_,prod_accum_57__39_,prod_accum_57__38_,prod_accum_57__37_,
  prod_accum_57__36_,prod_accum_57__35_,prod_accum_57__34_,prod_accum_57__33_,
  prod_accum_57__32_,prod_accum_57__31_,prod_accum_57__30_,prod_accum_57__29_,
  prod_accum_57__28_,prod_accum_57__27_,prod_accum_57__26_,prod_accum_57__25_,
  prod_accum_57__24_,prod_accum_57__23_,prod_accum_57__22_,prod_accum_57__21_,
  prod_accum_57__20_,prod_accum_57__19_,prod_accum_57__18_,prod_accum_57__17_,prod_accum_57__16_,
  prod_accum_57__15_,prod_accum_57__14_,prod_accum_57__13_,prod_accum_57__12_,
  prod_accum_57__11_,prod_accum_57__10_,prod_accum_57__9_,prod_accum_57__8_,
  prod_accum_57__7_,prod_accum_57__6_,prod_accum_57__5_,prod_accum_57__4_,prod_accum_57__3_,
  prod_accum_57__2_,prod_accum_57__1_,prod_accum_57__0_,prod_accum_56__57_,
  prod_accum_56__56_,prod_accum_56__55_,prod_accum_56__54_,prod_accum_56__53_,
  prod_accum_56__52_,prod_accum_56__51_,prod_accum_56__50_,prod_accum_56__49_,
  prod_accum_56__48_,prod_accum_56__47_,prod_accum_56__46_,prod_accum_56__45_,prod_accum_56__44_,
  prod_accum_56__43_,prod_accum_56__42_,prod_accum_56__41_,prod_accum_56__40_,
  prod_accum_56__39_,prod_accum_56__38_,prod_accum_56__37_,prod_accum_56__36_,
  prod_accum_56__35_,prod_accum_56__34_,prod_accum_56__33_,prod_accum_56__32_,
  prod_accum_56__31_,prod_accum_56__30_,prod_accum_56__29_,prod_accum_56__28_,
  prod_accum_56__27_,prod_accum_56__26_,prod_accum_56__25_,prod_accum_56__24_,prod_accum_56__23_,
  prod_accum_56__22_,prod_accum_56__21_,prod_accum_56__20_,prod_accum_56__19_,
  prod_accum_56__18_,prod_accum_56__17_,prod_accum_56__16_,prod_accum_56__15_,
  prod_accum_56__14_,prod_accum_56__13_,prod_accum_56__12_,prod_accum_56__11_,
  prod_accum_56__10_,prod_accum_56__9_,prod_accum_56__8_,prod_accum_56__7_,prod_accum_56__6_,
  prod_accum_56__5_,prod_accum_56__4_,prod_accum_56__3_,prod_accum_56__2_,
  prod_accum_56__1_,prod_accum_56__0_,prod_accum_55__56_,prod_accum_55__55_,
  prod_accum_55__54_,prod_accum_55__53_,prod_accum_55__52_,prod_accum_55__51_,prod_accum_55__50_,
  prod_accum_55__49_,prod_accum_55__48_,prod_accum_55__47_,prod_accum_55__46_,
  prod_accum_55__45_,prod_accum_55__44_,prod_accum_55__43_,prod_accum_55__42_,
  prod_accum_55__41_,prod_accum_55__40_,prod_accum_55__39_,prod_accum_55__38_,
  prod_accum_55__37_,prod_accum_55__36_,prod_accum_55__35_,prod_accum_55__34_,
  prod_accum_55__33_,prod_accum_55__32_,prod_accum_55__31_,prod_accum_55__30_,prod_accum_55__29_,
  prod_accum_55__28_,prod_accum_55__27_,prod_accum_55__26_,prod_accum_55__25_,
  prod_accum_55__24_,prod_accum_55__23_,prod_accum_55__22_,prod_accum_55__21_,
  prod_accum_55__20_,prod_accum_55__19_,prod_accum_55__18_,prod_accum_55__17_,
  prod_accum_55__16_,prod_accum_55__15_,prod_accum_55__14_,prod_accum_55__13_,prod_accum_55__12_,
  prod_accum_55__11_,prod_accum_55__10_,prod_accum_55__9_,prod_accum_55__8_,
  prod_accum_55__7_,prod_accum_55__6_,prod_accum_55__5_,prod_accum_55__4_,
  prod_accum_55__3_,prod_accum_55__2_,prod_accum_55__1_,prod_accum_55__0_,s_r_62__127_,
  s_r_62__126_,s_r_62__125_,s_r_62__124_,s_r_62__123_,s_r_62__122_,s_r_62__121_,
  s_r_62__120_,s_r_62__119_,s_r_62__118_,s_r_62__117_,s_r_62__116_,s_r_62__115_,s_r_62__114_,
  s_r_62__113_,s_r_62__112_,s_r_62__111_,s_r_62__110_,s_r_62__109_,s_r_62__108_,
  s_r_62__107_,s_r_62__106_,s_r_62__105_,s_r_62__104_,s_r_62__103_,s_r_62__102_,
  s_r_62__101_,s_r_62__100_,s_r_62__99_,s_r_62__98_,s_r_62__97_,s_r_62__96_,
  s_r_62__95_,s_r_62__94_,s_r_62__93_,s_r_62__92_,s_r_62__91_,s_r_62__90_,s_r_62__89_,
  s_r_62__88_,s_r_62__87_,s_r_62__86_,s_r_62__85_,s_r_62__84_,s_r_62__83_,s_r_62__82_,
  s_r_62__81_,s_r_62__80_,s_r_62__79_,s_r_62__78_,s_r_62__77_,s_r_62__76_,
  s_r_62__75_,s_r_62__74_,s_r_62__73_,s_r_62__72_,s_r_62__71_,s_r_62__70_,s_r_62__69_,
  s_r_62__68_,s_r_62__67_,s_r_62__66_,s_r_62__65_,s_r_62__64_,s_r_62__63_,s_r_62__62_,
  s_r_62__61_,s_r_62__60_,s_r_62__59_,s_r_62__58_,s_r_62__57_,s_r_62__56_,
  s_r_62__55_,s_r_62__54_,s_r_62__53_,s_r_62__52_,s_r_62__51_,s_r_62__50_,s_r_62__49_,
  s_r_62__48_,s_r_62__47_,s_r_62__46_,s_r_62__45_,s_r_62__44_,s_r_62__43_,s_r_62__42_,
  s_r_62__41_,s_r_62__40_,s_r_62__39_,s_r_62__38_,s_r_62__37_,s_r_62__36_,
  s_r_62__35_,s_r_62__34_,s_r_62__33_,s_r_62__32_,s_r_62__31_,s_r_62__30_,s_r_62__29_,
  s_r_62__28_,s_r_62__27_,s_r_62__26_,s_r_62__25_,s_r_62__24_,s_r_62__23_,s_r_62__22_,
  s_r_62__21_,s_r_62__20_,s_r_62__19_,s_r_62__18_,s_r_62__17_,s_r_62__16_,
  s_r_62__15_,s_r_62__14_,s_r_62__13_,s_r_62__12_,s_r_62__11_,s_r_62__10_,s_r_62__9_,
  s_r_62__8_,s_r_62__7_,s_r_62__6_,s_r_62__5_,s_r_62__4_,s_r_62__3_,s_r_62__2_,
  s_r_62__1_,s_r_62__0_,s_r_61__127_,s_r_61__126_,s_r_61__125_,s_r_61__124_,s_r_61__123_,
  s_r_61__122_,s_r_61__121_,s_r_61__120_,s_r_61__119_,s_r_61__118_,s_r_61__117_,
  s_r_61__116_,s_r_61__115_,s_r_61__114_,s_r_61__113_,s_r_61__112_,s_r_61__111_,
  s_r_61__110_,s_r_61__109_,s_r_61__108_,s_r_61__107_,s_r_61__106_,s_r_61__105_,
  s_r_61__104_,s_r_61__103_,s_r_61__102_,s_r_61__101_,s_r_61__100_,s_r_61__99_,s_r_61__98_,
  s_r_61__97_,s_r_61__96_,s_r_61__95_,s_r_61__94_,s_r_61__93_,s_r_61__92_,
  s_r_61__91_,s_r_61__90_,s_r_61__89_,s_r_61__88_,s_r_61__87_,s_r_61__86_,s_r_61__85_,
  s_r_61__84_,s_r_61__83_,s_r_61__82_,s_r_61__81_,s_r_61__80_,s_r_61__79_,s_r_61__78_,
  s_r_61__77_,s_r_61__76_,s_r_61__75_,s_r_61__74_,s_r_61__73_,s_r_61__72_,
  s_r_61__71_,s_r_61__70_,s_r_61__69_,s_r_61__68_,s_r_61__67_,s_r_61__66_,s_r_61__65_,
  s_r_61__64_,s_r_61__63_,s_r_61__62_,s_r_61__61_,s_r_61__60_,s_r_61__59_,s_r_61__58_,
  s_r_61__57_,s_r_61__56_,s_r_61__55_,s_r_61__54_,s_r_61__53_,s_r_61__52_,
  s_r_61__51_,s_r_61__50_,s_r_61__49_,s_r_61__48_,s_r_61__47_,s_r_61__46_,s_r_61__45_,
  s_r_61__44_,s_r_61__43_,s_r_61__42_,s_r_61__41_,s_r_61__40_,s_r_61__39_,s_r_61__38_,
  s_r_61__37_,s_r_61__36_,s_r_61__35_,s_r_61__34_,s_r_61__33_,s_r_61__32_,
  s_r_61__31_,s_r_61__30_,s_r_61__29_,s_r_61__28_,s_r_61__27_,s_r_61__26_,s_r_61__25_,
  s_r_61__24_,s_r_61__23_,s_r_61__22_,s_r_61__21_,s_r_61__20_,s_r_61__19_,s_r_61__18_,
  s_r_61__17_,s_r_61__16_,s_r_61__15_,s_r_61__14_,s_r_61__13_,s_r_61__12_,
  s_r_61__11_,s_r_61__10_,s_r_61__9_,s_r_61__8_,s_r_61__7_,s_r_61__6_,s_r_61__5_,
  s_r_61__4_,s_r_61__3_,s_r_61__2_,s_r_61__1_,s_r_61__0_,s_r_60__127_,s_r_60__126_,
  s_r_60__125_,s_r_60__124_,s_r_60__123_,s_r_60__122_,s_r_60__121_,s_r_60__120_,
  s_r_60__119_,s_r_60__118_,s_r_60__117_,s_r_60__116_,s_r_60__115_,s_r_60__114_,
  s_r_60__113_,s_r_60__112_,s_r_60__111_,s_r_60__110_,s_r_60__109_,s_r_60__108_,s_r_60__107_,
  s_r_60__106_,s_r_60__105_,s_r_60__104_,s_r_60__103_,s_r_60__102_,s_r_60__101_,
  s_r_60__100_,s_r_60__99_,s_r_60__98_,s_r_60__97_,s_r_60__96_,s_r_60__95_,
  s_r_60__94_,s_r_60__93_,s_r_60__92_,s_r_60__91_,s_r_60__90_,s_r_60__89_,s_r_60__88_,
  s_r_60__87_,s_r_60__86_,s_r_60__85_,s_r_60__84_,s_r_60__83_,s_r_60__82_,s_r_60__81_,
  s_r_60__80_,s_r_60__79_,s_r_60__78_,s_r_60__77_,s_r_60__76_,s_r_60__75_,
  s_r_60__74_,s_r_60__73_,s_r_60__72_,s_r_60__71_,s_r_60__70_,s_r_60__69_,s_r_60__68_,
  s_r_60__67_,s_r_60__66_,s_r_60__65_,s_r_60__64_,s_r_60__63_,s_r_60__62_,s_r_60__61_,
  s_r_60__60_,s_r_60__59_,s_r_60__58_,s_r_60__57_,s_r_60__56_,s_r_60__55_,
  s_r_60__54_,s_r_60__53_,s_r_60__52_,s_r_60__51_,s_r_60__50_,s_r_60__49_,s_r_60__48_,
  s_r_60__47_,s_r_60__46_,s_r_60__45_,s_r_60__44_,s_r_60__43_,s_r_60__42_,s_r_60__41_,
  s_r_60__40_,s_r_60__39_,s_r_60__38_,s_r_60__37_,s_r_60__36_,s_r_60__35_,
  s_r_60__34_,s_r_60__33_,s_r_60__32_,s_r_60__31_,s_r_60__30_,s_r_60__29_,s_r_60__28_,
  s_r_60__27_,s_r_60__26_,s_r_60__25_,s_r_60__24_,s_r_60__23_,s_r_60__22_,s_r_60__21_,
  s_r_60__20_,s_r_60__19_,s_r_60__18_,s_r_60__17_,s_r_60__16_,s_r_60__15_,
  s_r_60__14_,s_r_60__13_,s_r_60__12_,s_r_60__11_,s_r_60__10_,s_r_60__9_,s_r_60__8_,
  s_r_60__7_,s_r_60__6_,s_r_60__5_,s_r_60__4_,s_r_60__3_,s_r_60__2_,s_r_60__1_,s_r_60__0_,
  s_r_59__127_,s_r_59__126_,s_r_59__125_,s_r_59__124_,s_r_59__123_,s_r_59__122_,
  s_r_59__121_,s_r_59__120_,s_r_59__119_,s_r_59__118_,s_r_59__117_,s_r_59__116_,
  s_r_59__115_,s_r_59__114_,s_r_59__113_,s_r_59__112_,s_r_59__111_,s_r_59__110_,
  s_r_59__109_,s_r_59__108_,s_r_59__107_,s_r_59__106_,s_r_59__105_,s_r_59__104_,
  s_r_59__103_,s_r_59__102_,s_r_59__101_,s_r_59__100_,s_r_59__99_,s_r_59__98_,s_r_59__97_,
  s_r_59__96_,s_r_59__95_,s_r_59__94_,s_r_59__93_,s_r_59__92_,s_r_59__91_,
  s_r_59__90_,s_r_59__89_,s_r_59__88_,s_r_59__87_,s_r_59__86_,s_r_59__85_,s_r_59__84_,
  s_r_59__83_,s_r_59__82_,s_r_59__81_,s_r_59__80_,s_r_59__79_,s_r_59__78_,s_r_59__77_,
  s_r_59__76_,s_r_59__75_,s_r_59__74_,s_r_59__73_,s_r_59__72_,s_r_59__71_,
  s_r_59__70_,s_r_59__69_,s_r_59__68_,s_r_59__67_,s_r_59__66_,s_r_59__65_,s_r_59__64_,
  s_r_59__63_,s_r_59__62_,s_r_59__61_,s_r_59__60_,s_r_59__59_,s_r_59__58_,s_r_59__57_,
  s_r_59__56_,s_r_59__55_,s_r_59__54_,s_r_59__53_,s_r_59__52_,s_r_59__51_,
  s_r_59__50_,s_r_59__49_,s_r_59__48_,s_r_59__47_,s_r_59__46_,s_r_59__45_,s_r_59__44_,
  s_r_59__43_,s_r_59__42_,s_r_59__41_,s_r_59__40_,s_r_59__39_,s_r_59__38_,s_r_59__37_,
  s_r_59__36_,s_r_59__35_,s_r_59__34_,s_r_59__33_,s_r_59__32_,s_r_59__31_,
  s_r_59__30_,s_r_59__29_,s_r_59__28_,s_r_59__27_,s_r_59__26_,s_r_59__25_,s_r_59__24_,
  s_r_59__23_,s_r_59__22_,s_r_59__21_,s_r_59__20_,s_r_59__19_,s_r_59__18_,s_r_59__17_,
  s_r_59__16_,s_r_59__15_,s_r_59__14_,s_r_59__13_,s_r_59__12_,s_r_59__11_,
  s_r_59__10_,s_r_59__9_,s_r_59__8_,s_r_59__7_,s_r_59__6_,s_r_59__5_,s_r_59__4_,
  s_r_59__3_,s_r_59__2_,s_r_59__1_,s_r_59__0_,prod_accum_62__63_,prod_accum_62__62_,
  prod_accum_62__61_,prod_accum_62__60_,prod_accum_62__59_,prod_accum_62__58_,
  prod_accum_62__57_,prod_accum_62__56_,prod_accum_62__55_,prod_accum_62__54_,
  prod_accum_62__53_,prod_accum_62__52_,prod_accum_62__51_,prod_accum_62__50_,prod_accum_62__49_,
  prod_accum_62__48_,prod_accum_62__47_,prod_accum_62__46_,prod_accum_62__45_,
  prod_accum_62__44_,prod_accum_62__43_,prod_accum_62__42_,prod_accum_62__41_,
  prod_accum_62__40_,prod_accum_62__39_,prod_accum_62__38_,prod_accum_62__37_,
  prod_accum_62__36_,prod_accum_62__35_,prod_accum_62__34_,prod_accum_62__33_,
  prod_accum_62__32_,prod_accum_62__31_,prod_accum_62__30_,prod_accum_62__29_,prod_accum_62__28_,
  prod_accum_62__27_,prod_accum_62__26_,prod_accum_62__25_,prod_accum_62__24_,
  prod_accum_62__23_,prod_accum_62__22_,prod_accum_62__21_,prod_accum_62__20_,
  prod_accum_62__19_,prod_accum_62__18_,prod_accum_62__17_,prod_accum_62__16_,
  prod_accum_62__15_,prod_accum_62__14_,prod_accum_62__13_,prod_accum_62__12_,
  prod_accum_62__11_,prod_accum_62__10_,prod_accum_62__9_,prod_accum_62__8_,prod_accum_62__7_,
  prod_accum_62__6_,prod_accum_62__5_,prod_accum_62__4_,prod_accum_62__3_,
  prod_accum_62__2_,prod_accum_62__1_,prod_accum_62__0_,prod_accum_61__62_,prod_accum_61__61_,
  prod_accum_61__60_,prod_accum_61__59_,prod_accum_61__58_,prod_accum_61__57_,
  prod_accum_61__56_,prod_accum_61__55_,prod_accum_61__54_,prod_accum_61__53_,
  prod_accum_61__52_,prod_accum_61__51_,prod_accum_61__50_,prod_accum_61__49_,
  prod_accum_61__48_,prod_accum_61__47_,prod_accum_61__46_,prod_accum_61__45_,
  prod_accum_61__44_,prod_accum_61__43_,prod_accum_61__42_,prod_accum_61__41_,prod_accum_61__40_,
  prod_accum_61__39_,prod_accum_61__38_,prod_accum_61__37_,prod_accum_61__36_,
  prod_accum_61__35_,prod_accum_61__34_,prod_accum_61__33_,prod_accum_61__32_,
  prod_accum_61__31_,prod_accum_61__30_,prod_accum_61__29_,prod_accum_61__28_,
  prod_accum_61__27_,prod_accum_61__26_,prod_accum_61__25_,prod_accum_61__24_,prod_accum_61__23_,
  prod_accum_61__22_,prod_accum_61__21_,prod_accum_61__20_,prod_accum_61__19_,
  prod_accum_61__18_,prod_accum_61__17_,prod_accum_61__16_,prod_accum_61__15_,
  prod_accum_61__14_,prod_accum_61__13_,prod_accum_61__12_,prod_accum_61__11_,
  prod_accum_61__10_,prod_accum_61__9_,prod_accum_61__8_,prod_accum_61__7_,prod_accum_61__6_,
  prod_accum_61__5_,prod_accum_61__4_,prod_accum_61__3_,prod_accum_61__2_,
  prod_accum_61__1_,prod_accum_61__0_,prod_accum_60__61_,prod_accum_60__60_,
  prod_accum_60__59_,prod_accum_60__58_,prod_accum_60__57_,prod_accum_60__56_,prod_accum_60__55_,
  prod_accum_60__54_,prod_accum_60__53_,prod_accum_60__52_,prod_accum_60__51_,
  prod_accum_60__50_,prod_accum_60__49_,prod_accum_60__48_,prod_accum_60__47_,
  prod_accum_60__46_,prod_accum_60__45_,prod_accum_60__44_,prod_accum_60__43_,
  prod_accum_60__42_,prod_accum_60__41_,prod_accum_60__40_,prod_accum_60__39_,
  prod_accum_60__38_,prod_accum_60__37_,prod_accum_60__36_,prod_accum_60__35_,prod_accum_60__34_,
  prod_accum_60__33_,prod_accum_60__32_,prod_accum_60__31_,prod_accum_60__30_,
  prod_accum_60__29_,prod_accum_60__28_,prod_accum_60__27_,prod_accum_60__26_,
  prod_accum_60__25_,prod_accum_60__24_,prod_accum_60__23_,prod_accum_60__22_,
  prod_accum_60__21_,prod_accum_60__20_,prod_accum_60__19_,prod_accum_60__18_,
  prod_accum_60__17_,prod_accum_60__16_,prod_accum_60__15_,prod_accum_60__14_,prod_accum_60__13_,
  prod_accum_60__12_,prod_accum_60__11_,prod_accum_60__10_,prod_accum_60__9_,
  prod_accum_60__8_,prod_accum_60__7_,prod_accum_60__6_,prod_accum_60__5_,
  prod_accum_60__4_,prod_accum_60__3_,prod_accum_60__2_,prod_accum_60__1_,prod_accum_60__0_,
  prod_accum_59__60_,prod_accum_59__59_,prod_accum_59__58_,prod_accum_59__57_,
  prod_accum_59__56_,prod_accum_59__55_,prod_accum_59__54_,prod_accum_59__53_,
  prod_accum_59__52_,prod_accum_59__51_,prod_accum_59__50_,prod_accum_59__49_,
  prod_accum_59__48_,prod_accum_59__47_,prod_accum_59__46_,prod_accum_59__45_,prod_accum_59__44_,
  prod_accum_59__43_,prod_accum_59__42_,prod_accum_59__41_,prod_accum_59__40_,
  prod_accum_59__39_,prod_accum_59__38_,prod_accum_59__37_,prod_accum_59__36_,
  prod_accum_59__35_,prod_accum_59__34_,prod_accum_59__33_,prod_accum_59__32_,
  prod_accum_59__31_,prod_accum_59__30_,prod_accum_59__29_,prod_accum_59__28_,
  prod_accum_59__27_,prod_accum_59__26_,prod_accum_59__25_,prod_accum_59__24_,prod_accum_59__23_,
  prod_accum_59__22_,prod_accum_59__21_,prod_accum_59__20_,prod_accum_59__19_,
  prod_accum_59__18_,prod_accum_59__17_,prod_accum_59__16_,prod_accum_59__15_,
  prod_accum_59__14_,prod_accum_59__13_,prod_accum_59__12_,prod_accum_59__11_,
  prod_accum_59__10_,prod_accum_59__9_,prod_accum_59__8_,prod_accum_59__7_,prod_accum_59__6_,
  prod_accum_59__5_,prod_accum_59__4_,prod_accum_59__3_,prod_accum_59__2_,
  prod_accum_59__1_,prod_accum_59__0_,s_r_66__127_,s_r_66__126_,s_r_66__125_,s_r_66__124_,
  s_r_66__123_,s_r_66__122_,s_r_66__121_,s_r_66__120_,s_r_66__119_,s_r_66__118_,
  s_r_66__117_,s_r_66__116_,s_r_66__115_,s_r_66__114_,s_r_66__113_,s_r_66__112_,
  s_r_66__111_,s_r_66__110_,s_r_66__109_,s_r_66__108_,s_r_66__107_,s_r_66__106_,
  s_r_66__105_,s_r_66__104_,s_r_66__103_,s_r_66__102_,s_r_66__101_,s_r_66__100_,s_r_66__99_,
  s_r_66__98_,s_r_66__97_,s_r_66__96_,s_r_66__95_,s_r_66__94_,s_r_66__93_,
  s_r_66__92_,s_r_66__91_,s_r_66__90_,s_r_66__89_,s_r_66__88_,s_r_66__87_,s_r_66__86_,
  s_r_66__85_,s_r_66__84_,s_r_66__83_,s_r_66__82_,s_r_66__81_,s_r_66__80_,s_r_66__79_,
  s_r_66__78_,s_r_66__77_,s_r_66__76_,s_r_66__75_,s_r_66__74_,s_r_66__73_,
  s_r_66__72_,s_r_66__71_,s_r_66__70_,s_r_66__69_,s_r_66__68_,s_r_66__67_,s_r_66__66_,
  s_r_66__65_,s_r_66__64_,s_r_66__63_,s_r_66__62_,s_r_66__61_,s_r_66__60_,s_r_66__59_,
  s_r_66__58_,s_r_66__57_,s_r_66__56_,s_r_66__55_,s_r_66__54_,s_r_66__53_,
  s_r_66__52_,s_r_66__51_,s_r_66__50_,s_r_66__49_,s_r_66__48_,s_r_66__47_,s_r_66__46_,
  s_r_66__45_,s_r_66__44_,s_r_66__43_,s_r_66__42_,s_r_66__41_,s_r_66__40_,s_r_66__39_,
  s_r_66__38_,s_r_66__37_,s_r_66__36_,s_r_66__35_,s_r_66__34_,s_r_66__33_,
  s_r_66__32_,s_r_66__31_,s_r_66__30_,s_r_66__29_,s_r_66__28_,s_r_66__27_,s_r_66__26_,
  s_r_66__25_,s_r_66__24_,s_r_66__23_,s_r_66__22_,s_r_66__21_,s_r_66__20_,s_r_66__19_,
  s_r_66__18_,s_r_66__17_,s_r_66__16_,s_r_66__15_,s_r_66__14_,s_r_66__13_,
  s_r_66__12_,s_r_66__11_,s_r_66__10_,s_r_66__9_,s_r_66__8_,s_r_66__7_,s_r_66__6_,
  s_r_66__5_,s_r_66__4_,s_r_66__3_,s_r_66__2_,s_r_66__1_,s_r_66__0_,s_r_65__127_,
  s_r_65__126_,s_r_65__125_,s_r_65__124_,s_r_65__123_,s_r_65__122_,s_r_65__121_,
  s_r_65__120_,s_r_65__119_,s_r_65__118_,s_r_65__117_,s_r_65__116_,s_r_65__115_,s_r_65__114_,
  s_r_65__113_,s_r_65__112_,s_r_65__111_,s_r_65__110_,s_r_65__109_,s_r_65__108_,
  s_r_65__107_,s_r_65__106_,s_r_65__105_,s_r_65__104_,s_r_65__103_,s_r_65__102_,
  s_r_65__101_,s_r_65__100_,s_r_65__99_,s_r_65__98_,s_r_65__97_,s_r_65__96_,
  s_r_65__95_,s_r_65__94_,s_r_65__93_,s_r_65__92_,s_r_65__91_,s_r_65__90_,s_r_65__89_,
  s_r_65__88_,s_r_65__87_,s_r_65__86_,s_r_65__85_,s_r_65__84_,s_r_65__83_,s_r_65__82_,
  s_r_65__81_,s_r_65__80_,s_r_65__79_,s_r_65__78_,s_r_65__77_,s_r_65__76_,
  s_r_65__75_,s_r_65__74_,s_r_65__73_,s_r_65__72_,s_r_65__71_,s_r_65__70_,s_r_65__69_,
  s_r_65__68_,s_r_65__67_,s_r_65__66_,s_r_65__65_,s_r_65__64_,s_r_65__63_,s_r_65__62_,
  s_r_65__61_,s_r_65__60_,s_r_65__59_,s_r_65__58_,s_r_65__57_,s_r_65__56_,
  s_r_65__55_,s_r_65__54_,s_r_65__53_,s_r_65__52_,s_r_65__51_,s_r_65__50_,s_r_65__49_,
  s_r_65__48_,s_r_65__47_,s_r_65__46_,s_r_65__45_,s_r_65__44_,s_r_65__43_,s_r_65__42_,
  s_r_65__41_,s_r_65__40_,s_r_65__39_,s_r_65__38_,s_r_65__37_,s_r_65__36_,
  s_r_65__35_,s_r_65__34_,s_r_65__33_,s_r_65__32_,s_r_65__31_,s_r_65__30_,s_r_65__29_,
  s_r_65__28_,s_r_65__27_,s_r_65__26_,s_r_65__25_,s_r_65__24_,s_r_65__23_,s_r_65__22_,
  s_r_65__21_,s_r_65__20_,s_r_65__19_,s_r_65__18_,s_r_65__17_,s_r_65__16_,
  s_r_65__15_,s_r_65__14_,s_r_65__13_,s_r_65__12_,s_r_65__11_,s_r_65__10_,s_r_65__9_,
  s_r_65__8_,s_r_65__7_,s_r_65__6_,s_r_65__5_,s_r_65__4_,s_r_65__3_,s_r_65__2_,
  s_r_65__1_,s_r_65__0_,s_r_64__127_,s_r_64__126_,s_r_64__125_,s_r_64__124_,s_r_64__123_,
  s_r_64__122_,s_r_64__121_,s_r_64__120_,s_r_64__119_,s_r_64__118_,s_r_64__117_,
  s_r_64__116_,s_r_64__115_,s_r_64__114_,s_r_64__113_,s_r_64__112_,s_r_64__111_,
  s_r_64__110_,s_r_64__109_,s_r_64__108_,s_r_64__107_,s_r_64__106_,s_r_64__105_,
  s_r_64__104_,s_r_64__103_,s_r_64__102_,s_r_64__101_,s_r_64__100_,s_r_64__99_,s_r_64__98_,
  s_r_64__97_,s_r_64__96_,s_r_64__95_,s_r_64__94_,s_r_64__93_,s_r_64__92_,
  s_r_64__91_,s_r_64__90_,s_r_64__89_,s_r_64__88_,s_r_64__87_,s_r_64__86_,s_r_64__85_,
  s_r_64__84_,s_r_64__83_,s_r_64__82_,s_r_64__81_,s_r_64__80_,s_r_64__79_,s_r_64__78_,
  s_r_64__77_,s_r_64__76_,s_r_64__75_,s_r_64__74_,s_r_64__73_,s_r_64__72_,
  s_r_64__71_,s_r_64__70_,s_r_64__69_,s_r_64__68_,s_r_64__67_,s_r_64__66_,s_r_64__65_,
  s_r_64__64_,s_r_64__63_,s_r_64__62_,s_r_64__61_,s_r_64__60_,s_r_64__59_,s_r_64__58_,
  s_r_64__57_,s_r_64__56_,s_r_64__55_,s_r_64__54_,s_r_64__53_,s_r_64__52_,
  s_r_64__51_,s_r_64__50_,s_r_64__49_,s_r_64__48_,s_r_64__47_,s_r_64__46_,s_r_64__45_,
  s_r_64__44_,s_r_64__43_,s_r_64__42_,s_r_64__41_,s_r_64__40_,s_r_64__39_,s_r_64__38_,
  s_r_64__37_,s_r_64__36_,s_r_64__35_,s_r_64__34_,s_r_64__33_,s_r_64__32_,
  s_r_64__31_,s_r_64__30_,s_r_64__29_,s_r_64__28_,s_r_64__27_,s_r_64__26_,s_r_64__25_,
  s_r_64__24_,s_r_64__23_,s_r_64__22_,s_r_64__21_,s_r_64__20_,s_r_64__19_,s_r_64__18_,
  s_r_64__17_,s_r_64__16_,s_r_64__15_,s_r_64__14_,s_r_64__13_,s_r_64__12_,
  s_r_64__11_,s_r_64__10_,s_r_64__9_,s_r_64__8_,s_r_64__7_,s_r_64__6_,s_r_64__5_,
  s_r_64__4_,s_r_64__3_,s_r_64__2_,s_r_64__1_,s_r_64__0_,s_r_63__127_,s_r_63__126_,
  s_r_63__125_,s_r_63__124_,s_r_63__123_,s_r_63__122_,s_r_63__121_,s_r_63__120_,
  s_r_63__119_,s_r_63__118_,s_r_63__117_,s_r_63__116_,s_r_63__115_,s_r_63__114_,
  s_r_63__113_,s_r_63__112_,s_r_63__111_,s_r_63__110_,s_r_63__109_,s_r_63__108_,s_r_63__107_,
  s_r_63__106_,s_r_63__105_,s_r_63__104_,s_r_63__103_,s_r_63__102_,s_r_63__101_,
  s_r_63__100_,s_r_63__99_,s_r_63__98_,s_r_63__97_,s_r_63__96_,s_r_63__95_,
  s_r_63__94_,s_r_63__93_,s_r_63__92_,s_r_63__91_,s_r_63__90_,s_r_63__89_,s_r_63__88_,
  s_r_63__87_,s_r_63__86_,s_r_63__85_,s_r_63__84_,s_r_63__83_,s_r_63__82_,s_r_63__81_,
  s_r_63__80_,s_r_63__79_,s_r_63__78_,s_r_63__77_,s_r_63__76_,s_r_63__75_,
  s_r_63__74_,s_r_63__73_,s_r_63__72_,s_r_63__71_,s_r_63__70_,s_r_63__69_,s_r_63__68_,
  s_r_63__67_,s_r_63__66_,s_r_63__65_,s_r_63__64_,s_r_63__63_,s_r_63__62_,s_r_63__61_,
  s_r_63__60_,s_r_63__59_,s_r_63__58_,s_r_63__57_,s_r_63__56_,s_r_63__55_,
  s_r_63__54_,s_r_63__53_,s_r_63__52_,s_r_63__51_,s_r_63__50_,s_r_63__49_,s_r_63__48_,
  s_r_63__47_,s_r_63__46_,s_r_63__45_,s_r_63__44_,s_r_63__43_,s_r_63__42_,s_r_63__41_,
  s_r_63__40_,s_r_63__39_,s_r_63__38_,s_r_63__37_,s_r_63__36_,s_r_63__35_,
  s_r_63__34_,s_r_63__33_,s_r_63__32_,s_r_63__31_,s_r_63__30_,s_r_63__29_,s_r_63__28_,
  s_r_63__27_,s_r_63__26_,s_r_63__25_,s_r_63__24_,s_r_63__23_,s_r_63__22_,s_r_63__21_,
  s_r_63__20_,s_r_63__19_,s_r_63__18_,s_r_63__17_,s_r_63__16_,s_r_63__15_,
  s_r_63__14_,s_r_63__13_,s_r_63__12_,s_r_63__11_,s_r_63__10_,s_r_63__9_,s_r_63__8_,
  s_r_63__7_,s_r_63__6_,s_r_63__5_,s_r_63__4_,s_r_63__3_,s_r_63__2_,s_r_63__1_,s_r_63__0_,
  prod_accum_66__67_,prod_accum_66__66_,prod_accum_66__65_,prod_accum_66__64_,
  prod_accum_66__63_,prod_accum_66__62_,prod_accum_66__61_,prod_accum_66__60_,
  prod_accum_66__59_,prod_accum_66__58_,prod_accum_66__57_,prod_accum_66__56_,
  prod_accum_66__55_,prod_accum_66__54_,prod_accum_66__53_,prod_accum_66__52_,
  prod_accum_66__51_,prod_accum_66__50_,prod_accum_66__49_,prod_accum_66__48_,prod_accum_66__47_,
  prod_accum_66__46_,prod_accum_66__45_,prod_accum_66__44_,prod_accum_66__43_,
  prod_accum_66__42_,prod_accum_66__41_,prod_accum_66__40_,prod_accum_66__39_,
  prod_accum_66__38_,prod_accum_66__37_,prod_accum_66__36_,prod_accum_66__35_,
  prod_accum_66__34_,prod_accum_66__33_,prod_accum_66__32_,prod_accum_66__31_,
  prod_accum_66__30_,prod_accum_66__29_,prod_accum_66__28_,prod_accum_66__27_,prod_accum_66__26_,
  prod_accum_66__25_,prod_accum_66__24_,prod_accum_66__23_,prod_accum_66__22_,
  prod_accum_66__21_,prod_accum_66__20_,prod_accum_66__19_,prod_accum_66__18_,
  prod_accum_66__17_,prod_accum_66__16_,prod_accum_66__15_,prod_accum_66__14_,
  prod_accum_66__13_,prod_accum_66__12_,prod_accum_66__11_,prod_accum_66__10_,prod_accum_66__9_,
  prod_accum_66__8_,prod_accum_66__7_,prod_accum_66__6_,prod_accum_66__5_,
  prod_accum_66__4_,prod_accum_66__3_,prod_accum_66__2_,prod_accum_66__1_,
  prod_accum_66__0_,prod_accum_65__66_,prod_accum_65__65_,prod_accum_65__64_,prod_accum_65__63_,
  prod_accum_65__62_,prod_accum_65__61_,prod_accum_65__60_,prod_accum_65__59_,
  prod_accum_65__58_,prod_accum_65__57_,prod_accum_65__56_,prod_accum_65__55_,
  prod_accum_65__54_,prod_accum_65__53_,prod_accum_65__52_,prod_accum_65__51_,
  prod_accum_65__50_,prod_accum_65__49_,prod_accum_65__48_,prod_accum_65__47_,
  prod_accum_65__46_,prod_accum_65__45_,prod_accum_65__44_,prod_accum_65__43_,prod_accum_65__42_,
  prod_accum_65__41_,prod_accum_65__40_,prod_accum_65__39_,prod_accum_65__38_,
  prod_accum_65__37_,prod_accum_65__36_,prod_accum_65__35_,prod_accum_65__34_,
  prod_accum_65__33_,prod_accum_65__32_,prod_accum_65__31_,prod_accum_65__30_,
  prod_accum_65__29_,prod_accum_65__28_,prod_accum_65__27_,prod_accum_65__26_,prod_accum_65__25_,
  prod_accum_65__24_,prod_accum_65__23_,prod_accum_65__22_,prod_accum_65__21_,
  prod_accum_65__20_,prod_accum_65__19_,prod_accum_65__18_,prod_accum_65__17_,
  prod_accum_65__16_,prod_accum_65__15_,prod_accum_65__14_,prod_accum_65__13_,
  prod_accum_65__12_,prod_accum_65__11_,prod_accum_65__10_,prod_accum_65__9_,
  prod_accum_65__8_,prod_accum_65__7_,prod_accum_65__6_,prod_accum_65__5_,prod_accum_65__4_,
  prod_accum_65__3_,prod_accum_65__2_,prod_accum_65__1_,prod_accum_65__0_,
  prod_accum_64__65_,prod_accum_64__64_,prod_accum_64__63_,prod_accum_64__62_,prod_accum_64__61_,
  prod_accum_64__60_,prod_accum_64__59_,prod_accum_64__58_,prod_accum_64__57_,
  prod_accum_64__56_,prod_accum_64__55_,prod_accum_64__54_,prod_accum_64__53_,
  prod_accum_64__52_,prod_accum_64__51_,prod_accum_64__50_,prod_accum_64__49_,
  prod_accum_64__48_,prod_accum_64__47_,prod_accum_64__46_,prod_accum_64__45_,
  prod_accum_64__44_,prod_accum_64__43_,prod_accum_64__42_,prod_accum_64__41_,prod_accum_64__40_,
  prod_accum_64__39_,prod_accum_64__38_,prod_accum_64__37_,prod_accum_64__36_,
  prod_accum_64__35_,prod_accum_64__34_,prod_accum_64__33_,prod_accum_64__32_,
  prod_accum_64__31_,prod_accum_64__30_,prod_accum_64__29_,prod_accum_64__28_,
  prod_accum_64__27_,prod_accum_64__26_,prod_accum_64__25_,prod_accum_64__24_,
  prod_accum_64__23_,prod_accum_64__22_,prod_accum_64__21_,prod_accum_64__20_,prod_accum_64__19_,
  prod_accum_64__18_,prod_accum_64__17_,prod_accum_64__16_,prod_accum_64__15_,
  prod_accum_64__14_,prod_accum_64__13_,prod_accum_64__12_,prod_accum_64__11_,
  prod_accum_64__10_,prod_accum_64__9_,prod_accum_64__8_,prod_accum_64__7_,
  prod_accum_64__6_,prod_accum_64__5_,prod_accum_64__4_,prod_accum_64__3_,prod_accum_64__2_,
  prod_accum_64__1_,prod_accum_64__0_,prod_accum_63__64_,prod_accum_63__63_,
  prod_accum_63__62_,prod_accum_63__61_,prod_accum_63__60_,prod_accum_63__59_,
  prod_accum_63__58_,prod_accum_63__57_,prod_accum_63__56_,prod_accum_63__55_,prod_accum_63__54_,
  prod_accum_63__53_,prod_accum_63__52_,prod_accum_63__51_,prod_accum_63__50_,
  prod_accum_63__49_,prod_accum_63__48_,prod_accum_63__47_,prod_accum_63__46_,
  prod_accum_63__45_,prod_accum_63__44_,prod_accum_63__43_,prod_accum_63__42_,
  prod_accum_63__41_,prod_accum_63__40_,prod_accum_63__39_,prod_accum_63__38_,
  prod_accum_63__37_,prod_accum_63__36_,prod_accum_63__35_,prod_accum_63__34_,prod_accum_63__33_,
  prod_accum_63__32_,prod_accum_63__31_,prod_accum_63__30_,prod_accum_63__29_,
  prod_accum_63__28_,prod_accum_63__27_,prod_accum_63__26_,prod_accum_63__25_,
  prod_accum_63__24_,prod_accum_63__23_,prod_accum_63__22_,prod_accum_63__21_,
  prod_accum_63__20_,prod_accum_63__19_,prod_accum_63__18_,prod_accum_63__17_,prod_accum_63__16_,
  prod_accum_63__15_,prod_accum_63__14_,prod_accum_63__13_,prod_accum_63__12_,
  prod_accum_63__11_,prod_accum_63__10_,prod_accum_63__9_,prod_accum_63__8_,
  prod_accum_63__7_,prod_accum_63__6_,prod_accum_63__5_,prod_accum_63__4_,prod_accum_63__3_,
  prod_accum_63__2_,prod_accum_63__1_,prod_accum_63__0_,s_r_70__127_,s_r_70__126_,
  s_r_70__125_,s_r_70__124_,s_r_70__123_,s_r_70__122_,s_r_70__121_,s_r_70__120_,
  s_r_70__119_,s_r_70__118_,s_r_70__117_,s_r_70__116_,s_r_70__115_,s_r_70__114_,
  s_r_70__113_,s_r_70__112_,s_r_70__111_,s_r_70__110_,s_r_70__109_,s_r_70__108_,
  s_r_70__107_,s_r_70__106_,s_r_70__105_,s_r_70__104_,s_r_70__103_,s_r_70__102_,
  s_r_70__101_,s_r_70__100_,s_r_70__99_,s_r_70__98_,s_r_70__97_,s_r_70__96_,s_r_70__95_,
  s_r_70__94_,s_r_70__93_,s_r_70__92_,s_r_70__91_,s_r_70__90_,s_r_70__89_,
  s_r_70__88_,s_r_70__87_,s_r_70__86_,s_r_70__85_,s_r_70__84_,s_r_70__83_,s_r_70__82_,
  s_r_70__81_,s_r_70__80_,s_r_70__79_,s_r_70__78_,s_r_70__77_,s_r_70__76_,s_r_70__75_,
  s_r_70__74_,s_r_70__73_,s_r_70__72_,s_r_70__71_,s_r_70__70_,s_r_70__69_,
  s_r_70__68_,s_r_70__67_,s_r_70__66_,s_r_70__65_,s_r_70__64_,s_r_70__63_,s_r_70__62_,
  s_r_70__61_,s_r_70__60_,s_r_70__59_,s_r_70__58_,s_r_70__57_,s_r_70__56_,s_r_70__55_,
  s_r_70__54_,s_r_70__53_,s_r_70__52_,s_r_70__51_,s_r_70__50_,s_r_70__49_,
  s_r_70__48_,s_r_70__47_,s_r_70__46_,s_r_70__45_,s_r_70__44_,s_r_70__43_,s_r_70__42_,
  s_r_70__41_,s_r_70__40_,s_r_70__39_,s_r_70__38_,s_r_70__37_,s_r_70__36_,s_r_70__35_,
  s_r_70__34_,s_r_70__33_,s_r_70__32_,s_r_70__31_,s_r_70__30_,s_r_70__29_,
  s_r_70__28_,s_r_70__27_,s_r_70__26_,s_r_70__25_,s_r_70__24_,s_r_70__23_,s_r_70__22_,
  s_r_70__21_,s_r_70__20_,s_r_70__19_,s_r_70__18_,s_r_70__17_,s_r_70__16_,s_r_70__15_,
  s_r_70__14_,s_r_70__13_,s_r_70__12_,s_r_70__11_,s_r_70__10_,s_r_70__9_,s_r_70__8_,
  s_r_70__7_,s_r_70__6_,s_r_70__5_,s_r_70__4_,s_r_70__3_,s_r_70__2_,s_r_70__1_,
  s_r_70__0_,s_r_69__127_,s_r_69__126_,s_r_69__125_,s_r_69__124_,s_r_69__123_,
  s_r_69__122_,s_r_69__121_,s_r_69__120_,s_r_69__119_,s_r_69__118_,s_r_69__117_,
  s_r_69__116_,s_r_69__115_,s_r_69__114_,s_r_69__113_,s_r_69__112_,s_r_69__111_,
  s_r_69__110_,s_r_69__109_,s_r_69__108_,s_r_69__107_,s_r_69__106_,s_r_69__105_,s_r_69__104_,
  s_r_69__103_,s_r_69__102_,s_r_69__101_,s_r_69__100_,s_r_69__99_,s_r_69__98_,
  s_r_69__97_,s_r_69__96_,s_r_69__95_,s_r_69__94_,s_r_69__93_,s_r_69__92_,s_r_69__91_,
  s_r_69__90_,s_r_69__89_,s_r_69__88_,s_r_69__87_,s_r_69__86_,s_r_69__85_,
  s_r_69__84_,s_r_69__83_,s_r_69__82_,s_r_69__81_,s_r_69__80_,s_r_69__79_,s_r_69__78_,
  s_r_69__77_,s_r_69__76_,s_r_69__75_,s_r_69__74_,s_r_69__73_,s_r_69__72_,s_r_69__71_,
  s_r_69__70_,s_r_69__69_,s_r_69__68_,s_r_69__67_,s_r_69__66_,s_r_69__65_,
  s_r_69__64_,s_r_69__63_,s_r_69__62_,s_r_69__61_,s_r_69__60_,s_r_69__59_,s_r_69__58_,
  s_r_69__57_,s_r_69__56_,s_r_69__55_,s_r_69__54_,s_r_69__53_,s_r_69__52_,s_r_69__51_,
  s_r_69__50_,s_r_69__49_,s_r_69__48_,s_r_69__47_,s_r_69__46_,s_r_69__45_,
  s_r_69__44_,s_r_69__43_,s_r_69__42_,s_r_69__41_,s_r_69__40_,s_r_69__39_,s_r_69__38_,
  s_r_69__37_,s_r_69__36_,s_r_69__35_,s_r_69__34_,s_r_69__33_,s_r_69__32_,s_r_69__31_,
  s_r_69__30_,s_r_69__29_,s_r_69__28_,s_r_69__27_,s_r_69__26_,s_r_69__25_,
  s_r_69__24_,s_r_69__23_,s_r_69__22_,s_r_69__21_,s_r_69__20_,s_r_69__19_,s_r_69__18_,
  s_r_69__17_,s_r_69__16_,s_r_69__15_,s_r_69__14_,s_r_69__13_,s_r_69__12_,s_r_69__11_,
  s_r_69__10_,s_r_69__9_,s_r_69__8_,s_r_69__7_,s_r_69__6_,s_r_69__5_,s_r_69__4_,
  s_r_69__3_,s_r_69__2_,s_r_69__1_,s_r_69__0_,s_r_68__127_,s_r_68__126_,
  s_r_68__125_,s_r_68__124_,s_r_68__123_,s_r_68__122_,s_r_68__121_,s_r_68__120_,s_r_68__119_,
  s_r_68__118_,s_r_68__117_,s_r_68__116_,s_r_68__115_,s_r_68__114_,s_r_68__113_,
  s_r_68__112_,s_r_68__111_,s_r_68__110_,s_r_68__109_,s_r_68__108_,s_r_68__107_,
  s_r_68__106_,s_r_68__105_,s_r_68__104_,s_r_68__103_,s_r_68__102_,s_r_68__101_,
  s_r_68__100_,s_r_68__99_,s_r_68__98_,s_r_68__97_,s_r_68__96_,s_r_68__95_,s_r_68__94_,
  s_r_68__93_,s_r_68__92_,s_r_68__91_,s_r_68__90_,s_r_68__89_,s_r_68__88_,
  s_r_68__87_,s_r_68__86_,s_r_68__85_,s_r_68__84_,s_r_68__83_,s_r_68__82_,s_r_68__81_,
  s_r_68__80_,s_r_68__79_,s_r_68__78_,s_r_68__77_,s_r_68__76_,s_r_68__75_,s_r_68__74_,
  s_r_68__73_,s_r_68__72_,s_r_68__71_,s_r_68__70_,s_r_68__69_,s_r_68__68_,
  s_r_68__67_,s_r_68__66_,s_r_68__65_,s_r_68__64_,s_r_68__63_,s_r_68__62_,s_r_68__61_,
  s_r_68__60_,s_r_68__59_,s_r_68__58_,s_r_68__57_,s_r_68__56_,s_r_68__55_,s_r_68__54_,
  s_r_68__53_,s_r_68__52_,s_r_68__51_,s_r_68__50_,s_r_68__49_,s_r_68__48_,
  s_r_68__47_,s_r_68__46_,s_r_68__45_,s_r_68__44_,s_r_68__43_,s_r_68__42_,s_r_68__41_,
  s_r_68__40_,s_r_68__39_,s_r_68__38_,s_r_68__37_,s_r_68__36_,s_r_68__35_,s_r_68__34_,
  s_r_68__33_,s_r_68__32_,s_r_68__31_,s_r_68__30_,s_r_68__29_,s_r_68__28_,
  s_r_68__27_,s_r_68__26_,s_r_68__25_,s_r_68__24_,s_r_68__23_,s_r_68__22_,s_r_68__21_,
  s_r_68__20_,s_r_68__19_,s_r_68__18_,s_r_68__17_,s_r_68__16_,s_r_68__15_,s_r_68__14_,
  s_r_68__13_,s_r_68__12_,s_r_68__11_,s_r_68__10_,s_r_68__9_,s_r_68__8_,s_r_68__7_,
  s_r_68__6_,s_r_68__5_,s_r_68__4_,s_r_68__3_,s_r_68__2_,s_r_68__1_,s_r_68__0_,
  s_r_67__127_,s_r_67__126_,s_r_67__125_,s_r_67__124_,s_r_67__123_,s_r_67__122_,
  s_r_67__121_,s_r_67__120_,s_r_67__119_,s_r_67__118_,s_r_67__117_,s_r_67__116_,
  s_r_67__115_,s_r_67__114_,s_r_67__113_,s_r_67__112_,s_r_67__111_,s_r_67__110_,
  s_r_67__109_,s_r_67__108_,s_r_67__107_,s_r_67__106_,s_r_67__105_,s_r_67__104_,
  s_r_67__103_,s_r_67__102_,s_r_67__101_,s_r_67__100_,s_r_67__99_,s_r_67__98_,s_r_67__97_,
  s_r_67__96_,s_r_67__95_,s_r_67__94_,s_r_67__93_,s_r_67__92_,s_r_67__91_,s_r_67__90_,
  s_r_67__89_,s_r_67__88_,s_r_67__87_,s_r_67__86_,s_r_67__85_,s_r_67__84_,
  s_r_67__83_,s_r_67__82_,s_r_67__81_,s_r_67__80_,s_r_67__79_,s_r_67__78_,s_r_67__77_,
  s_r_67__76_,s_r_67__75_,s_r_67__74_,s_r_67__73_,s_r_67__72_,s_r_67__71_,s_r_67__70_,
  s_r_67__69_,s_r_67__68_,s_r_67__67_,s_r_67__66_,s_r_67__65_,s_r_67__64_,
  s_r_67__63_,s_r_67__62_,s_r_67__61_,s_r_67__60_,s_r_67__59_,s_r_67__58_,s_r_67__57_,
  s_r_67__56_,s_r_67__55_,s_r_67__54_,s_r_67__53_,s_r_67__52_,s_r_67__51_,s_r_67__50_,
  s_r_67__49_,s_r_67__48_,s_r_67__47_,s_r_67__46_,s_r_67__45_,s_r_67__44_,
  s_r_67__43_,s_r_67__42_,s_r_67__41_,s_r_67__40_,s_r_67__39_,s_r_67__38_,s_r_67__37_,
  s_r_67__36_,s_r_67__35_,s_r_67__34_,s_r_67__33_,s_r_67__32_,s_r_67__31_,s_r_67__30_,
  s_r_67__29_,s_r_67__28_,s_r_67__27_,s_r_67__26_,s_r_67__25_,s_r_67__24_,
  s_r_67__23_,s_r_67__22_,s_r_67__21_,s_r_67__20_,s_r_67__19_,s_r_67__18_,s_r_67__17_,
  s_r_67__16_,s_r_67__15_,s_r_67__14_,s_r_67__13_,s_r_67__12_,s_r_67__11_,s_r_67__10_,
  s_r_67__9_,s_r_67__8_,s_r_67__7_,s_r_67__6_,s_r_67__5_,s_r_67__4_,s_r_67__3_,
  s_r_67__2_,s_r_67__1_,s_r_67__0_,prod_accum_70__71_,prod_accum_70__70_,
  prod_accum_70__69_,prod_accum_70__68_,prod_accum_70__67_,prod_accum_70__66_,
  prod_accum_70__65_,prod_accum_70__64_,prod_accum_70__63_,prod_accum_70__62_,prod_accum_70__61_,
  prod_accum_70__60_,prod_accum_70__59_,prod_accum_70__58_,prod_accum_70__57_,
  prod_accum_70__56_,prod_accum_70__55_,prod_accum_70__54_,prod_accum_70__53_,
  prod_accum_70__52_,prod_accum_70__51_,prod_accum_70__50_,prod_accum_70__49_,
  prod_accum_70__48_,prod_accum_70__47_,prod_accum_70__46_,prod_accum_70__45_,
  prod_accum_70__44_,prod_accum_70__43_,prod_accum_70__42_,prod_accum_70__41_,prod_accum_70__40_,
  prod_accum_70__39_,prod_accum_70__38_,prod_accum_70__37_,prod_accum_70__36_,
  prod_accum_70__35_,prod_accum_70__34_,prod_accum_70__33_,prod_accum_70__32_,
  prod_accum_70__31_,prod_accum_70__30_,prod_accum_70__29_,prod_accum_70__28_,
  prod_accum_70__27_,prod_accum_70__26_,prod_accum_70__25_,prod_accum_70__24_,
  prod_accum_70__23_,prod_accum_70__22_,prod_accum_70__21_,prod_accum_70__20_,prod_accum_70__19_,
  prod_accum_70__18_,prod_accum_70__17_,prod_accum_70__16_,prod_accum_70__15_,
  prod_accum_70__14_,prod_accum_70__13_,prod_accum_70__12_,prod_accum_70__11_,
  prod_accum_70__10_,prod_accum_70__9_,prod_accum_70__8_,prod_accum_70__7_,prod_accum_70__6_,
  prod_accum_70__5_,prod_accum_70__4_,prod_accum_70__3_,prod_accum_70__2_,
  prod_accum_70__1_,prod_accum_70__0_,prod_accum_69__70_,prod_accum_69__69_,
  prod_accum_69__68_,prod_accum_69__67_,prod_accum_69__66_,prod_accum_69__65_,
  prod_accum_69__64_,prod_accum_69__63_,prod_accum_69__62_,prod_accum_69__61_,prod_accum_69__60_,
  prod_accum_69__59_,prod_accum_69__58_,prod_accum_69__57_,prod_accum_69__56_,
  prod_accum_69__55_,prod_accum_69__54_,prod_accum_69__53_,prod_accum_69__52_,
  prod_accum_69__51_,prod_accum_69__50_,prod_accum_69__49_,prod_accum_69__48_,
  prod_accum_69__47_,prod_accum_69__46_,prod_accum_69__45_,prod_accum_69__44_,prod_accum_69__43_,
  prod_accum_69__42_,prod_accum_69__41_,prod_accum_69__40_,prod_accum_69__39_,
  prod_accum_69__38_,prod_accum_69__37_,prod_accum_69__36_,prod_accum_69__35_,
  prod_accum_69__34_,prod_accum_69__33_,prod_accum_69__32_,prod_accum_69__31_,
  prod_accum_69__30_,prod_accum_69__29_,prod_accum_69__28_,prod_accum_69__27_,
  prod_accum_69__26_,prod_accum_69__25_,prod_accum_69__24_,prod_accum_69__23_,prod_accum_69__22_,
  prod_accum_69__21_,prod_accum_69__20_,prod_accum_69__19_,prod_accum_69__18_,
  prod_accum_69__17_,prod_accum_69__16_,prod_accum_69__15_,prod_accum_69__14_,
  prod_accum_69__13_,prod_accum_69__12_,prod_accum_69__11_,prod_accum_69__10_,
  prod_accum_69__9_,prod_accum_69__8_,prod_accum_69__7_,prod_accum_69__6_,prod_accum_69__5_,
  prod_accum_69__4_,prod_accum_69__3_,prod_accum_69__2_,prod_accum_69__1_,
  prod_accum_69__0_,prod_accum_68__69_,prod_accum_68__68_,prod_accum_68__67_,
  prod_accum_68__66_,prod_accum_68__65_,prod_accum_68__64_,prod_accum_68__63_,prod_accum_68__62_,
  prod_accum_68__61_,prod_accum_68__60_,prod_accum_68__59_,prod_accum_68__58_,
  prod_accum_68__57_,prod_accum_68__56_,prod_accum_68__55_,prod_accum_68__54_,
  prod_accum_68__53_,prod_accum_68__52_,prod_accum_68__51_,prod_accum_68__50_,
  prod_accum_68__49_,prod_accum_68__48_,prod_accum_68__47_,prod_accum_68__46_,
  prod_accum_68__45_,prod_accum_68__44_,prod_accum_68__43_,prod_accum_68__42_,prod_accum_68__41_,
  prod_accum_68__40_,prod_accum_68__39_,prod_accum_68__38_,prod_accum_68__37_,
  prod_accum_68__36_,prod_accum_68__35_,prod_accum_68__34_,prod_accum_68__33_,
  prod_accum_68__32_,prod_accum_68__31_,prod_accum_68__30_,prod_accum_68__29_,
  prod_accum_68__28_,prod_accum_68__27_,prod_accum_68__26_,prod_accum_68__25_,
  prod_accum_68__24_,prod_accum_68__23_,prod_accum_68__22_,prod_accum_68__21_,prod_accum_68__20_,
  prod_accum_68__19_,prod_accum_68__18_,prod_accum_68__17_,prod_accum_68__16_,
  prod_accum_68__15_,prod_accum_68__14_,prod_accum_68__13_,prod_accum_68__12_,
  prod_accum_68__11_,prod_accum_68__10_,prod_accum_68__9_,prod_accum_68__8_,
  prod_accum_68__7_,prod_accum_68__6_,prod_accum_68__5_,prod_accum_68__4_,prod_accum_68__3_,
  prod_accum_68__2_,prod_accum_68__1_,prod_accum_68__0_,prod_accum_67__68_,
  prod_accum_67__67_,prod_accum_67__66_,prod_accum_67__65_,prod_accum_67__64_,
  prod_accum_67__63_,prod_accum_67__62_,prod_accum_67__61_,prod_accum_67__60_,prod_accum_67__59_,
  prod_accum_67__58_,prod_accum_67__57_,prod_accum_67__56_,prod_accum_67__55_,
  prod_accum_67__54_,prod_accum_67__53_,prod_accum_67__52_,prod_accum_67__51_,
  prod_accum_67__50_,prod_accum_67__49_,prod_accum_67__48_,prod_accum_67__47_,
  prod_accum_67__46_,prod_accum_67__45_,prod_accum_67__44_,prod_accum_67__43_,prod_accum_67__42_,
  prod_accum_67__41_,prod_accum_67__40_,prod_accum_67__39_,prod_accum_67__38_,
  prod_accum_67__37_,prod_accum_67__36_,prod_accum_67__35_,prod_accum_67__34_,
  prod_accum_67__33_,prod_accum_67__32_,prod_accum_67__31_,prod_accum_67__30_,
  prod_accum_67__29_,prod_accum_67__28_,prod_accum_67__27_,prod_accum_67__26_,
  prod_accum_67__25_,prod_accum_67__24_,prod_accum_67__23_,prod_accum_67__22_,prod_accum_67__21_,
  prod_accum_67__20_,prod_accum_67__19_,prod_accum_67__18_,prod_accum_67__17_,
  prod_accum_67__16_,prod_accum_67__15_,prod_accum_67__14_,prod_accum_67__13_,
  prod_accum_67__12_,prod_accum_67__11_,prod_accum_67__10_,prod_accum_67__9_,
  prod_accum_67__8_,prod_accum_67__7_,prod_accum_67__6_,prod_accum_67__5_,prod_accum_67__4_,
  prod_accum_67__3_,prod_accum_67__2_,prod_accum_67__1_,prod_accum_67__0_,
  s_r_74__127_,s_r_74__126_,s_r_74__125_,s_r_74__124_,s_r_74__123_,s_r_74__122_,s_r_74__121_,
  s_r_74__120_,s_r_74__119_,s_r_74__118_,s_r_74__117_,s_r_74__116_,s_r_74__115_,
  s_r_74__114_,s_r_74__113_,s_r_74__112_,s_r_74__111_,s_r_74__110_,s_r_74__109_,
  s_r_74__108_,s_r_74__107_,s_r_74__106_,s_r_74__105_,s_r_74__104_,s_r_74__103_,
  s_r_74__102_,s_r_74__101_,s_r_74__100_,s_r_74__99_,s_r_74__98_,s_r_74__97_,s_r_74__96_,
  s_r_74__95_,s_r_74__94_,s_r_74__93_,s_r_74__92_,s_r_74__91_,s_r_74__90_,
  s_r_74__89_,s_r_74__88_,s_r_74__87_,s_r_74__86_,s_r_74__85_,s_r_74__84_,s_r_74__83_,
  s_r_74__82_,s_r_74__81_,s_r_74__80_,s_r_74__79_,s_r_74__78_,s_r_74__77_,s_r_74__76_,
  s_r_74__75_,s_r_74__74_,s_r_74__73_,s_r_74__72_,s_r_74__71_,s_r_74__70_,
  s_r_74__69_,s_r_74__68_,s_r_74__67_,s_r_74__66_,s_r_74__65_,s_r_74__64_,s_r_74__63_,
  s_r_74__62_,s_r_74__61_,s_r_74__60_,s_r_74__59_,s_r_74__58_,s_r_74__57_,s_r_74__56_,
  s_r_74__55_,s_r_74__54_,s_r_74__53_,s_r_74__52_,s_r_74__51_,s_r_74__50_,
  s_r_74__49_,s_r_74__48_,s_r_74__47_,s_r_74__46_,s_r_74__45_,s_r_74__44_,s_r_74__43_,
  s_r_74__42_,s_r_74__41_,s_r_74__40_,s_r_74__39_,s_r_74__38_,s_r_74__37_,s_r_74__36_,
  s_r_74__35_,s_r_74__34_,s_r_74__33_,s_r_74__32_,s_r_74__31_,s_r_74__30_,
  s_r_74__29_,s_r_74__28_,s_r_74__27_,s_r_74__26_,s_r_74__25_,s_r_74__24_,s_r_74__23_,
  s_r_74__22_,s_r_74__21_,s_r_74__20_,s_r_74__19_,s_r_74__18_,s_r_74__17_,s_r_74__16_,
  s_r_74__15_,s_r_74__14_,s_r_74__13_,s_r_74__12_,s_r_74__11_,s_r_74__10_,
  s_r_74__9_,s_r_74__8_,s_r_74__7_,s_r_74__6_,s_r_74__5_,s_r_74__4_,s_r_74__3_,s_r_74__2_,
  s_r_74__1_,s_r_74__0_,s_r_73__127_,s_r_73__126_,s_r_73__125_,s_r_73__124_,
  s_r_73__123_,s_r_73__122_,s_r_73__121_,s_r_73__120_,s_r_73__119_,s_r_73__118_,
  s_r_73__117_,s_r_73__116_,s_r_73__115_,s_r_73__114_,s_r_73__113_,s_r_73__112_,
  s_r_73__111_,s_r_73__110_,s_r_73__109_,s_r_73__108_,s_r_73__107_,s_r_73__106_,
  s_r_73__105_,s_r_73__104_,s_r_73__103_,s_r_73__102_,s_r_73__101_,s_r_73__100_,s_r_73__99_,
  s_r_73__98_,s_r_73__97_,s_r_73__96_,s_r_73__95_,s_r_73__94_,s_r_73__93_,
  s_r_73__92_,s_r_73__91_,s_r_73__90_,s_r_73__89_,s_r_73__88_,s_r_73__87_,s_r_73__86_,
  s_r_73__85_,s_r_73__84_,s_r_73__83_,s_r_73__82_,s_r_73__81_,s_r_73__80_,s_r_73__79_,
  s_r_73__78_,s_r_73__77_,s_r_73__76_,s_r_73__75_,s_r_73__74_,s_r_73__73_,
  s_r_73__72_,s_r_73__71_,s_r_73__70_,s_r_73__69_,s_r_73__68_,s_r_73__67_,s_r_73__66_,
  s_r_73__65_,s_r_73__64_,s_r_73__63_,s_r_73__62_,s_r_73__61_,s_r_73__60_,s_r_73__59_,
  s_r_73__58_,s_r_73__57_,s_r_73__56_,s_r_73__55_,s_r_73__54_,s_r_73__53_,
  s_r_73__52_,s_r_73__51_,s_r_73__50_,s_r_73__49_,s_r_73__48_,s_r_73__47_,s_r_73__46_,
  s_r_73__45_,s_r_73__44_,s_r_73__43_,s_r_73__42_,s_r_73__41_,s_r_73__40_,s_r_73__39_,
  s_r_73__38_,s_r_73__37_,s_r_73__36_,s_r_73__35_,s_r_73__34_,s_r_73__33_,
  s_r_73__32_,s_r_73__31_,s_r_73__30_,s_r_73__29_,s_r_73__28_,s_r_73__27_,s_r_73__26_,
  s_r_73__25_,s_r_73__24_,s_r_73__23_,s_r_73__22_,s_r_73__21_,s_r_73__20_,s_r_73__19_,
  s_r_73__18_,s_r_73__17_,s_r_73__16_,s_r_73__15_,s_r_73__14_,s_r_73__13_,
  s_r_73__12_,s_r_73__11_,s_r_73__10_,s_r_73__9_,s_r_73__8_,s_r_73__7_,s_r_73__6_,
  s_r_73__5_,s_r_73__4_,s_r_73__3_,s_r_73__2_,s_r_73__1_,s_r_73__0_,s_r_72__127_,
  s_r_72__126_,s_r_72__125_,s_r_72__124_,s_r_72__123_,s_r_72__122_,s_r_72__121_,s_r_72__120_,
  s_r_72__119_,s_r_72__118_,s_r_72__117_,s_r_72__116_,s_r_72__115_,s_r_72__114_,
  s_r_72__113_,s_r_72__112_,s_r_72__111_,s_r_72__110_,s_r_72__109_,s_r_72__108_,
  s_r_72__107_,s_r_72__106_,s_r_72__105_,s_r_72__104_,s_r_72__103_,s_r_72__102_,
  s_r_72__101_,s_r_72__100_,s_r_72__99_,s_r_72__98_,s_r_72__97_,s_r_72__96_,s_r_72__95_,
  s_r_72__94_,s_r_72__93_,s_r_72__92_,s_r_72__91_,s_r_72__90_,s_r_72__89_,
  s_r_72__88_,s_r_72__87_,s_r_72__86_,s_r_72__85_,s_r_72__84_,s_r_72__83_,s_r_72__82_,
  s_r_72__81_,s_r_72__80_,s_r_72__79_,s_r_72__78_,s_r_72__77_,s_r_72__76_,s_r_72__75_,
  s_r_72__74_,s_r_72__73_,s_r_72__72_,s_r_72__71_,s_r_72__70_,s_r_72__69_,
  s_r_72__68_,s_r_72__67_,s_r_72__66_,s_r_72__65_,s_r_72__64_,s_r_72__63_,s_r_72__62_,
  s_r_72__61_,s_r_72__60_,s_r_72__59_,s_r_72__58_,s_r_72__57_,s_r_72__56_,s_r_72__55_,
  s_r_72__54_,s_r_72__53_,s_r_72__52_,s_r_72__51_,s_r_72__50_,s_r_72__49_,
  s_r_72__48_,s_r_72__47_,s_r_72__46_,s_r_72__45_,s_r_72__44_,s_r_72__43_,s_r_72__42_,
  s_r_72__41_,s_r_72__40_,s_r_72__39_,s_r_72__38_,s_r_72__37_,s_r_72__36_,s_r_72__35_,
  s_r_72__34_,s_r_72__33_,s_r_72__32_,s_r_72__31_,s_r_72__30_,s_r_72__29_,
  s_r_72__28_,s_r_72__27_,s_r_72__26_,s_r_72__25_,s_r_72__24_,s_r_72__23_,s_r_72__22_,
  s_r_72__21_,s_r_72__20_,s_r_72__19_,s_r_72__18_,s_r_72__17_,s_r_72__16_,s_r_72__15_,
  s_r_72__14_,s_r_72__13_,s_r_72__12_,s_r_72__11_,s_r_72__10_,s_r_72__9_,
  s_r_72__8_,s_r_72__7_,s_r_72__6_,s_r_72__5_,s_r_72__4_,s_r_72__3_,s_r_72__2_,s_r_72__1_,
  s_r_72__0_,s_r_71__127_,s_r_71__126_,s_r_71__125_,s_r_71__124_,s_r_71__123_,
  s_r_71__122_,s_r_71__121_,s_r_71__120_,s_r_71__119_,s_r_71__118_,s_r_71__117_,
  s_r_71__116_,s_r_71__115_,s_r_71__114_,s_r_71__113_,s_r_71__112_,s_r_71__111_,
  s_r_71__110_,s_r_71__109_,s_r_71__108_,s_r_71__107_,s_r_71__106_,s_r_71__105_,
  s_r_71__104_,s_r_71__103_,s_r_71__102_,s_r_71__101_,s_r_71__100_,s_r_71__99_,s_r_71__98_,
  s_r_71__97_,s_r_71__96_,s_r_71__95_,s_r_71__94_,s_r_71__93_,s_r_71__92_,
  s_r_71__91_,s_r_71__90_,s_r_71__89_,s_r_71__88_,s_r_71__87_,s_r_71__86_,s_r_71__85_,
  s_r_71__84_,s_r_71__83_,s_r_71__82_,s_r_71__81_,s_r_71__80_,s_r_71__79_,s_r_71__78_,
  s_r_71__77_,s_r_71__76_,s_r_71__75_,s_r_71__74_,s_r_71__73_,s_r_71__72_,
  s_r_71__71_,s_r_71__70_,s_r_71__69_,s_r_71__68_,s_r_71__67_,s_r_71__66_,s_r_71__65_,
  s_r_71__64_,s_r_71__63_,s_r_71__62_,s_r_71__61_,s_r_71__60_,s_r_71__59_,s_r_71__58_,
  s_r_71__57_,s_r_71__56_,s_r_71__55_,s_r_71__54_,s_r_71__53_,s_r_71__52_,
  s_r_71__51_,s_r_71__50_,s_r_71__49_,s_r_71__48_,s_r_71__47_,s_r_71__46_,s_r_71__45_,
  s_r_71__44_,s_r_71__43_,s_r_71__42_,s_r_71__41_,s_r_71__40_,s_r_71__39_,s_r_71__38_,
  s_r_71__37_,s_r_71__36_,s_r_71__35_,s_r_71__34_,s_r_71__33_,s_r_71__32_,
  s_r_71__31_,s_r_71__30_,s_r_71__29_,s_r_71__28_,s_r_71__27_,s_r_71__26_,s_r_71__25_,
  s_r_71__24_,s_r_71__23_,s_r_71__22_,s_r_71__21_,s_r_71__20_,s_r_71__19_,s_r_71__18_,
  s_r_71__17_,s_r_71__16_,s_r_71__15_,s_r_71__14_,s_r_71__13_,s_r_71__12_,
  s_r_71__11_,s_r_71__10_,s_r_71__9_,s_r_71__8_,s_r_71__7_,s_r_71__6_,s_r_71__5_,s_r_71__4_,
  s_r_71__3_,s_r_71__2_,s_r_71__1_,s_r_71__0_,prod_accum_74__75_,
  prod_accum_74__74_,prod_accum_74__73_,prod_accum_74__72_,prod_accum_74__71_,prod_accum_74__70_,
  prod_accum_74__69_,prod_accum_74__68_,prod_accum_74__67_,prod_accum_74__66_,
  prod_accum_74__65_,prod_accum_74__64_,prod_accum_74__63_,prod_accum_74__62_,
  prod_accum_74__61_,prod_accum_74__60_,prod_accum_74__59_,prod_accum_74__58_,
  prod_accum_74__57_,prod_accum_74__56_,prod_accum_74__55_,prod_accum_74__54_,
  prod_accum_74__53_,prod_accum_74__52_,prod_accum_74__51_,prod_accum_74__50_,prod_accum_74__49_,
  prod_accum_74__48_,prod_accum_74__47_,prod_accum_74__46_,prod_accum_74__45_,
  prod_accum_74__44_,prod_accum_74__43_,prod_accum_74__42_,prod_accum_74__41_,
  prod_accum_74__40_,prod_accum_74__39_,prod_accum_74__38_,prod_accum_74__37_,
  prod_accum_74__36_,prod_accum_74__35_,prod_accum_74__34_,prod_accum_74__33_,prod_accum_74__32_,
  prod_accum_74__31_,prod_accum_74__30_,prod_accum_74__29_,prod_accum_74__28_,
  prod_accum_74__27_,prod_accum_74__26_,prod_accum_74__25_,prod_accum_74__24_,
  prod_accum_74__23_,prod_accum_74__22_,prod_accum_74__21_,prod_accum_74__20_,
  prod_accum_74__19_,prod_accum_74__18_,prod_accum_74__17_,prod_accum_74__16_,
  prod_accum_74__15_,prod_accum_74__14_,prod_accum_74__13_,prod_accum_74__12_,prod_accum_74__11_,
  prod_accum_74__10_,prod_accum_74__9_,prod_accum_74__8_,prod_accum_74__7_,
  prod_accum_74__6_,prod_accum_74__5_,prod_accum_74__4_,prod_accum_74__3_,
  prod_accum_74__2_,prod_accum_74__1_,prod_accum_74__0_,prod_accum_73__74_,prod_accum_73__73_,
  prod_accum_73__72_,prod_accum_73__71_,prod_accum_73__70_,prod_accum_73__69_,
  prod_accum_73__68_,prod_accum_73__67_,prod_accum_73__66_,prod_accum_73__65_,
  prod_accum_73__64_,prod_accum_73__63_,prod_accum_73__62_,prod_accum_73__61_,
  prod_accum_73__60_,prod_accum_73__59_,prod_accum_73__58_,prod_accum_73__57_,prod_accum_73__56_,
  prod_accum_73__55_,prod_accum_73__54_,prod_accum_73__53_,prod_accum_73__52_,
  prod_accum_73__51_,prod_accum_73__50_,prod_accum_73__49_,prod_accum_73__48_,
  prod_accum_73__47_,prod_accum_73__46_,prod_accum_73__45_,prod_accum_73__44_,
  prod_accum_73__43_,prod_accum_73__42_,prod_accum_73__41_,prod_accum_73__40_,
  prod_accum_73__39_,prod_accum_73__38_,prod_accum_73__37_,prod_accum_73__36_,prod_accum_73__35_,
  prod_accum_73__34_,prod_accum_73__33_,prod_accum_73__32_,prod_accum_73__31_,
  prod_accum_73__30_,prod_accum_73__29_,prod_accum_73__28_,prod_accum_73__27_,
  prod_accum_73__26_,prod_accum_73__25_,prod_accum_73__24_,prod_accum_73__23_,
  prod_accum_73__22_,prod_accum_73__21_,prod_accum_73__20_,prod_accum_73__19_,
  prod_accum_73__18_,prod_accum_73__17_,prod_accum_73__16_,prod_accum_73__15_,prod_accum_73__14_,
  prod_accum_73__13_,prod_accum_73__12_,prod_accum_73__11_,prod_accum_73__10_,
  prod_accum_73__9_,prod_accum_73__8_,prod_accum_73__7_,prod_accum_73__6_,
  prod_accum_73__5_,prod_accum_73__4_,prod_accum_73__3_,prod_accum_73__2_,prod_accum_73__1_,
  prod_accum_73__0_,prod_accum_72__73_,prod_accum_72__72_,prod_accum_72__71_,
  prod_accum_72__70_,prod_accum_72__69_,prod_accum_72__68_,prod_accum_72__67_,
  prod_accum_72__66_,prod_accum_72__65_,prod_accum_72__64_,prod_accum_72__63_,
  prod_accum_72__62_,prod_accum_72__61_,prod_accum_72__60_,prod_accum_72__59_,prod_accum_72__58_,
  prod_accum_72__57_,prod_accum_72__56_,prod_accum_72__55_,prod_accum_72__54_,
  prod_accum_72__53_,prod_accum_72__52_,prod_accum_72__51_,prod_accum_72__50_,
  prod_accum_72__49_,prod_accum_72__48_,prod_accum_72__47_,prod_accum_72__46_,
  prod_accum_72__45_,prod_accum_72__44_,prod_accum_72__43_,prod_accum_72__42_,prod_accum_72__41_,
  prod_accum_72__40_,prod_accum_72__39_,prod_accum_72__38_,prod_accum_72__37_,
  prod_accum_72__36_,prod_accum_72__35_,prod_accum_72__34_,prod_accum_72__33_,
  prod_accum_72__32_,prod_accum_72__31_,prod_accum_72__30_,prod_accum_72__29_,
  prod_accum_72__28_,prod_accum_72__27_,prod_accum_72__26_,prod_accum_72__25_,
  prod_accum_72__24_,prod_accum_72__23_,prod_accum_72__22_,prod_accum_72__21_,prod_accum_72__20_,
  prod_accum_72__19_,prod_accum_72__18_,prod_accum_72__17_,prod_accum_72__16_,
  prod_accum_72__15_,prod_accum_72__14_,prod_accum_72__13_,prod_accum_72__12_,
  prod_accum_72__11_,prod_accum_72__10_,prod_accum_72__9_,prod_accum_72__8_,
  prod_accum_72__7_,prod_accum_72__6_,prod_accum_72__5_,prod_accum_72__4_,prod_accum_72__3_,
  prod_accum_72__2_,prod_accum_72__1_,prod_accum_72__0_,prod_accum_71__72_,
  prod_accum_71__71_,prod_accum_71__70_,prod_accum_71__69_,prod_accum_71__68_,
  prod_accum_71__67_,prod_accum_71__66_,prod_accum_71__65_,prod_accum_71__64_,prod_accum_71__63_,
  prod_accum_71__62_,prod_accum_71__61_,prod_accum_71__60_,prod_accum_71__59_,
  prod_accum_71__58_,prod_accum_71__57_,prod_accum_71__56_,prod_accum_71__55_,
  prod_accum_71__54_,prod_accum_71__53_,prod_accum_71__52_,prod_accum_71__51_,
  prod_accum_71__50_,prod_accum_71__49_,prod_accum_71__48_,prod_accum_71__47_,
  prod_accum_71__46_,prod_accum_71__45_,prod_accum_71__44_,prod_accum_71__43_,prod_accum_71__42_,
  prod_accum_71__41_,prod_accum_71__40_,prod_accum_71__39_,prod_accum_71__38_,
  prod_accum_71__37_,prod_accum_71__36_,prod_accum_71__35_,prod_accum_71__34_,
  prod_accum_71__33_,prod_accum_71__32_,prod_accum_71__31_,prod_accum_71__30_,
  prod_accum_71__29_,prod_accum_71__28_,prod_accum_71__27_,prod_accum_71__26_,
  prod_accum_71__25_,prod_accum_71__24_,prod_accum_71__23_,prod_accum_71__22_,prod_accum_71__21_,
  prod_accum_71__20_,prod_accum_71__19_,prod_accum_71__18_,prod_accum_71__17_,
  prod_accum_71__16_,prod_accum_71__15_,prod_accum_71__14_,prod_accum_71__13_,
  prod_accum_71__12_,prod_accum_71__11_,prod_accum_71__10_,prod_accum_71__9_,
  prod_accum_71__8_,prod_accum_71__7_,prod_accum_71__6_,prod_accum_71__5_,prod_accum_71__4_,
  prod_accum_71__3_,prod_accum_71__2_,prod_accum_71__1_,prod_accum_71__0_,s_r_78__127_,
  s_r_78__126_,s_r_78__125_,s_r_78__124_,s_r_78__123_,s_r_78__122_,s_r_78__121_,
  s_r_78__120_,s_r_78__119_,s_r_78__118_,s_r_78__117_,s_r_78__116_,s_r_78__115_,
  s_r_78__114_,s_r_78__113_,s_r_78__112_,s_r_78__111_,s_r_78__110_,s_r_78__109_,
  s_r_78__108_,s_r_78__107_,s_r_78__106_,s_r_78__105_,s_r_78__104_,s_r_78__103_,
  s_r_78__102_,s_r_78__101_,s_r_78__100_,s_r_78__99_,s_r_78__98_,s_r_78__97_,s_r_78__96_,
  s_r_78__95_,s_r_78__94_,s_r_78__93_,s_r_78__92_,s_r_78__91_,s_r_78__90_,
  s_r_78__89_,s_r_78__88_,s_r_78__87_,s_r_78__86_,s_r_78__85_,s_r_78__84_,s_r_78__83_,
  s_r_78__82_,s_r_78__81_,s_r_78__80_,s_r_78__79_,s_r_78__78_,s_r_78__77_,s_r_78__76_,
  s_r_78__75_,s_r_78__74_,s_r_78__73_,s_r_78__72_,s_r_78__71_,s_r_78__70_,
  s_r_78__69_,s_r_78__68_,s_r_78__67_,s_r_78__66_,s_r_78__65_,s_r_78__64_,s_r_78__63_,
  s_r_78__62_,s_r_78__61_,s_r_78__60_,s_r_78__59_,s_r_78__58_,s_r_78__57_,s_r_78__56_,
  s_r_78__55_,s_r_78__54_,s_r_78__53_,s_r_78__52_,s_r_78__51_,s_r_78__50_,
  s_r_78__49_,s_r_78__48_,s_r_78__47_,s_r_78__46_,s_r_78__45_,s_r_78__44_,s_r_78__43_,
  s_r_78__42_,s_r_78__41_,s_r_78__40_,s_r_78__39_,s_r_78__38_,s_r_78__37_,s_r_78__36_,
  s_r_78__35_,s_r_78__34_,s_r_78__33_,s_r_78__32_,s_r_78__31_,s_r_78__30_,
  s_r_78__29_,s_r_78__28_,s_r_78__27_,s_r_78__26_,s_r_78__25_,s_r_78__24_,s_r_78__23_,
  s_r_78__22_,s_r_78__21_,s_r_78__20_,s_r_78__19_,s_r_78__18_,s_r_78__17_,s_r_78__16_,
  s_r_78__15_,s_r_78__14_,s_r_78__13_,s_r_78__12_,s_r_78__11_,s_r_78__10_,
  s_r_78__9_,s_r_78__8_,s_r_78__7_,s_r_78__6_,s_r_78__5_,s_r_78__4_,s_r_78__3_,s_r_78__2_,
  s_r_78__1_,s_r_78__0_,s_r_77__127_,s_r_77__126_,s_r_77__125_,s_r_77__124_,
  s_r_77__123_,s_r_77__122_,s_r_77__121_,s_r_77__120_,s_r_77__119_,s_r_77__118_,
  s_r_77__117_,s_r_77__116_,s_r_77__115_,s_r_77__114_,s_r_77__113_,s_r_77__112_,
  s_r_77__111_,s_r_77__110_,s_r_77__109_,s_r_77__108_,s_r_77__107_,s_r_77__106_,s_r_77__105_,
  s_r_77__104_,s_r_77__103_,s_r_77__102_,s_r_77__101_,s_r_77__100_,s_r_77__99_,
  s_r_77__98_,s_r_77__97_,s_r_77__96_,s_r_77__95_,s_r_77__94_,s_r_77__93_,s_r_77__92_,
  s_r_77__91_,s_r_77__90_,s_r_77__89_,s_r_77__88_,s_r_77__87_,s_r_77__86_,
  s_r_77__85_,s_r_77__84_,s_r_77__83_,s_r_77__82_,s_r_77__81_,s_r_77__80_,s_r_77__79_,
  s_r_77__78_,s_r_77__77_,s_r_77__76_,s_r_77__75_,s_r_77__74_,s_r_77__73_,s_r_77__72_,
  s_r_77__71_,s_r_77__70_,s_r_77__69_,s_r_77__68_,s_r_77__67_,s_r_77__66_,
  s_r_77__65_,s_r_77__64_,s_r_77__63_,s_r_77__62_,s_r_77__61_,s_r_77__60_,s_r_77__59_,
  s_r_77__58_,s_r_77__57_,s_r_77__56_,s_r_77__55_,s_r_77__54_,s_r_77__53_,s_r_77__52_,
  s_r_77__51_,s_r_77__50_,s_r_77__49_,s_r_77__48_,s_r_77__47_,s_r_77__46_,
  s_r_77__45_,s_r_77__44_,s_r_77__43_,s_r_77__42_,s_r_77__41_,s_r_77__40_,s_r_77__39_,
  s_r_77__38_,s_r_77__37_,s_r_77__36_,s_r_77__35_,s_r_77__34_,s_r_77__33_,s_r_77__32_,
  s_r_77__31_,s_r_77__30_,s_r_77__29_,s_r_77__28_,s_r_77__27_,s_r_77__26_,
  s_r_77__25_,s_r_77__24_,s_r_77__23_,s_r_77__22_,s_r_77__21_,s_r_77__20_,s_r_77__19_,
  s_r_77__18_,s_r_77__17_,s_r_77__16_,s_r_77__15_,s_r_77__14_,s_r_77__13_,s_r_77__12_,
  s_r_77__11_,s_r_77__10_,s_r_77__9_,s_r_77__8_,s_r_77__7_,s_r_77__6_,s_r_77__5_,
  s_r_77__4_,s_r_77__3_,s_r_77__2_,s_r_77__1_,s_r_77__0_,s_r_76__127_,s_r_76__126_,
  s_r_76__125_,s_r_76__124_,s_r_76__123_,s_r_76__122_,s_r_76__121_,s_r_76__120_,
  s_r_76__119_,s_r_76__118_,s_r_76__117_,s_r_76__116_,s_r_76__115_,s_r_76__114_,
  s_r_76__113_,s_r_76__112_,s_r_76__111_,s_r_76__110_,s_r_76__109_,s_r_76__108_,
  s_r_76__107_,s_r_76__106_,s_r_76__105_,s_r_76__104_,s_r_76__103_,s_r_76__102_,
  s_r_76__101_,s_r_76__100_,s_r_76__99_,s_r_76__98_,s_r_76__97_,s_r_76__96_,s_r_76__95_,
  s_r_76__94_,s_r_76__93_,s_r_76__92_,s_r_76__91_,s_r_76__90_,s_r_76__89_,
  s_r_76__88_,s_r_76__87_,s_r_76__86_,s_r_76__85_,s_r_76__84_,s_r_76__83_,s_r_76__82_,
  s_r_76__81_,s_r_76__80_,s_r_76__79_,s_r_76__78_,s_r_76__77_,s_r_76__76_,s_r_76__75_,
  s_r_76__74_,s_r_76__73_,s_r_76__72_,s_r_76__71_,s_r_76__70_,s_r_76__69_,
  s_r_76__68_,s_r_76__67_,s_r_76__66_,s_r_76__65_,s_r_76__64_,s_r_76__63_,s_r_76__62_,
  s_r_76__61_,s_r_76__60_,s_r_76__59_,s_r_76__58_,s_r_76__57_,s_r_76__56_,s_r_76__55_,
  s_r_76__54_,s_r_76__53_,s_r_76__52_,s_r_76__51_,s_r_76__50_,s_r_76__49_,
  s_r_76__48_,s_r_76__47_,s_r_76__46_,s_r_76__45_,s_r_76__44_,s_r_76__43_,s_r_76__42_,
  s_r_76__41_,s_r_76__40_,s_r_76__39_,s_r_76__38_,s_r_76__37_,s_r_76__36_,s_r_76__35_,
  s_r_76__34_,s_r_76__33_,s_r_76__32_,s_r_76__31_,s_r_76__30_,s_r_76__29_,
  s_r_76__28_,s_r_76__27_,s_r_76__26_,s_r_76__25_,s_r_76__24_,s_r_76__23_,s_r_76__22_,
  s_r_76__21_,s_r_76__20_,s_r_76__19_,s_r_76__18_,s_r_76__17_,s_r_76__16_,s_r_76__15_,
  s_r_76__14_,s_r_76__13_,s_r_76__12_,s_r_76__11_,s_r_76__10_,s_r_76__9_,s_r_76__8_,
  s_r_76__7_,s_r_76__6_,s_r_76__5_,s_r_76__4_,s_r_76__3_,s_r_76__2_,s_r_76__1_,
  s_r_76__0_,s_r_75__127_,s_r_75__126_,s_r_75__125_,s_r_75__124_,s_r_75__123_,
  s_r_75__122_,s_r_75__121_,s_r_75__120_,s_r_75__119_,s_r_75__118_,s_r_75__117_,
  s_r_75__116_,s_r_75__115_,s_r_75__114_,s_r_75__113_,s_r_75__112_,s_r_75__111_,
  s_r_75__110_,s_r_75__109_,s_r_75__108_,s_r_75__107_,s_r_75__106_,s_r_75__105_,s_r_75__104_,
  s_r_75__103_,s_r_75__102_,s_r_75__101_,s_r_75__100_,s_r_75__99_,s_r_75__98_,
  s_r_75__97_,s_r_75__96_,s_r_75__95_,s_r_75__94_,s_r_75__93_,s_r_75__92_,s_r_75__91_,
  s_r_75__90_,s_r_75__89_,s_r_75__88_,s_r_75__87_,s_r_75__86_,s_r_75__85_,
  s_r_75__84_,s_r_75__83_,s_r_75__82_,s_r_75__81_,s_r_75__80_,s_r_75__79_,s_r_75__78_,
  s_r_75__77_,s_r_75__76_,s_r_75__75_,s_r_75__74_,s_r_75__73_,s_r_75__72_,s_r_75__71_,
  s_r_75__70_,s_r_75__69_,s_r_75__68_,s_r_75__67_,s_r_75__66_,s_r_75__65_,
  s_r_75__64_,s_r_75__63_,s_r_75__62_,s_r_75__61_,s_r_75__60_,s_r_75__59_,s_r_75__58_,
  s_r_75__57_,s_r_75__56_,s_r_75__55_,s_r_75__54_,s_r_75__53_,s_r_75__52_,s_r_75__51_,
  s_r_75__50_,s_r_75__49_,s_r_75__48_,s_r_75__47_,s_r_75__46_,s_r_75__45_,
  s_r_75__44_,s_r_75__43_,s_r_75__42_,s_r_75__41_,s_r_75__40_,s_r_75__39_,s_r_75__38_,
  s_r_75__37_,s_r_75__36_,s_r_75__35_,s_r_75__34_,s_r_75__33_,s_r_75__32_,s_r_75__31_,
  s_r_75__30_,s_r_75__29_,s_r_75__28_,s_r_75__27_,s_r_75__26_,s_r_75__25_,
  s_r_75__24_,s_r_75__23_,s_r_75__22_,s_r_75__21_,s_r_75__20_,s_r_75__19_,s_r_75__18_,
  s_r_75__17_,s_r_75__16_,s_r_75__15_,s_r_75__14_,s_r_75__13_,s_r_75__12_,s_r_75__11_,
  s_r_75__10_,s_r_75__9_,s_r_75__8_,s_r_75__7_,s_r_75__6_,s_r_75__5_,s_r_75__4_,
  s_r_75__3_,s_r_75__2_,s_r_75__1_,s_r_75__0_,prod_accum_78__79_,prod_accum_78__78_,
  prod_accum_78__77_,prod_accum_78__76_,prod_accum_78__75_,prod_accum_78__74_,
  prod_accum_78__73_,prod_accum_78__72_,prod_accum_78__71_,prod_accum_78__70_,
  prod_accum_78__69_,prod_accum_78__68_,prod_accum_78__67_,prod_accum_78__66_,
  prod_accum_78__65_,prod_accum_78__64_,prod_accum_78__63_,prod_accum_78__62_,
  prod_accum_78__61_,prod_accum_78__60_,prod_accum_78__59_,prod_accum_78__58_,prod_accum_78__57_,
  prod_accum_78__56_,prod_accum_78__55_,prod_accum_78__54_,prod_accum_78__53_,
  prod_accum_78__52_,prod_accum_78__51_,prod_accum_78__50_,prod_accum_78__49_,
  prod_accum_78__48_,prod_accum_78__47_,prod_accum_78__46_,prod_accum_78__45_,
  prod_accum_78__44_,prod_accum_78__43_,prod_accum_78__42_,prod_accum_78__41_,
  prod_accum_78__40_,prod_accum_78__39_,prod_accum_78__38_,prod_accum_78__37_,prod_accum_78__36_,
  prod_accum_78__35_,prod_accum_78__34_,prod_accum_78__33_,prod_accum_78__32_,
  prod_accum_78__31_,prod_accum_78__30_,prod_accum_78__29_,prod_accum_78__28_,
  prod_accum_78__27_,prod_accum_78__26_,prod_accum_78__25_,prod_accum_78__24_,
  prod_accum_78__23_,prod_accum_78__22_,prod_accum_78__21_,prod_accum_78__20_,
  prod_accum_78__19_,prod_accum_78__18_,prod_accum_78__17_,prod_accum_78__16_,prod_accum_78__15_,
  prod_accum_78__14_,prod_accum_78__13_,prod_accum_78__12_,prod_accum_78__11_,
  prod_accum_78__10_,prod_accum_78__9_,prod_accum_78__8_,prod_accum_78__7_,
  prod_accum_78__6_,prod_accum_78__5_,prod_accum_78__4_,prod_accum_78__3_,prod_accum_78__2_,
  prod_accum_78__1_,prod_accum_78__0_,prod_accum_77__78_,prod_accum_77__77_,
  prod_accum_77__76_,prod_accum_77__75_,prod_accum_77__74_,prod_accum_77__73_,
  prod_accum_77__72_,prod_accum_77__71_,prod_accum_77__70_,prod_accum_77__69_,
  prod_accum_77__68_,prod_accum_77__67_,prod_accum_77__66_,prod_accum_77__65_,prod_accum_77__64_,
  prod_accum_77__63_,prod_accum_77__62_,prod_accum_77__61_,prod_accum_77__60_,
  prod_accum_77__59_,prod_accum_77__58_,prod_accum_77__57_,prod_accum_77__56_,
  prod_accum_77__55_,prod_accum_77__54_,prod_accum_77__53_,prod_accum_77__52_,
  prod_accum_77__51_,prod_accum_77__50_,prod_accum_77__49_,prod_accum_77__48_,prod_accum_77__47_,
  prod_accum_77__46_,prod_accum_77__45_,prod_accum_77__44_,prod_accum_77__43_,
  prod_accum_77__42_,prod_accum_77__41_,prod_accum_77__40_,prod_accum_77__39_,
  prod_accum_77__38_,prod_accum_77__37_,prod_accum_77__36_,prod_accum_77__35_,
  prod_accum_77__34_,prod_accum_77__33_,prod_accum_77__32_,prod_accum_77__31_,
  prod_accum_77__30_,prod_accum_77__29_,prod_accum_77__28_,prod_accum_77__27_,prod_accum_77__26_,
  prod_accum_77__25_,prod_accum_77__24_,prod_accum_77__23_,prod_accum_77__22_,
  prod_accum_77__21_,prod_accum_77__20_,prod_accum_77__19_,prod_accum_77__18_,
  prod_accum_77__17_,prod_accum_77__16_,prod_accum_77__15_,prod_accum_77__14_,
  prod_accum_77__13_,prod_accum_77__12_,prod_accum_77__11_,prod_accum_77__10_,
  prod_accum_77__9_,prod_accum_77__8_,prod_accum_77__7_,prod_accum_77__6_,prod_accum_77__5_,
  prod_accum_77__4_,prod_accum_77__3_,prod_accum_77__2_,prod_accum_77__1_,
  prod_accum_77__0_,prod_accum_76__77_,prod_accum_76__76_,prod_accum_76__75_,prod_accum_76__74_,
  prod_accum_76__73_,prod_accum_76__72_,prod_accum_76__71_,prod_accum_76__70_,
  prod_accum_76__69_,prod_accum_76__68_,prod_accum_76__67_,prod_accum_76__66_,
  prod_accum_76__65_,prod_accum_76__64_,prod_accum_76__63_,prod_accum_76__62_,
  prod_accum_76__61_,prod_accum_76__60_,prod_accum_76__59_,prod_accum_76__58_,
  prod_accum_76__57_,prod_accum_76__56_,prod_accum_76__55_,prod_accum_76__54_,prod_accum_76__53_,
  prod_accum_76__52_,prod_accum_76__51_,prod_accum_76__50_,prod_accum_76__49_,
  prod_accum_76__48_,prod_accum_76__47_,prod_accum_76__46_,prod_accum_76__45_,
  prod_accum_76__44_,prod_accum_76__43_,prod_accum_76__42_,prod_accum_76__41_,
  prod_accum_76__40_,prod_accum_76__39_,prod_accum_76__38_,prod_accum_76__37_,
  prod_accum_76__36_,prod_accum_76__35_,prod_accum_76__34_,prod_accum_76__33_,prod_accum_76__32_,
  prod_accum_76__31_,prod_accum_76__30_,prod_accum_76__29_,prod_accum_76__28_,
  prod_accum_76__27_,prod_accum_76__26_,prod_accum_76__25_,prod_accum_76__24_,
  prod_accum_76__23_,prod_accum_76__22_,prod_accum_76__21_,prod_accum_76__20_,
  prod_accum_76__19_,prod_accum_76__18_,prod_accum_76__17_,prod_accum_76__16_,prod_accum_76__15_,
  prod_accum_76__14_,prod_accum_76__13_,prod_accum_76__12_,prod_accum_76__11_,
  prod_accum_76__10_,prod_accum_76__9_,prod_accum_76__8_,prod_accum_76__7_,
  prod_accum_76__6_,prod_accum_76__5_,prod_accum_76__4_,prod_accum_76__3_,prod_accum_76__2_,
  prod_accum_76__1_,prod_accum_76__0_,prod_accum_75__76_,prod_accum_75__75_,
  prod_accum_75__74_,prod_accum_75__73_,prod_accum_75__72_,prod_accum_75__71_,
  prod_accum_75__70_,prod_accum_75__69_,prod_accum_75__68_,prod_accum_75__67_,
  prod_accum_75__66_,prod_accum_75__65_,prod_accum_75__64_,prod_accum_75__63_,prod_accum_75__62_,
  prod_accum_75__61_,prod_accum_75__60_,prod_accum_75__59_,prod_accum_75__58_,
  prod_accum_75__57_,prod_accum_75__56_,prod_accum_75__55_,prod_accum_75__54_,
  prod_accum_75__53_,prod_accum_75__52_,prod_accum_75__51_,prod_accum_75__50_,
  prod_accum_75__49_,prod_accum_75__48_,prod_accum_75__47_,prod_accum_75__46_,
  prod_accum_75__45_,prod_accum_75__44_,prod_accum_75__43_,prod_accum_75__42_,prod_accum_75__41_,
  prod_accum_75__40_,prod_accum_75__39_,prod_accum_75__38_,prod_accum_75__37_,
  prod_accum_75__36_,prod_accum_75__35_,prod_accum_75__34_,prod_accum_75__33_,
  prod_accum_75__32_,prod_accum_75__31_,prod_accum_75__30_,prod_accum_75__29_,
  prod_accum_75__28_,prod_accum_75__27_,prod_accum_75__26_,prod_accum_75__25_,
  prod_accum_75__24_,prod_accum_75__23_,prod_accum_75__22_,prod_accum_75__21_,prod_accum_75__20_,
  prod_accum_75__19_,prod_accum_75__18_,prod_accum_75__17_,prod_accum_75__16_,
  prod_accum_75__15_,prod_accum_75__14_,prod_accum_75__13_,prod_accum_75__12_,
  prod_accum_75__11_,prod_accum_75__10_,prod_accum_75__9_,prod_accum_75__8_,
  prod_accum_75__7_,prod_accum_75__6_,prod_accum_75__5_,prod_accum_75__4_,prod_accum_75__3_,
  prod_accum_75__2_,prod_accum_75__1_,prod_accum_75__0_,s_r_82__127_,s_r_82__126_,
  s_r_82__125_,s_r_82__124_,s_r_82__123_,s_r_82__122_,s_r_82__121_,s_r_82__120_,
  s_r_82__119_,s_r_82__118_,s_r_82__117_,s_r_82__116_,s_r_82__115_,s_r_82__114_,
  s_r_82__113_,s_r_82__112_,s_r_82__111_,s_r_82__110_,s_r_82__109_,s_r_82__108_,
  s_r_82__107_,s_r_82__106_,s_r_82__105_,s_r_82__104_,s_r_82__103_,s_r_82__102_,s_r_82__101_,
  s_r_82__100_,s_r_82__99_,s_r_82__98_,s_r_82__97_,s_r_82__96_,s_r_82__95_,
  s_r_82__94_,s_r_82__93_,s_r_82__92_,s_r_82__91_,s_r_82__90_,s_r_82__89_,s_r_82__88_,
  s_r_82__87_,s_r_82__86_,s_r_82__85_,s_r_82__84_,s_r_82__83_,s_r_82__82_,s_r_82__81_,
  s_r_82__80_,s_r_82__79_,s_r_82__78_,s_r_82__77_,s_r_82__76_,s_r_82__75_,
  s_r_82__74_,s_r_82__73_,s_r_82__72_,s_r_82__71_,s_r_82__70_,s_r_82__69_,s_r_82__68_,
  s_r_82__67_,s_r_82__66_,s_r_82__65_,s_r_82__64_,s_r_82__63_,s_r_82__62_,s_r_82__61_,
  s_r_82__60_,s_r_82__59_,s_r_82__58_,s_r_82__57_,s_r_82__56_,s_r_82__55_,
  s_r_82__54_,s_r_82__53_,s_r_82__52_,s_r_82__51_,s_r_82__50_,s_r_82__49_,s_r_82__48_,
  s_r_82__47_,s_r_82__46_,s_r_82__45_,s_r_82__44_,s_r_82__43_,s_r_82__42_,s_r_82__41_,
  s_r_82__40_,s_r_82__39_,s_r_82__38_,s_r_82__37_,s_r_82__36_,s_r_82__35_,
  s_r_82__34_,s_r_82__33_,s_r_82__32_,s_r_82__31_,s_r_82__30_,s_r_82__29_,s_r_82__28_,
  s_r_82__27_,s_r_82__26_,s_r_82__25_,s_r_82__24_,s_r_82__23_,s_r_82__22_,s_r_82__21_,
  s_r_82__20_,s_r_82__19_,s_r_82__18_,s_r_82__17_,s_r_82__16_,s_r_82__15_,
  s_r_82__14_,s_r_82__13_,s_r_82__12_,s_r_82__11_,s_r_82__10_,s_r_82__9_,s_r_82__8_,
  s_r_82__7_,s_r_82__6_,s_r_82__5_,s_r_82__4_,s_r_82__3_,s_r_82__2_,s_r_82__1_,
  s_r_82__0_,s_r_81__127_,s_r_81__126_,s_r_81__125_,s_r_81__124_,s_r_81__123_,s_r_81__122_,
  s_r_81__121_,s_r_81__120_,s_r_81__119_,s_r_81__118_,s_r_81__117_,s_r_81__116_,
  s_r_81__115_,s_r_81__114_,s_r_81__113_,s_r_81__112_,s_r_81__111_,s_r_81__110_,
  s_r_81__109_,s_r_81__108_,s_r_81__107_,s_r_81__106_,s_r_81__105_,s_r_81__104_,
  s_r_81__103_,s_r_81__102_,s_r_81__101_,s_r_81__100_,s_r_81__99_,s_r_81__98_,
  s_r_81__97_,s_r_81__96_,s_r_81__95_,s_r_81__94_,s_r_81__93_,s_r_81__92_,s_r_81__91_,
  s_r_81__90_,s_r_81__89_,s_r_81__88_,s_r_81__87_,s_r_81__86_,s_r_81__85_,s_r_81__84_,
  s_r_81__83_,s_r_81__82_,s_r_81__81_,s_r_81__80_,s_r_81__79_,s_r_81__78_,
  s_r_81__77_,s_r_81__76_,s_r_81__75_,s_r_81__74_,s_r_81__73_,s_r_81__72_,s_r_81__71_,
  s_r_81__70_,s_r_81__69_,s_r_81__68_,s_r_81__67_,s_r_81__66_,s_r_81__65_,s_r_81__64_,
  s_r_81__63_,s_r_81__62_,s_r_81__61_,s_r_81__60_,s_r_81__59_,s_r_81__58_,
  s_r_81__57_,s_r_81__56_,s_r_81__55_,s_r_81__54_,s_r_81__53_,s_r_81__52_,s_r_81__51_,
  s_r_81__50_,s_r_81__49_,s_r_81__48_,s_r_81__47_,s_r_81__46_,s_r_81__45_,s_r_81__44_,
  s_r_81__43_,s_r_81__42_,s_r_81__41_,s_r_81__40_,s_r_81__39_,s_r_81__38_,
  s_r_81__37_,s_r_81__36_,s_r_81__35_,s_r_81__34_,s_r_81__33_,s_r_81__32_,s_r_81__31_,
  s_r_81__30_,s_r_81__29_,s_r_81__28_,s_r_81__27_,s_r_81__26_,s_r_81__25_,s_r_81__24_,
  s_r_81__23_,s_r_81__22_,s_r_81__21_,s_r_81__20_,s_r_81__19_,s_r_81__18_,
  s_r_81__17_,s_r_81__16_,s_r_81__15_,s_r_81__14_,s_r_81__13_,s_r_81__12_,s_r_81__11_,
  s_r_81__10_,s_r_81__9_,s_r_81__8_,s_r_81__7_,s_r_81__6_,s_r_81__5_,s_r_81__4_,
  s_r_81__3_,s_r_81__2_,s_r_81__1_,s_r_81__0_,s_r_80__127_,s_r_80__126_,s_r_80__125_,
  s_r_80__124_,s_r_80__123_,s_r_80__122_,s_r_80__121_,s_r_80__120_,s_r_80__119_,
  s_r_80__118_,s_r_80__117_,s_r_80__116_,s_r_80__115_,s_r_80__114_,s_r_80__113_,
  s_r_80__112_,s_r_80__111_,s_r_80__110_,s_r_80__109_,s_r_80__108_,s_r_80__107_,
  s_r_80__106_,s_r_80__105_,s_r_80__104_,s_r_80__103_,s_r_80__102_,s_r_80__101_,s_r_80__100_,
  s_r_80__99_,s_r_80__98_,s_r_80__97_,s_r_80__96_,s_r_80__95_,s_r_80__94_,
  s_r_80__93_,s_r_80__92_,s_r_80__91_,s_r_80__90_,s_r_80__89_,s_r_80__88_,s_r_80__87_,
  s_r_80__86_,s_r_80__85_,s_r_80__84_,s_r_80__83_,s_r_80__82_,s_r_80__81_,s_r_80__80_,
  s_r_80__79_,s_r_80__78_,s_r_80__77_,s_r_80__76_,s_r_80__75_,s_r_80__74_,
  s_r_80__73_,s_r_80__72_,s_r_80__71_,s_r_80__70_,s_r_80__69_,s_r_80__68_,s_r_80__67_,
  s_r_80__66_,s_r_80__65_,s_r_80__64_,s_r_80__63_,s_r_80__62_,s_r_80__61_,s_r_80__60_,
  s_r_80__59_,s_r_80__58_,s_r_80__57_,s_r_80__56_,s_r_80__55_,s_r_80__54_,
  s_r_80__53_,s_r_80__52_,s_r_80__51_,s_r_80__50_,s_r_80__49_,s_r_80__48_,s_r_80__47_,
  s_r_80__46_,s_r_80__45_,s_r_80__44_,s_r_80__43_,s_r_80__42_,s_r_80__41_,s_r_80__40_,
  s_r_80__39_,s_r_80__38_,s_r_80__37_,s_r_80__36_,s_r_80__35_,s_r_80__34_,
  s_r_80__33_,s_r_80__32_,s_r_80__31_,s_r_80__30_,s_r_80__29_,s_r_80__28_,s_r_80__27_,
  s_r_80__26_,s_r_80__25_,s_r_80__24_,s_r_80__23_,s_r_80__22_,s_r_80__21_,s_r_80__20_,
  s_r_80__19_,s_r_80__18_,s_r_80__17_,s_r_80__16_,s_r_80__15_,s_r_80__14_,
  s_r_80__13_,s_r_80__12_,s_r_80__11_,s_r_80__10_,s_r_80__9_,s_r_80__8_,s_r_80__7_,
  s_r_80__6_,s_r_80__5_,s_r_80__4_,s_r_80__3_,s_r_80__2_,s_r_80__1_,s_r_80__0_,
  s_r_79__127_,s_r_79__126_,s_r_79__125_,s_r_79__124_,s_r_79__123_,s_r_79__122_,
  s_r_79__121_,s_r_79__120_,s_r_79__119_,s_r_79__118_,s_r_79__117_,s_r_79__116_,s_r_79__115_,
  s_r_79__114_,s_r_79__113_,s_r_79__112_,s_r_79__111_,s_r_79__110_,s_r_79__109_,
  s_r_79__108_,s_r_79__107_,s_r_79__106_,s_r_79__105_,s_r_79__104_,s_r_79__103_,
  s_r_79__102_,s_r_79__101_,s_r_79__100_,s_r_79__99_,s_r_79__98_,s_r_79__97_,
  s_r_79__96_,s_r_79__95_,s_r_79__94_,s_r_79__93_,s_r_79__92_,s_r_79__91_,s_r_79__90_,
  s_r_79__89_,s_r_79__88_,s_r_79__87_,s_r_79__86_,s_r_79__85_,s_r_79__84_,s_r_79__83_,
  s_r_79__82_,s_r_79__81_,s_r_79__80_,s_r_79__79_,s_r_79__78_,s_r_79__77_,
  s_r_79__76_,s_r_79__75_,s_r_79__74_,s_r_79__73_,s_r_79__72_,s_r_79__71_,s_r_79__70_,
  s_r_79__69_,s_r_79__68_,s_r_79__67_,s_r_79__66_,s_r_79__65_,s_r_79__64_,s_r_79__63_,
  s_r_79__62_,s_r_79__61_,s_r_79__60_,s_r_79__59_,s_r_79__58_,s_r_79__57_,
  s_r_79__56_,s_r_79__55_,s_r_79__54_,s_r_79__53_,s_r_79__52_,s_r_79__51_,s_r_79__50_,
  s_r_79__49_,s_r_79__48_,s_r_79__47_,s_r_79__46_,s_r_79__45_,s_r_79__44_,s_r_79__43_,
  s_r_79__42_,s_r_79__41_,s_r_79__40_,s_r_79__39_,s_r_79__38_,s_r_79__37_,
  s_r_79__36_,s_r_79__35_,s_r_79__34_,s_r_79__33_,s_r_79__32_,s_r_79__31_,s_r_79__30_,
  s_r_79__29_,s_r_79__28_,s_r_79__27_,s_r_79__26_,s_r_79__25_,s_r_79__24_,s_r_79__23_,
  s_r_79__22_,s_r_79__21_,s_r_79__20_,s_r_79__19_,s_r_79__18_,s_r_79__17_,
  s_r_79__16_,s_r_79__15_,s_r_79__14_,s_r_79__13_,s_r_79__12_,s_r_79__11_,s_r_79__10_,
  s_r_79__9_,s_r_79__8_,s_r_79__7_,s_r_79__6_,s_r_79__5_,s_r_79__4_,s_r_79__3_,
  s_r_79__2_,s_r_79__1_,s_r_79__0_,prod_accum_82__83_,prod_accum_82__82_,
  prod_accum_82__81_,prod_accum_82__80_,prod_accum_82__79_,prod_accum_82__78_,prod_accum_82__77_,
  prod_accum_82__76_,prod_accum_82__75_,prod_accum_82__74_,prod_accum_82__73_,
  prod_accum_82__72_,prod_accum_82__71_,prod_accum_82__70_,prod_accum_82__69_,
  prod_accum_82__68_,prod_accum_82__67_,prod_accum_82__66_,prod_accum_82__65_,
  prod_accum_82__64_,prod_accum_82__63_,prod_accum_82__62_,prod_accum_82__61_,prod_accum_82__60_,
  prod_accum_82__59_,prod_accum_82__58_,prod_accum_82__57_,prod_accum_82__56_,
  prod_accum_82__55_,prod_accum_82__54_,prod_accum_82__53_,prod_accum_82__52_,
  prod_accum_82__51_,prod_accum_82__50_,prod_accum_82__49_,prod_accum_82__48_,
  prod_accum_82__47_,prod_accum_82__46_,prod_accum_82__45_,prod_accum_82__44_,
  prod_accum_82__43_,prod_accum_82__42_,prod_accum_82__41_,prod_accum_82__40_,prod_accum_82__39_,
  prod_accum_82__38_,prod_accum_82__37_,prod_accum_82__36_,prod_accum_82__35_,
  prod_accum_82__34_,prod_accum_82__33_,prod_accum_82__32_,prod_accum_82__31_,
  prod_accum_82__30_,prod_accum_82__29_,prod_accum_82__28_,prod_accum_82__27_,
  prod_accum_82__26_,prod_accum_82__25_,prod_accum_82__24_,prod_accum_82__23_,
  prod_accum_82__22_,prod_accum_82__21_,prod_accum_82__20_,prod_accum_82__19_,prod_accum_82__18_,
  prod_accum_82__17_,prod_accum_82__16_,prod_accum_82__15_,prod_accum_82__14_,
  prod_accum_82__13_,prod_accum_82__12_,prod_accum_82__11_,prod_accum_82__10_,
  prod_accum_82__9_,prod_accum_82__8_,prod_accum_82__7_,prod_accum_82__6_,prod_accum_82__5_,
  prod_accum_82__4_,prod_accum_82__3_,prod_accum_82__2_,prod_accum_82__1_,
  prod_accum_82__0_,prod_accum_81__82_,prod_accum_81__81_,prod_accum_81__80_,
  prod_accum_81__79_,prod_accum_81__78_,prod_accum_81__77_,prod_accum_81__76_,
  prod_accum_81__75_,prod_accum_81__74_,prod_accum_81__73_,prod_accum_81__72_,prod_accum_81__71_,
  prod_accum_81__70_,prod_accum_81__69_,prod_accum_81__68_,prod_accum_81__67_,
  prod_accum_81__66_,prod_accum_81__65_,prod_accum_81__64_,prod_accum_81__63_,
  prod_accum_81__62_,prod_accum_81__61_,prod_accum_81__60_,prod_accum_81__59_,
  prod_accum_81__58_,prod_accum_81__57_,prod_accum_81__56_,prod_accum_81__55_,
  prod_accum_81__54_,prod_accum_81__53_,prod_accum_81__52_,prod_accum_81__51_,prod_accum_81__50_,
  prod_accum_81__49_,prod_accum_81__48_,prod_accum_81__47_,prod_accum_81__46_,
  prod_accum_81__45_,prod_accum_81__44_,prod_accum_81__43_,prod_accum_81__42_,
  prod_accum_81__41_,prod_accum_81__40_,prod_accum_81__39_,prod_accum_81__38_,
  prod_accum_81__37_,prod_accum_81__36_,prod_accum_81__35_,prod_accum_81__34_,prod_accum_81__33_,
  prod_accum_81__32_,prod_accum_81__31_,prod_accum_81__30_,prod_accum_81__29_,
  prod_accum_81__28_,prod_accum_81__27_,prod_accum_81__26_,prod_accum_81__25_,
  prod_accum_81__24_,prod_accum_81__23_,prod_accum_81__22_,prod_accum_81__21_,
  prod_accum_81__20_,prod_accum_81__19_,prod_accum_81__18_,prod_accum_81__17_,
  prod_accum_81__16_,prod_accum_81__15_,prod_accum_81__14_,prod_accum_81__13_,prod_accum_81__12_,
  prod_accum_81__11_,prod_accum_81__10_,prod_accum_81__9_,prod_accum_81__8_,
  prod_accum_81__7_,prod_accum_81__6_,prod_accum_81__5_,prod_accum_81__4_,
  prod_accum_81__3_,prod_accum_81__2_,prod_accum_81__1_,prod_accum_81__0_,prod_accum_80__81_,
  prod_accum_80__80_,prod_accum_80__79_,prod_accum_80__78_,prod_accum_80__77_,
  prod_accum_80__76_,prod_accum_80__75_,prod_accum_80__74_,prod_accum_80__73_,
  prod_accum_80__72_,prod_accum_80__71_,prod_accum_80__70_,prod_accum_80__69_,
  prod_accum_80__68_,prod_accum_80__67_,prod_accum_80__66_,prod_accum_80__65_,prod_accum_80__64_,
  prod_accum_80__63_,prod_accum_80__62_,prod_accum_80__61_,prod_accum_80__60_,
  prod_accum_80__59_,prod_accum_80__58_,prod_accum_80__57_,prod_accum_80__56_,
  prod_accum_80__55_,prod_accum_80__54_,prod_accum_80__53_,prod_accum_80__52_,
  prod_accum_80__51_,prod_accum_80__50_,prod_accum_80__49_,prod_accum_80__48_,
  prod_accum_80__47_,prod_accum_80__46_,prod_accum_80__45_,prod_accum_80__44_,prod_accum_80__43_,
  prod_accum_80__42_,prod_accum_80__41_,prod_accum_80__40_,prod_accum_80__39_,
  prod_accum_80__38_,prod_accum_80__37_,prod_accum_80__36_,prod_accum_80__35_,
  prod_accum_80__34_,prod_accum_80__33_,prod_accum_80__32_,prod_accum_80__31_,
  prod_accum_80__30_,prod_accum_80__29_,prod_accum_80__28_,prod_accum_80__27_,
  prod_accum_80__26_,prod_accum_80__25_,prod_accum_80__24_,prod_accum_80__23_,prod_accum_80__22_,
  prod_accum_80__21_,prod_accum_80__20_,prod_accum_80__19_,prod_accum_80__18_,
  prod_accum_80__17_,prod_accum_80__16_,prod_accum_80__15_,prod_accum_80__14_,
  prod_accum_80__13_,prod_accum_80__12_,prod_accum_80__11_,prod_accum_80__10_,
  prod_accum_80__9_,prod_accum_80__8_,prod_accum_80__7_,prod_accum_80__6_,prod_accum_80__5_,
  prod_accum_80__4_,prod_accum_80__3_,prod_accum_80__2_,prod_accum_80__1_,
  prod_accum_80__0_,prod_accum_79__80_,prod_accum_79__79_,prod_accum_79__78_,
  prod_accum_79__77_,prod_accum_79__76_,prod_accum_79__75_,prod_accum_79__74_,prod_accum_79__73_,
  prod_accum_79__72_,prod_accum_79__71_,prod_accum_79__70_,prod_accum_79__69_,
  prod_accum_79__68_,prod_accum_79__67_,prod_accum_79__66_,prod_accum_79__65_,
  prod_accum_79__64_,prod_accum_79__63_,prod_accum_79__62_,prod_accum_79__61_,
  prod_accum_79__60_,prod_accum_79__59_,prod_accum_79__58_,prod_accum_79__57_,prod_accum_79__56_,
  prod_accum_79__55_,prod_accum_79__54_,prod_accum_79__53_,prod_accum_79__52_,
  prod_accum_79__51_,prod_accum_79__50_,prod_accum_79__49_,prod_accum_79__48_,
  prod_accum_79__47_,prod_accum_79__46_,prod_accum_79__45_,prod_accum_79__44_,
  prod_accum_79__43_,prod_accum_79__42_,prod_accum_79__41_,prod_accum_79__40_,
  prod_accum_79__39_,prod_accum_79__38_,prod_accum_79__37_,prod_accum_79__36_,prod_accum_79__35_,
  prod_accum_79__34_,prod_accum_79__33_,prod_accum_79__32_,prod_accum_79__31_,
  prod_accum_79__30_,prod_accum_79__29_,prod_accum_79__28_,prod_accum_79__27_,
  prod_accum_79__26_,prod_accum_79__25_,prod_accum_79__24_,prod_accum_79__23_,
  prod_accum_79__22_,prod_accum_79__21_,prod_accum_79__20_,prod_accum_79__19_,
  prod_accum_79__18_,prod_accum_79__17_,prod_accum_79__16_,prod_accum_79__15_,prod_accum_79__14_,
  prod_accum_79__13_,prod_accum_79__12_,prod_accum_79__11_,prod_accum_79__10_,
  prod_accum_79__9_,prod_accum_79__8_,prod_accum_79__7_,prod_accum_79__6_,
  prod_accum_79__5_,prod_accum_79__4_,prod_accum_79__3_,prod_accum_79__2_,prod_accum_79__1_,
  prod_accum_79__0_,s_r_86__127_,s_r_86__126_,s_r_86__125_,s_r_86__124_,s_r_86__123_,
  s_r_86__122_,s_r_86__121_,s_r_86__120_,s_r_86__119_,s_r_86__118_,s_r_86__117_,
  s_r_86__116_,s_r_86__115_,s_r_86__114_,s_r_86__113_,s_r_86__112_,s_r_86__111_,
  s_r_86__110_,s_r_86__109_,s_r_86__108_,s_r_86__107_,s_r_86__106_,s_r_86__105_,
  s_r_86__104_,s_r_86__103_,s_r_86__102_,s_r_86__101_,s_r_86__100_,s_r_86__99_,
  s_r_86__98_,s_r_86__97_,s_r_86__96_,s_r_86__95_,s_r_86__94_,s_r_86__93_,s_r_86__92_,
  s_r_86__91_,s_r_86__90_,s_r_86__89_,s_r_86__88_,s_r_86__87_,s_r_86__86_,s_r_86__85_,
  s_r_86__84_,s_r_86__83_,s_r_86__82_,s_r_86__81_,s_r_86__80_,s_r_86__79_,
  s_r_86__78_,s_r_86__77_,s_r_86__76_,s_r_86__75_,s_r_86__74_,s_r_86__73_,s_r_86__72_,
  s_r_86__71_,s_r_86__70_,s_r_86__69_,s_r_86__68_,s_r_86__67_,s_r_86__66_,s_r_86__65_,
  s_r_86__64_,s_r_86__63_,s_r_86__62_,s_r_86__61_,s_r_86__60_,s_r_86__59_,
  s_r_86__58_,s_r_86__57_,s_r_86__56_,s_r_86__55_,s_r_86__54_,s_r_86__53_,s_r_86__52_,
  s_r_86__51_,s_r_86__50_,s_r_86__49_,s_r_86__48_,s_r_86__47_,s_r_86__46_,s_r_86__45_,
  s_r_86__44_,s_r_86__43_,s_r_86__42_,s_r_86__41_,s_r_86__40_,s_r_86__39_,
  s_r_86__38_,s_r_86__37_,s_r_86__36_,s_r_86__35_,s_r_86__34_,s_r_86__33_,s_r_86__32_,
  s_r_86__31_,s_r_86__30_,s_r_86__29_,s_r_86__28_,s_r_86__27_,s_r_86__26_,s_r_86__25_,
  s_r_86__24_,s_r_86__23_,s_r_86__22_,s_r_86__21_,s_r_86__20_,s_r_86__19_,
  s_r_86__18_,s_r_86__17_,s_r_86__16_,s_r_86__15_,s_r_86__14_,s_r_86__13_,s_r_86__12_,
  s_r_86__11_,s_r_86__10_,s_r_86__9_,s_r_86__8_,s_r_86__7_,s_r_86__6_,s_r_86__5_,
  s_r_86__4_,s_r_86__3_,s_r_86__2_,s_r_86__1_,s_r_86__0_,s_r_85__127_,s_r_85__126_,
  s_r_85__125_,s_r_85__124_,s_r_85__123_,s_r_85__122_,s_r_85__121_,s_r_85__120_,
  s_r_85__119_,s_r_85__118_,s_r_85__117_,s_r_85__116_,s_r_85__115_,s_r_85__114_,
  s_r_85__113_,s_r_85__112_,s_r_85__111_,s_r_85__110_,s_r_85__109_,s_r_85__108_,
  s_r_85__107_,s_r_85__106_,s_r_85__105_,s_r_85__104_,s_r_85__103_,s_r_85__102_,s_r_85__101_,
  s_r_85__100_,s_r_85__99_,s_r_85__98_,s_r_85__97_,s_r_85__96_,s_r_85__95_,
  s_r_85__94_,s_r_85__93_,s_r_85__92_,s_r_85__91_,s_r_85__90_,s_r_85__89_,s_r_85__88_,
  s_r_85__87_,s_r_85__86_,s_r_85__85_,s_r_85__84_,s_r_85__83_,s_r_85__82_,s_r_85__81_,
  s_r_85__80_,s_r_85__79_,s_r_85__78_,s_r_85__77_,s_r_85__76_,s_r_85__75_,
  s_r_85__74_,s_r_85__73_,s_r_85__72_,s_r_85__71_,s_r_85__70_,s_r_85__69_,s_r_85__68_,
  s_r_85__67_,s_r_85__66_,s_r_85__65_,s_r_85__64_,s_r_85__63_,s_r_85__62_,s_r_85__61_,
  s_r_85__60_,s_r_85__59_,s_r_85__58_,s_r_85__57_,s_r_85__56_,s_r_85__55_,
  s_r_85__54_,s_r_85__53_,s_r_85__52_,s_r_85__51_,s_r_85__50_,s_r_85__49_,s_r_85__48_,
  s_r_85__47_,s_r_85__46_,s_r_85__45_,s_r_85__44_,s_r_85__43_,s_r_85__42_,s_r_85__41_,
  s_r_85__40_,s_r_85__39_,s_r_85__38_,s_r_85__37_,s_r_85__36_,s_r_85__35_,
  s_r_85__34_,s_r_85__33_,s_r_85__32_,s_r_85__31_,s_r_85__30_,s_r_85__29_,s_r_85__28_,
  s_r_85__27_,s_r_85__26_,s_r_85__25_,s_r_85__24_,s_r_85__23_,s_r_85__22_,s_r_85__21_,
  s_r_85__20_,s_r_85__19_,s_r_85__18_,s_r_85__17_,s_r_85__16_,s_r_85__15_,
  s_r_85__14_,s_r_85__13_,s_r_85__12_,s_r_85__11_,s_r_85__10_,s_r_85__9_,s_r_85__8_,
  s_r_85__7_,s_r_85__6_,s_r_85__5_,s_r_85__4_,s_r_85__3_,s_r_85__2_,s_r_85__1_,
  s_r_85__0_,s_r_84__127_,s_r_84__126_,s_r_84__125_,s_r_84__124_,s_r_84__123_,s_r_84__122_,
  s_r_84__121_,s_r_84__120_,s_r_84__119_,s_r_84__118_,s_r_84__117_,s_r_84__116_,
  s_r_84__115_,s_r_84__114_,s_r_84__113_,s_r_84__112_,s_r_84__111_,s_r_84__110_,
  s_r_84__109_,s_r_84__108_,s_r_84__107_,s_r_84__106_,s_r_84__105_,s_r_84__104_,
  s_r_84__103_,s_r_84__102_,s_r_84__101_,s_r_84__100_,s_r_84__99_,s_r_84__98_,
  s_r_84__97_,s_r_84__96_,s_r_84__95_,s_r_84__94_,s_r_84__93_,s_r_84__92_,s_r_84__91_,
  s_r_84__90_,s_r_84__89_,s_r_84__88_,s_r_84__87_,s_r_84__86_,s_r_84__85_,s_r_84__84_,
  s_r_84__83_,s_r_84__82_,s_r_84__81_,s_r_84__80_,s_r_84__79_,s_r_84__78_,
  s_r_84__77_,s_r_84__76_,s_r_84__75_,s_r_84__74_,s_r_84__73_,s_r_84__72_,s_r_84__71_,
  s_r_84__70_,s_r_84__69_,s_r_84__68_,s_r_84__67_,s_r_84__66_,s_r_84__65_,s_r_84__64_,
  s_r_84__63_,s_r_84__62_,s_r_84__61_,s_r_84__60_,s_r_84__59_,s_r_84__58_,
  s_r_84__57_,s_r_84__56_,s_r_84__55_,s_r_84__54_,s_r_84__53_,s_r_84__52_,s_r_84__51_,
  s_r_84__50_,s_r_84__49_,s_r_84__48_,s_r_84__47_,s_r_84__46_,s_r_84__45_,s_r_84__44_,
  s_r_84__43_,s_r_84__42_,s_r_84__41_,s_r_84__40_,s_r_84__39_,s_r_84__38_,
  s_r_84__37_,s_r_84__36_,s_r_84__35_,s_r_84__34_,s_r_84__33_,s_r_84__32_,s_r_84__31_,
  s_r_84__30_,s_r_84__29_,s_r_84__28_,s_r_84__27_,s_r_84__26_,s_r_84__25_,s_r_84__24_,
  s_r_84__23_,s_r_84__22_,s_r_84__21_,s_r_84__20_,s_r_84__19_,s_r_84__18_,
  s_r_84__17_,s_r_84__16_,s_r_84__15_,s_r_84__14_,s_r_84__13_,s_r_84__12_,s_r_84__11_,
  s_r_84__10_,s_r_84__9_,s_r_84__8_,s_r_84__7_,s_r_84__6_,s_r_84__5_,s_r_84__4_,
  s_r_84__3_,s_r_84__2_,s_r_84__1_,s_r_84__0_,s_r_83__127_,s_r_83__126_,s_r_83__125_,
  s_r_83__124_,s_r_83__123_,s_r_83__122_,s_r_83__121_,s_r_83__120_,s_r_83__119_,
  s_r_83__118_,s_r_83__117_,s_r_83__116_,s_r_83__115_,s_r_83__114_,s_r_83__113_,
  s_r_83__112_,s_r_83__111_,s_r_83__110_,s_r_83__109_,s_r_83__108_,s_r_83__107_,
  s_r_83__106_,s_r_83__105_,s_r_83__104_,s_r_83__103_,s_r_83__102_,s_r_83__101_,s_r_83__100_,
  s_r_83__99_,s_r_83__98_,s_r_83__97_,s_r_83__96_,s_r_83__95_,s_r_83__94_,
  s_r_83__93_,s_r_83__92_,s_r_83__91_,s_r_83__90_,s_r_83__89_,s_r_83__88_,s_r_83__87_,
  s_r_83__86_,s_r_83__85_,s_r_83__84_,s_r_83__83_,s_r_83__82_,s_r_83__81_,s_r_83__80_,
  s_r_83__79_,s_r_83__78_,s_r_83__77_,s_r_83__76_,s_r_83__75_,s_r_83__74_,
  s_r_83__73_,s_r_83__72_,s_r_83__71_,s_r_83__70_,s_r_83__69_,s_r_83__68_,s_r_83__67_,
  s_r_83__66_,s_r_83__65_,s_r_83__64_,s_r_83__63_,s_r_83__62_,s_r_83__61_,s_r_83__60_,
  s_r_83__59_,s_r_83__58_,s_r_83__57_,s_r_83__56_,s_r_83__55_,s_r_83__54_,
  s_r_83__53_,s_r_83__52_,s_r_83__51_,s_r_83__50_,s_r_83__49_,s_r_83__48_,s_r_83__47_,
  s_r_83__46_,s_r_83__45_,s_r_83__44_,s_r_83__43_,s_r_83__42_,s_r_83__41_,s_r_83__40_,
  s_r_83__39_,s_r_83__38_,s_r_83__37_,s_r_83__36_,s_r_83__35_,s_r_83__34_,
  s_r_83__33_,s_r_83__32_,s_r_83__31_,s_r_83__30_,s_r_83__29_,s_r_83__28_,s_r_83__27_,
  s_r_83__26_,s_r_83__25_,s_r_83__24_,s_r_83__23_,s_r_83__22_,s_r_83__21_,s_r_83__20_,
  s_r_83__19_,s_r_83__18_,s_r_83__17_,s_r_83__16_,s_r_83__15_,s_r_83__14_,
  s_r_83__13_,s_r_83__12_,s_r_83__11_,s_r_83__10_,s_r_83__9_,s_r_83__8_,s_r_83__7_,
  s_r_83__6_,s_r_83__5_,s_r_83__4_,s_r_83__3_,s_r_83__2_,s_r_83__1_,s_r_83__0_,
  prod_accum_86__87_,prod_accum_86__86_,prod_accum_86__85_,prod_accum_86__84_,
  prod_accum_86__83_,prod_accum_86__82_,prod_accum_86__81_,prod_accum_86__80_,
  prod_accum_86__79_,prod_accum_86__78_,prod_accum_86__77_,prod_accum_86__76_,prod_accum_86__75_,
  prod_accum_86__74_,prod_accum_86__73_,prod_accum_86__72_,prod_accum_86__71_,
  prod_accum_86__70_,prod_accum_86__69_,prod_accum_86__68_,prod_accum_86__67_,
  prod_accum_86__66_,prod_accum_86__65_,prod_accum_86__64_,prod_accum_86__63_,
  prod_accum_86__62_,prod_accum_86__61_,prod_accum_86__60_,prod_accum_86__59_,prod_accum_86__58_,
  prod_accum_86__57_,prod_accum_86__56_,prod_accum_86__55_,prod_accum_86__54_,
  prod_accum_86__53_,prod_accum_86__52_,prod_accum_86__51_,prod_accum_86__50_,
  prod_accum_86__49_,prod_accum_86__48_,prod_accum_86__47_,prod_accum_86__46_,
  prod_accum_86__45_,prod_accum_86__44_,prod_accum_86__43_,prod_accum_86__42_,
  prod_accum_86__41_,prod_accum_86__40_,prod_accum_86__39_,prod_accum_86__38_,prod_accum_86__37_,
  prod_accum_86__36_,prod_accum_86__35_,prod_accum_86__34_,prod_accum_86__33_,
  prod_accum_86__32_,prod_accum_86__31_,prod_accum_86__30_,prod_accum_86__29_,
  prod_accum_86__28_,prod_accum_86__27_,prod_accum_86__26_,prod_accum_86__25_,
  prod_accum_86__24_,prod_accum_86__23_,prod_accum_86__22_,prod_accum_86__21_,
  prod_accum_86__20_,prod_accum_86__19_,prod_accum_86__18_,prod_accum_86__17_,prod_accum_86__16_,
  prod_accum_86__15_,prod_accum_86__14_,prod_accum_86__13_,prod_accum_86__12_,
  prod_accum_86__11_,prod_accum_86__10_,prod_accum_86__9_,prod_accum_86__8_,
  prod_accum_86__7_,prod_accum_86__6_,prod_accum_86__5_,prod_accum_86__4_,prod_accum_86__3_,
  prod_accum_86__2_,prod_accum_86__1_,prod_accum_86__0_,prod_accum_85__86_,
  prod_accum_85__85_,prod_accum_85__84_,prod_accum_85__83_,prod_accum_85__82_,
  prod_accum_85__81_,prod_accum_85__80_,prod_accum_85__79_,prod_accum_85__78_,
  prod_accum_85__77_,prod_accum_85__76_,prod_accum_85__75_,prod_accum_85__74_,prod_accum_85__73_,
  prod_accum_85__72_,prod_accum_85__71_,prod_accum_85__70_,prod_accum_85__69_,
  prod_accum_85__68_,prod_accum_85__67_,prod_accum_85__66_,prod_accum_85__65_,
  prod_accum_85__64_,prod_accum_85__63_,prod_accum_85__62_,prod_accum_85__61_,
  prod_accum_85__60_,prod_accum_85__59_,prod_accum_85__58_,prod_accum_85__57_,
  prod_accum_85__56_,prod_accum_85__55_,prod_accum_85__54_,prod_accum_85__53_,prod_accum_85__52_,
  prod_accum_85__51_,prod_accum_85__50_,prod_accum_85__49_,prod_accum_85__48_,
  prod_accum_85__47_,prod_accum_85__46_,prod_accum_85__45_,prod_accum_85__44_,
  prod_accum_85__43_,prod_accum_85__42_,prod_accum_85__41_,prod_accum_85__40_,
  prod_accum_85__39_,prod_accum_85__38_,prod_accum_85__37_,prod_accum_85__36_,prod_accum_85__35_,
  prod_accum_85__34_,prod_accum_85__33_,prod_accum_85__32_,prod_accum_85__31_,
  prod_accum_85__30_,prod_accum_85__29_,prod_accum_85__28_,prod_accum_85__27_,
  prod_accum_85__26_,prod_accum_85__25_,prod_accum_85__24_,prod_accum_85__23_,
  prod_accum_85__22_,prod_accum_85__21_,prod_accum_85__20_,prod_accum_85__19_,
  prod_accum_85__18_,prod_accum_85__17_,prod_accum_85__16_,prod_accum_85__15_,prod_accum_85__14_,
  prod_accum_85__13_,prod_accum_85__12_,prod_accum_85__11_,prod_accum_85__10_,
  prod_accum_85__9_,prod_accum_85__8_,prod_accum_85__7_,prod_accum_85__6_,
  prod_accum_85__5_,prod_accum_85__4_,prod_accum_85__3_,prod_accum_85__2_,prod_accum_85__1_,
  prod_accum_85__0_,prod_accum_84__85_,prod_accum_84__84_,prod_accum_84__83_,
  prod_accum_84__82_,prod_accum_84__81_,prod_accum_84__80_,prod_accum_84__79_,
  prod_accum_84__78_,prod_accum_84__77_,prod_accum_84__76_,prod_accum_84__75_,
  prod_accum_84__74_,prod_accum_84__73_,prod_accum_84__72_,prod_accum_84__71_,prod_accum_84__70_,
  prod_accum_84__69_,prod_accum_84__68_,prod_accum_84__67_,prod_accum_84__66_,
  prod_accum_84__65_,prod_accum_84__64_,prod_accum_84__63_,prod_accum_84__62_,
  prod_accum_84__61_,prod_accum_84__60_,prod_accum_84__59_,prod_accum_84__58_,
  prod_accum_84__57_,prod_accum_84__56_,prod_accum_84__55_,prod_accum_84__54_,
  prod_accum_84__53_,prod_accum_84__52_,prod_accum_84__51_,prod_accum_84__50_,prod_accum_84__49_,
  prod_accum_84__48_,prod_accum_84__47_,prod_accum_84__46_,prod_accum_84__45_,
  prod_accum_84__44_,prod_accum_84__43_,prod_accum_84__42_,prod_accum_84__41_,
  prod_accum_84__40_,prod_accum_84__39_,prod_accum_84__38_,prod_accum_84__37_,
  prod_accum_84__36_,prod_accum_84__35_,prod_accum_84__34_,prod_accum_84__33_,
  prod_accum_84__32_,prod_accum_84__31_,prod_accum_84__30_,prod_accum_84__29_,prod_accum_84__28_,
  prod_accum_84__27_,prod_accum_84__26_,prod_accum_84__25_,prod_accum_84__24_,
  prod_accum_84__23_,prod_accum_84__22_,prod_accum_84__21_,prod_accum_84__20_,
  prod_accum_84__19_,prod_accum_84__18_,prod_accum_84__17_,prod_accum_84__16_,
  prod_accum_84__15_,prod_accum_84__14_,prod_accum_84__13_,prod_accum_84__12_,prod_accum_84__11_,
  prod_accum_84__10_,prod_accum_84__9_,prod_accum_84__8_,prod_accum_84__7_,
  prod_accum_84__6_,prod_accum_84__5_,prod_accum_84__4_,prod_accum_84__3_,
  prod_accum_84__2_,prod_accum_84__1_,prod_accum_84__0_,prod_accum_83__84_,prod_accum_83__83_,
  prod_accum_83__82_,prod_accum_83__81_,prod_accum_83__80_,prod_accum_83__79_,
  prod_accum_83__78_,prod_accum_83__77_,prod_accum_83__76_,prod_accum_83__75_,
  prod_accum_83__74_,prod_accum_83__73_,prod_accum_83__72_,prod_accum_83__71_,
  prod_accum_83__70_,prod_accum_83__69_,prod_accum_83__68_,prod_accum_83__67_,prod_accum_83__66_,
  prod_accum_83__65_,prod_accum_83__64_,prod_accum_83__63_,prod_accum_83__62_,
  prod_accum_83__61_,prod_accum_83__60_,prod_accum_83__59_,prod_accum_83__58_,
  prod_accum_83__57_,prod_accum_83__56_,prod_accum_83__55_,prod_accum_83__54_,
  prod_accum_83__53_,prod_accum_83__52_,prod_accum_83__51_,prod_accum_83__50_,
  prod_accum_83__49_,prod_accum_83__48_,prod_accum_83__47_,prod_accum_83__46_,prod_accum_83__45_,
  prod_accum_83__44_,prod_accum_83__43_,prod_accum_83__42_,prod_accum_83__41_,
  prod_accum_83__40_,prod_accum_83__39_,prod_accum_83__38_,prod_accum_83__37_,
  prod_accum_83__36_,prod_accum_83__35_,prod_accum_83__34_,prod_accum_83__33_,
  prod_accum_83__32_,prod_accum_83__31_,prod_accum_83__30_,prod_accum_83__29_,
  prod_accum_83__28_,prod_accum_83__27_,prod_accum_83__26_,prod_accum_83__25_,prod_accum_83__24_,
  prod_accum_83__23_,prod_accum_83__22_,prod_accum_83__21_,prod_accum_83__20_,
  prod_accum_83__19_,prod_accum_83__18_,prod_accum_83__17_,prod_accum_83__16_,
  prod_accum_83__15_,prod_accum_83__14_,prod_accum_83__13_,prod_accum_83__12_,
  prod_accum_83__11_,prod_accum_83__10_,prod_accum_83__9_,prod_accum_83__8_,prod_accum_83__7_,
  prod_accum_83__6_,prod_accum_83__5_,prod_accum_83__4_,prod_accum_83__3_,
  prod_accum_83__2_,prod_accum_83__1_,prod_accum_83__0_,s_r_90__127_,s_r_90__126_,
  s_r_90__125_,s_r_90__124_,s_r_90__123_,s_r_90__122_,s_r_90__121_,s_r_90__120_,
  s_r_90__119_,s_r_90__118_,s_r_90__117_,s_r_90__116_,s_r_90__115_,s_r_90__114_,s_r_90__113_,
  s_r_90__112_,s_r_90__111_,s_r_90__110_,s_r_90__109_,s_r_90__108_,s_r_90__107_,
  s_r_90__106_,s_r_90__105_,s_r_90__104_,s_r_90__103_,s_r_90__102_,s_r_90__101_,
  s_r_90__100_,s_r_90__99_,s_r_90__98_,s_r_90__97_,s_r_90__96_,s_r_90__95_,s_r_90__94_,
  s_r_90__93_,s_r_90__92_,s_r_90__91_,s_r_90__90_,s_r_90__89_,s_r_90__88_,
  s_r_90__87_,s_r_90__86_,s_r_90__85_,s_r_90__84_,s_r_90__83_,s_r_90__82_,s_r_90__81_,
  s_r_90__80_,s_r_90__79_,s_r_90__78_,s_r_90__77_,s_r_90__76_,s_r_90__75_,s_r_90__74_,
  s_r_90__73_,s_r_90__72_,s_r_90__71_,s_r_90__70_,s_r_90__69_,s_r_90__68_,
  s_r_90__67_,s_r_90__66_,s_r_90__65_,s_r_90__64_,s_r_90__63_,s_r_90__62_,s_r_90__61_,
  s_r_90__60_,s_r_90__59_,s_r_90__58_,s_r_90__57_,s_r_90__56_,s_r_90__55_,s_r_90__54_,
  s_r_90__53_,s_r_90__52_,s_r_90__51_,s_r_90__50_,s_r_90__49_,s_r_90__48_,
  s_r_90__47_,s_r_90__46_,s_r_90__45_,s_r_90__44_,s_r_90__43_,s_r_90__42_,s_r_90__41_,
  s_r_90__40_,s_r_90__39_,s_r_90__38_,s_r_90__37_,s_r_90__36_,s_r_90__35_,s_r_90__34_,
  s_r_90__33_,s_r_90__32_,s_r_90__31_,s_r_90__30_,s_r_90__29_,s_r_90__28_,
  s_r_90__27_,s_r_90__26_,s_r_90__25_,s_r_90__24_,s_r_90__23_,s_r_90__22_,s_r_90__21_,
  s_r_90__20_,s_r_90__19_,s_r_90__18_,s_r_90__17_,s_r_90__16_,s_r_90__15_,s_r_90__14_,
  s_r_90__13_,s_r_90__12_,s_r_90__11_,s_r_90__10_,s_r_90__9_,s_r_90__8_,
  s_r_90__7_,s_r_90__6_,s_r_90__5_,s_r_90__4_,s_r_90__3_,s_r_90__2_,s_r_90__1_,s_r_90__0_,
  s_r_89__127_,s_r_89__126_,s_r_89__125_,s_r_89__124_,s_r_89__123_,s_r_89__122_,
  s_r_89__121_,s_r_89__120_,s_r_89__119_,s_r_89__118_,s_r_89__117_,s_r_89__116_,
  s_r_89__115_,s_r_89__114_,s_r_89__113_,s_r_89__112_,s_r_89__111_,s_r_89__110_,
  s_r_89__109_,s_r_89__108_,s_r_89__107_,s_r_89__106_,s_r_89__105_,s_r_89__104_,
  s_r_89__103_,s_r_89__102_,s_r_89__101_,s_r_89__100_,s_r_89__99_,s_r_89__98_,s_r_89__97_,
  s_r_89__96_,s_r_89__95_,s_r_89__94_,s_r_89__93_,s_r_89__92_,s_r_89__91_,
  s_r_89__90_,s_r_89__89_,s_r_89__88_,s_r_89__87_,s_r_89__86_,s_r_89__85_,s_r_89__84_,
  s_r_89__83_,s_r_89__82_,s_r_89__81_,s_r_89__80_,s_r_89__79_,s_r_89__78_,s_r_89__77_,
  s_r_89__76_,s_r_89__75_,s_r_89__74_,s_r_89__73_,s_r_89__72_,s_r_89__71_,
  s_r_89__70_,s_r_89__69_,s_r_89__68_,s_r_89__67_,s_r_89__66_,s_r_89__65_,s_r_89__64_,
  s_r_89__63_,s_r_89__62_,s_r_89__61_,s_r_89__60_,s_r_89__59_,s_r_89__58_,s_r_89__57_,
  s_r_89__56_,s_r_89__55_,s_r_89__54_,s_r_89__53_,s_r_89__52_,s_r_89__51_,
  s_r_89__50_,s_r_89__49_,s_r_89__48_,s_r_89__47_,s_r_89__46_,s_r_89__45_,s_r_89__44_,
  s_r_89__43_,s_r_89__42_,s_r_89__41_,s_r_89__40_,s_r_89__39_,s_r_89__38_,s_r_89__37_,
  s_r_89__36_,s_r_89__35_,s_r_89__34_,s_r_89__33_,s_r_89__32_,s_r_89__31_,
  s_r_89__30_,s_r_89__29_,s_r_89__28_,s_r_89__27_,s_r_89__26_,s_r_89__25_,s_r_89__24_,
  s_r_89__23_,s_r_89__22_,s_r_89__21_,s_r_89__20_,s_r_89__19_,s_r_89__18_,s_r_89__17_,
  s_r_89__16_,s_r_89__15_,s_r_89__14_,s_r_89__13_,s_r_89__12_,s_r_89__11_,
  s_r_89__10_,s_r_89__9_,s_r_89__8_,s_r_89__7_,s_r_89__6_,s_r_89__5_,s_r_89__4_,s_r_89__3_,
  s_r_89__2_,s_r_89__1_,s_r_89__0_,s_r_88__127_,s_r_88__126_,s_r_88__125_,
  s_r_88__124_,s_r_88__123_,s_r_88__122_,s_r_88__121_,s_r_88__120_,s_r_88__119_,
  s_r_88__118_,s_r_88__117_,s_r_88__116_,s_r_88__115_,s_r_88__114_,s_r_88__113_,s_r_88__112_,
  s_r_88__111_,s_r_88__110_,s_r_88__109_,s_r_88__108_,s_r_88__107_,s_r_88__106_,
  s_r_88__105_,s_r_88__104_,s_r_88__103_,s_r_88__102_,s_r_88__101_,s_r_88__100_,
  s_r_88__99_,s_r_88__98_,s_r_88__97_,s_r_88__96_,s_r_88__95_,s_r_88__94_,s_r_88__93_,
  s_r_88__92_,s_r_88__91_,s_r_88__90_,s_r_88__89_,s_r_88__88_,s_r_88__87_,
  s_r_88__86_,s_r_88__85_,s_r_88__84_,s_r_88__83_,s_r_88__82_,s_r_88__81_,s_r_88__80_,
  s_r_88__79_,s_r_88__78_,s_r_88__77_,s_r_88__76_,s_r_88__75_,s_r_88__74_,s_r_88__73_,
  s_r_88__72_,s_r_88__71_,s_r_88__70_,s_r_88__69_,s_r_88__68_,s_r_88__67_,
  s_r_88__66_,s_r_88__65_,s_r_88__64_,s_r_88__63_,s_r_88__62_,s_r_88__61_,s_r_88__60_,
  s_r_88__59_,s_r_88__58_,s_r_88__57_,s_r_88__56_,s_r_88__55_,s_r_88__54_,s_r_88__53_,
  s_r_88__52_,s_r_88__51_,s_r_88__50_,s_r_88__49_,s_r_88__48_,s_r_88__47_,
  s_r_88__46_,s_r_88__45_,s_r_88__44_,s_r_88__43_,s_r_88__42_,s_r_88__41_,s_r_88__40_,
  s_r_88__39_,s_r_88__38_,s_r_88__37_,s_r_88__36_,s_r_88__35_,s_r_88__34_,s_r_88__33_,
  s_r_88__32_,s_r_88__31_,s_r_88__30_,s_r_88__29_,s_r_88__28_,s_r_88__27_,
  s_r_88__26_,s_r_88__25_,s_r_88__24_,s_r_88__23_,s_r_88__22_,s_r_88__21_,s_r_88__20_,
  s_r_88__19_,s_r_88__18_,s_r_88__17_,s_r_88__16_,s_r_88__15_,s_r_88__14_,s_r_88__13_,
  s_r_88__12_,s_r_88__11_,s_r_88__10_,s_r_88__9_,s_r_88__8_,s_r_88__7_,s_r_88__6_,
  s_r_88__5_,s_r_88__4_,s_r_88__3_,s_r_88__2_,s_r_88__1_,s_r_88__0_,s_r_87__127_,
  s_r_87__126_,s_r_87__125_,s_r_87__124_,s_r_87__123_,s_r_87__122_,s_r_87__121_,
  s_r_87__120_,s_r_87__119_,s_r_87__118_,s_r_87__117_,s_r_87__116_,s_r_87__115_,
  s_r_87__114_,s_r_87__113_,s_r_87__112_,s_r_87__111_,s_r_87__110_,s_r_87__109_,
  s_r_87__108_,s_r_87__107_,s_r_87__106_,s_r_87__105_,s_r_87__104_,s_r_87__103_,
  s_r_87__102_,s_r_87__101_,s_r_87__100_,s_r_87__99_,s_r_87__98_,s_r_87__97_,s_r_87__96_,
  s_r_87__95_,s_r_87__94_,s_r_87__93_,s_r_87__92_,s_r_87__91_,s_r_87__90_,
  s_r_87__89_,s_r_87__88_,s_r_87__87_,s_r_87__86_,s_r_87__85_,s_r_87__84_,s_r_87__83_,
  s_r_87__82_,s_r_87__81_,s_r_87__80_,s_r_87__79_,s_r_87__78_,s_r_87__77_,s_r_87__76_,
  s_r_87__75_,s_r_87__74_,s_r_87__73_,s_r_87__72_,s_r_87__71_,s_r_87__70_,
  s_r_87__69_,s_r_87__68_,s_r_87__67_,s_r_87__66_,s_r_87__65_,s_r_87__64_,s_r_87__63_,
  s_r_87__62_,s_r_87__61_,s_r_87__60_,s_r_87__59_,s_r_87__58_,s_r_87__57_,s_r_87__56_,
  s_r_87__55_,s_r_87__54_,s_r_87__53_,s_r_87__52_,s_r_87__51_,s_r_87__50_,
  s_r_87__49_,s_r_87__48_,s_r_87__47_,s_r_87__46_,s_r_87__45_,s_r_87__44_,s_r_87__43_,
  s_r_87__42_,s_r_87__41_,s_r_87__40_,s_r_87__39_,s_r_87__38_,s_r_87__37_,s_r_87__36_,
  s_r_87__35_,s_r_87__34_,s_r_87__33_,s_r_87__32_,s_r_87__31_,s_r_87__30_,
  s_r_87__29_,s_r_87__28_,s_r_87__27_,s_r_87__26_,s_r_87__25_,s_r_87__24_,s_r_87__23_,
  s_r_87__22_,s_r_87__21_,s_r_87__20_,s_r_87__19_,s_r_87__18_,s_r_87__17_,s_r_87__16_,
  s_r_87__15_,s_r_87__14_,s_r_87__13_,s_r_87__12_,s_r_87__11_,s_r_87__10_,
  s_r_87__9_,s_r_87__8_,s_r_87__7_,s_r_87__6_,s_r_87__5_,s_r_87__4_,s_r_87__3_,s_r_87__2_,
  s_r_87__1_,s_r_87__0_,prod_accum_90__91_,prod_accum_90__90_,prod_accum_90__89_,
  prod_accum_90__88_,prod_accum_90__87_,prod_accum_90__86_,prod_accum_90__85_,
  prod_accum_90__84_,prod_accum_90__83_,prod_accum_90__82_,prod_accum_90__81_,
  prod_accum_90__80_,prod_accum_90__79_,prod_accum_90__78_,prod_accum_90__77_,
  prod_accum_90__76_,prod_accum_90__75_,prod_accum_90__74_,prod_accum_90__73_,prod_accum_90__72_,
  prod_accum_90__71_,prod_accum_90__70_,prod_accum_90__69_,prod_accum_90__68_,
  prod_accum_90__67_,prod_accum_90__66_,prod_accum_90__65_,prod_accum_90__64_,
  prod_accum_90__63_,prod_accum_90__62_,prod_accum_90__61_,prod_accum_90__60_,
  prod_accum_90__59_,prod_accum_90__58_,prod_accum_90__57_,prod_accum_90__56_,
  prod_accum_90__55_,prod_accum_90__54_,prod_accum_90__53_,prod_accum_90__52_,prod_accum_90__51_,
  prod_accum_90__50_,prod_accum_90__49_,prod_accum_90__48_,prod_accum_90__47_,
  prod_accum_90__46_,prod_accum_90__45_,prod_accum_90__44_,prod_accum_90__43_,
  prod_accum_90__42_,prod_accum_90__41_,prod_accum_90__40_,prod_accum_90__39_,
  prod_accum_90__38_,prod_accum_90__37_,prod_accum_90__36_,prod_accum_90__35_,
  prod_accum_90__34_,prod_accum_90__33_,prod_accum_90__32_,prod_accum_90__31_,prod_accum_90__30_,
  prod_accum_90__29_,prod_accum_90__28_,prod_accum_90__27_,prod_accum_90__26_,
  prod_accum_90__25_,prod_accum_90__24_,prod_accum_90__23_,prod_accum_90__22_,
  prod_accum_90__21_,prod_accum_90__20_,prod_accum_90__19_,prod_accum_90__18_,
  prod_accum_90__17_,prod_accum_90__16_,prod_accum_90__15_,prod_accum_90__14_,
  prod_accum_90__13_,prod_accum_90__12_,prod_accum_90__11_,prod_accum_90__10_,prod_accum_90__9_,
  prod_accum_90__8_,prod_accum_90__7_,prod_accum_90__6_,prod_accum_90__5_,
  prod_accum_90__4_,prod_accum_90__3_,prod_accum_90__2_,prod_accum_90__1_,prod_accum_90__0_,
  prod_accum_89__90_,prod_accum_89__89_,prod_accum_89__88_,prod_accum_89__87_,
  prod_accum_89__86_,prod_accum_89__85_,prod_accum_89__84_,prod_accum_89__83_,
  prod_accum_89__82_,prod_accum_89__81_,prod_accum_89__80_,prod_accum_89__79_,
  prod_accum_89__78_,prod_accum_89__77_,prod_accum_89__76_,prod_accum_89__75_,
  prod_accum_89__74_,prod_accum_89__73_,prod_accum_89__72_,prod_accum_89__71_,prod_accum_89__70_,
  prod_accum_89__69_,prod_accum_89__68_,prod_accum_89__67_,prod_accum_89__66_,
  prod_accum_89__65_,prod_accum_89__64_,prod_accum_89__63_,prod_accum_89__62_,
  prod_accum_89__61_,prod_accum_89__60_,prod_accum_89__59_,prod_accum_89__58_,
  prod_accum_89__57_,prod_accum_89__56_,prod_accum_89__55_,prod_accum_89__54_,prod_accum_89__53_,
  prod_accum_89__52_,prod_accum_89__51_,prod_accum_89__50_,prod_accum_89__49_,
  prod_accum_89__48_,prod_accum_89__47_,prod_accum_89__46_,prod_accum_89__45_,
  prod_accum_89__44_,prod_accum_89__43_,prod_accum_89__42_,prod_accum_89__41_,
  prod_accum_89__40_,prod_accum_89__39_,prod_accum_89__38_,prod_accum_89__37_,
  prod_accum_89__36_,prod_accum_89__35_,prod_accum_89__34_,prod_accum_89__33_,prod_accum_89__32_,
  prod_accum_89__31_,prod_accum_89__30_,prod_accum_89__29_,prod_accum_89__28_,
  prod_accum_89__27_,prod_accum_89__26_,prod_accum_89__25_,prod_accum_89__24_,
  prod_accum_89__23_,prod_accum_89__22_,prod_accum_89__21_,prod_accum_89__20_,
  prod_accum_89__19_,prod_accum_89__18_,prod_accum_89__17_,prod_accum_89__16_,
  prod_accum_89__15_,prod_accum_89__14_,prod_accum_89__13_,prod_accum_89__12_,prod_accum_89__11_,
  prod_accum_89__10_,prod_accum_89__9_,prod_accum_89__8_,prod_accum_89__7_,
  prod_accum_89__6_,prod_accum_89__5_,prod_accum_89__4_,prod_accum_89__3_,
  prod_accum_89__2_,prod_accum_89__1_,prod_accum_89__0_,prod_accum_88__89_,prod_accum_88__88_,
  prod_accum_88__87_,prod_accum_88__86_,prod_accum_88__85_,prod_accum_88__84_,
  prod_accum_88__83_,prod_accum_88__82_,prod_accum_88__81_,prod_accum_88__80_,
  prod_accum_88__79_,prod_accum_88__78_,prod_accum_88__77_,prod_accum_88__76_,
  prod_accum_88__75_,prod_accum_88__74_,prod_accum_88__73_,prod_accum_88__72_,prod_accum_88__71_,
  prod_accum_88__70_,prod_accum_88__69_,prod_accum_88__68_,prod_accum_88__67_,
  prod_accum_88__66_,prod_accum_88__65_,prod_accum_88__64_,prod_accum_88__63_,
  prod_accum_88__62_,prod_accum_88__61_,prod_accum_88__60_,prod_accum_88__59_,
  prod_accum_88__58_,prod_accum_88__57_,prod_accum_88__56_,prod_accum_88__55_,
  prod_accum_88__54_,prod_accum_88__53_,prod_accum_88__52_,prod_accum_88__51_,prod_accum_88__50_,
  prod_accum_88__49_,prod_accum_88__48_,prod_accum_88__47_,prod_accum_88__46_,
  prod_accum_88__45_,prod_accum_88__44_,prod_accum_88__43_,prod_accum_88__42_,
  prod_accum_88__41_,prod_accum_88__40_,prod_accum_88__39_,prod_accum_88__38_,
  prod_accum_88__37_,prod_accum_88__36_,prod_accum_88__35_,prod_accum_88__34_,prod_accum_88__33_,
  prod_accum_88__32_,prod_accum_88__31_,prod_accum_88__30_,prod_accum_88__29_,
  prod_accum_88__28_,prod_accum_88__27_,prod_accum_88__26_,prod_accum_88__25_,
  prod_accum_88__24_,prod_accum_88__23_,prod_accum_88__22_,prod_accum_88__21_,
  prod_accum_88__20_,prod_accum_88__19_,prod_accum_88__18_,prod_accum_88__17_,
  prod_accum_88__16_,prod_accum_88__15_,prod_accum_88__14_,prod_accum_88__13_,prod_accum_88__12_,
  prod_accum_88__11_,prod_accum_88__10_,prod_accum_88__9_,prod_accum_88__8_,
  prod_accum_88__7_,prod_accum_88__6_,prod_accum_88__5_,prod_accum_88__4_,
  prod_accum_88__3_,prod_accum_88__2_,prod_accum_88__1_,prod_accum_88__0_,prod_accum_87__88_,
  prod_accum_87__87_,prod_accum_87__86_,prod_accum_87__85_,prod_accum_87__84_,
  prod_accum_87__83_,prod_accum_87__82_,prod_accum_87__81_,prod_accum_87__80_,
  prod_accum_87__79_,prod_accum_87__78_,prod_accum_87__77_,prod_accum_87__76_,
  prod_accum_87__75_,prod_accum_87__74_,prod_accum_87__73_,prod_accum_87__72_,prod_accum_87__71_,
  prod_accum_87__70_,prod_accum_87__69_,prod_accum_87__68_,prod_accum_87__67_,
  prod_accum_87__66_,prod_accum_87__65_,prod_accum_87__64_,prod_accum_87__63_,
  prod_accum_87__62_,prod_accum_87__61_,prod_accum_87__60_,prod_accum_87__59_,
  prod_accum_87__58_,prod_accum_87__57_,prod_accum_87__56_,prod_accum_87__55_,
  prod_accum_87__54_,prod_accum_87__53_,prod_accum_87__52_,prod_accum_87__51_,prod_accum_87__50_,
  prod_accum_87__49_,prod_accum_87__48_,prod_accum_87__47_,prod_accum_87__46_,
  prod_accum_87__45_,prod_accum_87__44_,prod_accum_87__43_,prod_accum_87__42_,
  prod_accum_87__41_,prod_accum_87__40_,prod_accum_87__39_,prod_accum_87__38_,
  prod_accum_87__37_,prod_accum_87__36_,prod_accum_87__35_,prod_accum_87__34_,
  prod_accum_87__33_,prod_accum_87__32_,prod_accum_87__31_,prod_accum_87__30_,prod_accum_87__29_,
  prod_accum_87__28_,prod_accum_87__27_,prod_accum_87__26_,prod_accum_87__25_,
  prod_accum_87__24_,prod_accum_87__23_,prod_accum_87__22_,prod_accum_87__21_,
  prod_accum_87__20_,prod_accum_87__19_,prod_accum_87__18_,prod_accum_87__17_,
  prod_accum_87__16_,prod_accum_87__15_,prod_accum_87__14_,prod_accum_87__13_,prod_accum_87__12_,
  prod_accum_87__11_,prod_accum_87__10_,prod_accum_87__9_,prod_accum_87__8_,
  prod_accum_87__7_,prod_accum_87__6_,prod_accum_87__5_,prod_accum_87__4_,
  prod_accum_87__3_,prod_accum_87__2_,prod_accum_87__1_,prod_accum_87__0_,s_r_94__127_,
  s_r_94__126_,s_r_94__125_,s_r_94__124_,s_r_94__123_,s_r_94__122_,s_r_94__121_,
  s_r_94__120_,s_r_94__119_,s_r_94__118_,s_r_94__117_,s_r_94__116_,s_r_94__115_,s_r_94__114_,
  s_r_94__113_,s_r_94__112_,s_r_94__111_,s_r_94__110_,s_r_94__109_,s_r_94__108_,
  s_r_94__107_,s_r_94__106_,s_r_94__105_,s_r_94__104_,s_r_94__103_,s_r_94__102_,
  s_r_94__101_,s_r_94__100_,s_r_94__99_,s_r_94__98_,s_r_94__97_,s_r_94__96_,
  s_r_94__95_,s_r_94__94_,s_r_94__93_,s_r_94__92_,s_r_94__91_,s_r_94__90_,s_r_94__89_,
  s_r_94__88_,s_r_94__87_,s_r_94__86_,s_r_94__85_,s_r_94__84_,s_r_94__83_,s_r_94__82_,
  s_r_94__81_,s_r_94__80_,s_r_94__79_,s_r_94__78_,s_r_94__77_,s_r_94__76_,
  s_r_94__75_,s_r_94__74_,s_r_94__73_,s_r_94__72_,s_r_94__71_,s_r_94__70_,s_r_94__69_,
  s_r_94__68_,s_r_94__67_,s_r_94__66_,s_r_94__65_,s_r_94__64_,s_r_94__63_,s_r_94__62_,
  s_r_94__61_,s_r_94__60_,s_r_94__59_,s_r_94__58_,s_r_94__57_,s_r_94__56_,
  s_r_94__55_,s_r_94__54_,s_r_94__53_,s_r_94__52_,s_r_94__51_,s_r_94__50_,s_r_94__49_,
  s_r_94__48_,s_r_94__47_,s_r_94__46_,s_r_94__45_,s_r_94__44_,s_r_94__43_,s_r_94__42_,
  s_r_94__41_,s_r_94__40_,s_r_94__39_,s_r_94__38_,s_r_94__37_,s_r_94__36_,
  s_r_94__35_,s_r_94__34_,s_r_94__33_,s_r_94__32_,s_r_94__31_,s_r_94__30_,s_r_94__29_,
  s_r_94__28_,s_r_94__27_,s_r_94__26_,s_r_94__25_,s_r_94__24_,s_r_94__23_,s_r_94__22_,
  s_r_94__21_,s_r_94__20_,s_r_94__19_,s_r_94__18_,s_r_94__17_,s_r_94__16_,
  s_r_94__15_,s_r_94__14_,s_r_94__13_,s_r_94__12_,s_r_94__11_,s_r_94__10_,s_r_94__9_,
  s_r_94__8_,s_r_94__7_,s_r_94__6_,s_r_94__5_,s_r_94__4_,s_r_94__3_,s_r_94__2_,
  s_r_94__1_,s_r_94__0_,s_r_93__127_,s_r_93__126_,s_r_93__125_,s_r_93__124_,s_r_93__123_,
  s_r_93__122_,s_r_93__121_,s_r_93__120_,s_r_93__119_,s_r_93__118_,s_r_93__117_,
  s_r_93__116_,s_r_93__115_,s_r_93__114_,s_r_93__113_,s_r_93__112_,s_r_93__111_,
  s_r_93__110_,s_r_93__109_,s_r_93__108_,s_r_93__107_,s_r_93__106_,s_r_93__105_,
  s_r_93__104_,s_r_93__103_,s_r_93__102_,s_r_93__101_,s_r_93__100_,s_r_93__99_,s_r_93__98_,
  s_r_93__97_,s_r_93__96_,s_r_93__95_,s_r_93__94_,s_r_93__93_,s_r_93__92_,
  s_r_93__91_,s_r_93__90_,s_r_93__89_,s_r_93__88_,s_r_93__87_,s_r_93__86_,s_r_93__85_,
  s_r_93__84_,s_r_93__83_,s_r_93__82_,s_r_93__81_,s_r_93__80_,s_r_93__79_,s_r_93__78_,
  s_r_93__77_,s_r_93__76_,s_r_93__75_,s_r_93__74_,s_r_93__73_,s_r_93__72_,
  s_r_93__71_,s_r_93__70_,s_r_93__69_,s_r_93__68_,s_r_93__67_,s_r_93__66_,s_r_93__65_,
  s_r_93__64_,s_r_93__63_,s_r_93__62_,s_r_93__61_,s_r_93__60_,s_r_93__59_,s_r_93__58_,
  s_r_93__57_,s_r_93__56_,s_r_93__55_,s_r_93__54_,s_r_93__53_,s_r_93__52_,
  s_r_93__51_,s_r_93__50_,s_r_93__49_,s_r_93__48_,s_r_93__47_,s_r_93__46_,s_r_93__45_,
  s_r_93__44_,s_r_93__43_,s_r_93__42_,s_r_93__41_,s_r_93__40_,s_r_93__39_,s_r_93__38_,
  s_r_93__37_,s_r_93__36_,s_r_93__35_,s_r_93__34_,s_r_93__33_,s_r_93__32_,
  s_r_93__31_,s_r_93__30_,s_r_93__29_,s_r_93__28_,s_r_93__27_,s_r_93__26_,s_r_93__25_,
  s_r_93__24_,s_r_93__23_,s_r_93__22_,s_r_93__21_,s_r_93__20_,s_r_93__19_,s_r_93__18_,
  s_r_93__17_,s_r_93__16_,s_r_93__15_,s_r_93__14_,s_r_93__13_,s_r_93__12_,
  s_r_93__11_,s_r_93__10_,s_r_93__9_,s_r_93__8_,s_r_93__7_,s_r_93__6_,s_r_93__5_,
  s_r_93__4_,s_r_93__3_,s_r_93__2_,s_r_93__1_,s_r_93__0_,s_r_92__127_,s_r_92__126_,
  s_r_92__125_,s_r_92__124_,s_r_92__123_,s_r_92__122_,s_r_92__121_,s_r_92__120_,
  s_r_92__119_,s_r_92__118_,s_r_92__117_,s_r_92__116_,s_r_92__115_,s_r_92__114_,
  s_r_92__113_,s_r_92__112_,s_r_92__111_,s_r_92__110_,s_r_92__109_,s_r_92__108_,s_r_92__107_,
  s_r_92__106_,s_r_92__105_,s_r_92__104_,s_r_92__103_,s_r_92__102_,s_r_92__101_,
  s_r_92__100_,s_r_92__99_,s_r_92__98_,s_r_92__97_,s_r_92__96_,s_r_92__95_,
  s_r_92__94_,s_r_92__93_,s_r_92__92_,s_r_92__91_,s_r_92__90_,s_r_92__89_,s_r_92__88_,
  s_r_92__87_,s_r_92__86_,s_r_92__85_,s_r_92__84_,s_r_92__83_,s_r_92__82_,s_r_92__81_,
  s_r_92__80_,s_r_92__79_,s_r_92__78_,s_r_92__77_,s_r_92__76_,s_r_92__75_,
  s_r_92__74_,s_r_92__73_,s_r_92__72_,s_r_92__71_,s_r_92__70_,s_r_92__69_,s_r_92__68_,
  s_r_92__67_,s_r_92__66_,s_r_92__65_,s_r_92__64_,s_r_92__63_,s_r_92__62_,s_r_92__61_,
  s_r_92__60_,s_r_92__59_,s_r_92__58_,s_r_92__57_,s_r_92__56_,s_r_92__55_,
  s_r_92__54_,s_r_92__53_,s_r_92__52_,s_r_92__51_,s_r_92__50_,s_r_92__49_,s_r_92__48_,
  s_r_92__47_,s_r_92__46_,s_r_92__45_,s_r_92__44_,s_r_92__43_,s_r_92__42_,s_r_92__41_,
  s_r_92__40_,s_r_92__39_,s_r_92__38_,s_r_92__37_,s_r_92__36_,s_r_92__35_,
  s_r_92__34_,s_r_92__33_,s_r_92__32_,s_r_92__31_,s_r_92__30_,s_r_92__29_,s_r_92__28_,
  s_r_92__27_,s_r_92__26_,s_r_92__25_,s_r_92__24_,s_r_92__23_,s_r_92__22_,s_r_92__21_,
  s_r_92__20_,s_r_92__19_,s_r_92__18_,s_r_92__17_,s_r_92__16_,s_r_92__15_,
  s_r_92__14_,s_r_92__13_,s_r_92__12_,s_r_92__11_,s_r_92__10_,s_r_92__9_,s_r_92__8_,
  s_r_92__7_,s_r_92__6_,s_r_92__5_,s_r_92__4_,s_r_92__3_,s_r_92__2_,s_r_92__1_,s_r_92__0_,
  s_r_91__127_,s_r_91__126_,s_r_91__125_,s_r_91__124_,s_r_91__123_,s_r_91__122_,
  s_r_91__121_,s_r_91__120_,s_r_91__119_,s_r_91__118_,s_r_91__117_,s_r_91__116_,
  s_r_91__115_,s_r_91__114_,s_r_91__113_,s_r_91__112_,s_r_91__111_,s_r_91__110_,
  s_r_91__109_,s_r_91__108_,s_r_91__107_,s_r_91__106_,s_r_91__105_,s_r_91__104_,
  s_r_91__103_,s_r_91__102_,s_r_91__101_,s_r_91__100_,s_r_91__99_,s_r_91__98_,s_r_91__97_,
  s_r_91__96_,s_r_91__95_,s_r_91__94_,s_r_91__93_,s_r_91__92_,s_r_91__91_,
  s_r_91__90_,s_r_91__89_,s_r_91__88_,s_r_91__87_,s_r_91__86_,s_r_91__85_,s_r_91__84_,
  s_r_91__83_,s_r_91__82_,s_r_91__81_,s_r_91__80_,s_r_91__79_,s_r_91__78_,s_r_91__77_,
  s_r_91__76_,s_r_91__75_,s_r_91__74_,s_r_91__73_,s_r_91__72_,s_r_91__71_,
  s_r_91__70_,s_r_91__69_,s_r_91__68_,s_r_91__67_,s_r_91__66_,s_r_91__65_,s_r_91__64_,
  s_r_91__63_,s_r_91__62_,s_r_91__61_,s_r_91__60_,s_r_91__59_,s_r_91__58_,s_r_91__57_,
  s_r_91__56_,s_r_91__55_,s_r_91__54_,s_r_91__53_,s_r_91__52_,s_r_91__51_,
  s_r_91__50_,s_r_91__49_,s_r_91__48_,s_r_91__47_,s_r_91__46_,s_r_91__45_,s_r_91__44_,
  s_r_91__43_,s_r_91__42_,s_r_91__41_,s_r_91__40_,s_r_91__39_,s_r_91__38_,s_r_91__37_,
  s_r_91__36_,s_r_91__35_,s_r_91__34_,s_r_91__33_,s_r_91__32_,s_r_91__31_,
  s_r_91__30_,s_r_91__29_,s_r_91__28_,s_r_91__27_,s_r_91__26_,s_r_91__25_,s_r_91__24_,
  s_r_91__23_,s_r_91__22_,s_r_91__21_,s_r_91__20_,s_r_91__19_,s_r_91__18_,s_r_91__17_,
  s_r_91__16_,s_r_91__15_,s_r_91__14_,s_r_91__13_,s_r_91__12_,s_r_91__11_,
  s_r_91__10_,s_r_91__9_,s_r_91__8_,s_r_91__7_,s_r_91__6_,s_r_91__5_,s_r_91__4_,
  s_r_91__3_,s_r_91__2_,s_r_91__1_,s_r_91__0_,prod_accum_94__95_,prod_accum_94__94_,
  prod_accum_94__93_,prod_accum_94__92_,prod_accum_94__91_,prod_accum_94__90_,
  prod_accum_94__89_,prod_accum_94__88_,prod_accum_94__87_,prod_accum_94__86_,
  prod_accum_94__85_,prod_accum_94__84_,prod_accum_94__83_,prod_accum_94__82_,prod_accum_94__81_,
  prod_accum_94__80_,prod_accum_94__79_,prod_accum_94__78_,prod_accum_94__77_,
  prod_accum_94__76_,prod_accum_94__75_,prod_accum_94__74_,prod_accum_94__73_,
  prod_accum_94__72_,prod_accum_94__71_,prod_accum_94__70_,prod_accum_94__69_,
  prod_accum_94__68_,prod_accum_94__67_,prod_accum_94__66_,prod_accum_94__65_,
  prod_accum_94__64_,prod_accum_94__63_,prod_accum_94__62_,prod_accum_94__61_,prod_accum_94__60_,
  prod_accum_94__59_,prod_accum_94__58_,prod_accum_94__57_,prod_accum_94__56_,
  prod_accum_94__55_,prod_accum_94__54_,prod_accum_94__53_,prod_accum_94__52_,
  prod_accum_94__51_,prod_accum_94__50_,prod_accum_94__49_,prod_accum_94__48_,
  prod_accum_94__47_,prod_accum_94__46_,prod_accum_94__45_,prod_accum_94__44_,
  prod_accum_94__43_,prod_accum_94__42_,prod_accum_94__41_,prod_accum_94__40_,prod_accum_94__39_,
  prod_accum_94__38_,prod_accum_94__37_,prod_accum_94__36_,prod_accum_94__35_,
  prod_accum_94__34_,prod_accum_94__33_,prod_accum_94__32_,prod_accum_94__31_,
  prod_accum_94__30_,prod_accum_94__29_,prod_accum_94__28_,prod_accum_94__27_,
  prod_accum_94__26_,prod_accum_94__25_,prod_accum_94__24_,prod_accum_94__23_,prod_accum_94__22_,
  prod_accum_94__21_,prod_accum_94__20_,prod_accum_94__19_,prod_accum_94__18_,
  prod_accum_94__17_,prod_accum_94__16_,prod_accum_94__15_,prod_accum_94__14_,
  prod_accum_94__13_,prod_accum_94__12_,prod_accum_94__11_,prod_accum_94__10_,
  prod_accum_94__9_,prod_accum_94__8_,prod_accum_94__7_,prod_accum_94__6_,prod_accum_94__5_,
  prod_accum_94__4_,prod_accum_94__3_,prod_accum_94__2_,prod_accum_94__1_,
  prod_accum_94__0_,prod_accum_93__94_,prod_accum_93__93_,prod_accum_93__92_,
  prod_accum_93__91_,prod_accum_93__90_,prod_accum_93__89_,prod_accum_93__88_,prod_accum_93__87_,
  prod_accum_93__86_,prod_accum_93__85_,prod_accum_93__84_,prod_accum_93__83_,
  prod_accum_93__82_,prod_accum_93__81_,prod_accum_93__80_,prod_accum_93__79_,
  prod_accum_93__78_,prod_accum_93__77_,prod_accum_93__76_,prod_accum_93__75_,
  prod_accum_93__74_,prod_accum_93__73_,prod_accum_93__72_,prod_accum_93__71_,
  prod_accum_93__70_,prod_accum_93__69_,prod_accum_93__68_,prod_accum_93__67_,prod_accum_93__66_,
  prod_accum_93__65_,prod_accum_93__64_,prod_accum_93__63_,prod_accum_93__62_,
  prod_accum_93__61_,prod_accum_93__60_,prod_accum_93__59_,prod_accum_93__58_,
  prod_accum_93__57_,prod_accum_93__56_,prod_accum_93__55_,prod_accum_93__54_,
  prod_accum_93__53_,prod_accum_93__52_,prod_accum_93__51_,prod_accum_93__50_,
  prod_accum_93__49_,prod_accum_93__48_,prod_accum_93__47_,prod_accum_93__46_,prod_accum_93__45_,
  prod_accum_93__44_,prod_accum_93__43_,prod_accum_93__42_,prod_accum_93__41_,
  prod_accum_93__40_,prod_accum_93__39_,prod_accum_93__38_,prod_accum_93__37_,
  prod_accum_93__36_,prod_accum_93__35_,prod_accum_93__34_,prod_accum_93__33_,
  prod_accum_93__32_,prod_accum_93__31_,prod_accum_93__30_,prod_accum_93__29_,
  prod_accum_93__28_,prod_accum_93__27_,prod_accum_93__26_,prod_accum_93__25_,prod_accum_93__24_,
  prod_accum_93__23_,prod_accum_93__22_,prod_accum_93__21_,prod_accum_93__20_,
  prod_accum_93__19_,prod_accum_93__18_,prod_accum_93__17_,prod_accum_93__16_,
  prod_accum_93__15_,prod_accum_93__14_,prod_accum_93__13_,prod_accum_93__12_,
  prod_accum_93__11_,prod_accum_93__10_,prod_accum_93__9_,prod_accum_93__8_,prod_accum_93__7_,
  prod_accum_93__6_,prod_accum_93__5_,prod_accum_93__4_,prod_accum_93__3_,
  prod_accum_93__2_,prod_accum_93__1_,prod_accum_93__0_,prod_accum_92__93_,
  prod_accum_92__92_,prod_accum_92__91_,prod_accum_92__90_,prod_accum_92__89_,prod_accum_92__88_,
  prod_accum_92__87_,prod_accum_92__86_,prod_accum_92__85_,prod_accum_92__84_,
  prod_accum_92__83_,prod_accum_92__82_,prod_accum_92__81_,prod_accum_92__80_,
  prod_accum_92__79_,prod_accum_92__78_,prod_accum_92__77_,prod_accum_92__76_,
  prod_accum_92__75_,prod_accum_92__74_,prod_accum_92__73_,prod_accum_92__72_,prod_accum_92__71_,
  prod_accum_92__70_,prod_accum_92__69_,prod_accum_92__68_,prod_accum_92__67_,
  prod_accum_92__66_,prod_accum_92__65_,prod_accum_92__64_,prod_accum_92__63_,
  prod_accum_92__62_,prod_accum_92__61_,prod_accum_92__60_,prod_accum_92__59_,
  prod_accum_92__58_,prod_accum_92__57_,prod_accum_92__56_,prod_accum_92__55_,
  prod_accum_92__54_,prod_accum_92__53_,prod_accum_92__52_,prod_accum_92__51_,prod_accum_92__50_,
  prod_accum_92__49_,prod_accum_92__48_,prod_accum_92__47_,prod_accum_92__46_,
  prod_accum_92__45_,prod_accum_92__44_,prod_accum_92__43_,prod_accum_92__42_,
  prod_accum_92__41_,prod_accum_92__40_,prod_accum_92__39_,prod_accum_92__38_,
  prod_accum_92__37_,prod_accum_92__36_,prod_accum_92__35_,prod_accum_92__34_,
  prod_accum_92__33_,prod_accum_92__32_,prod_accum_92__31_,prod_accum_92__30_,prod_accum_92__29_,
  prod_accum_92__28_,prod_accum_92__27_,prod_accum_92__26_,prod_accum_92__25_,
  prod_accum_92__24_,prod_accum_92__23_,prod_accum_92__22_,prod_accum_92__21_,
  prod_accum_92__20_,prod_accum_92__19_,prod_accum_92__18_,prod_accum_92__17_,
  prod_accum_92__16_,prod_accum_92__15_,prod_accum_92__14_,prod_accum_92__13_,
  prod_accum_92__12_,prod_accum_92__11_,prod_accum_92__10_,prod_accum_92__9_,prod_accum_92__8_,
  prod_accum_92__7_,prod_accum_92__6_,prod_accum_92__5_,prod_accum_92__4_,
  prod_accum_92__3_,prod_accum_92__2_,prod_accum_92__1_,prod_accum_92__0_,prod_accum_91__92_,
  prod_accum_91__91_,prod_accum_91__90_,prod_accum_91__89_,prod_accum_91__88_,
  prod_accum_91__87_,prod_accum_91__86_,prod_accum_91__85_,prod_accum_91__84_,
  prod_accum_91__83_,prod_accum_91__82_,prod_accum_91__81_,prod_accum_91__80_,
  prod_accum_91__79_,prod_accum_91__78_,prod_accum_91__77_,prod_accum_91__76_,
  prod_accum_91__75_,prod_accum_91__74_,prod_accum_91__73_,prod_accum_91__72_,prod_accum_91__71_,
  prod_accum_91__70_,prod_accum_91__69_,prod_accum_91__68_,prod_accum_91__67_,
  prod_accum_91__66_,prod_accum_91__65_,prod_accum_91__64_,prod_accum_91__63_,
  prod_accum_91__62_,prod_accum_91__61_,prod_accum_91__60_,prod_accum_91__59_,
  prod_accum_91__58_,prod_accum_91__57_,prod_accum_91__56_,prod_accum_91__55_,prod_accum_91__54_,
  prod_accum_91__53_,prod_accum_91__52_,prod_accum_91__51_,prod_accum_91__50_,
  prod_accum_91__49_,prod_accum_91__48_,prod_accum_91__47_,prod_accum_91__46_,
  prod_accum_91__45_,prod_accum_91__44_,prod_accum_91__43_,prod_accum_91__42_,
  prod_accum_91__41_,prod_accum_91__40_,prod_accum_91__39_,prod_accum_91__38_,
  prod_accum_91__37_,prod_accum_91__36_,prod_accum_91__35_,prod_accum_91__34_,prod_accum_91__33_,
  prod_accum_91__32_,prod_accum_91__31_,prod_accum_91__30_,prod_accum_91__29_,
  prod_accum_91__28_,prod_accum_91__27_,prod_accum_91__26_,prod_accum_91__25_,
  prod_accum_91__24_,prod_accum_91__23_,prod_accum_91__22_,prod_accum_91__21_,
  prod_accum_91__20_,prod_accum_91__19_,prod_accum_91__18_,prod_accum_91__17_,
  prod_accum_91__16_,prod_accum_91__15_,prod_accum_91__14_,prod_accum_91__13_,prod_accum_91__12_,
  prod_accum_91__11_,prod_accum_91__10_,prod_accum_91__9_,prod_accum_91__8_,
  prod_accum_91__7_,prod_accum_91__6_,prod_accum_91__5_,prod_accum_91__4_,
  prod_accum_91__3_,prod_accum_91__2_,prod_accum_91__1_,prod_accum_91__0_,s_r_98__127_,
  s_r_98__126_,s_r_98__125_,s_r_98__124_,s_r_98__123_,s_r_98__122_,s_r_98__121_,s_r_98__120_,
  s_r_98__119_,s_r_98__118_,s_r_98__117_,s_r_98__116_,s_r_98__115_,s_r_98__114_,
  s_r_98__113_,s_r_98__112_,s_r_98__111_,s_r_98__110_,s_r_98__109_,s_r_98__108_,
  s_r_98__107_,s_r_98__106_,s_r_98__105_,s_r_98__104_,s_r_98__103_,s_r_98__102_,
  s_r_98__101_,s_r_98__100_,s_r_98__99_,s_r_98__98_,s_r_98__97_,s_r_98__96_,s_r_98__95_,
  s_r_98__94_,s_r_98__93_,s_r_98__92_,s_r_98__91_,s_r_98__90_,s_r_98__89_,
  s_r_98__88_,s_r_98__87_,s_r_98__86_,s_r_98__85_,s_r_98__84_,s_r_98__83_,s_r_98__82_,
  s_r_98__81_,s_r_98__80_,s_r_98__79_,s_r_98__78_,s_r_98__77_,s_r_98__76_,s_r_98__75_,
  s_r_98__74_,s_r_98__73_,s_r_98__72_,s_r_98__71_,s_r_98__70_,s_r_98__69_,
  s_r_98__68_,s_r_98__67_,s_r_98__66_,s_r_98__65_,s_r_98__64_,s_r_98__63_,s_r_98__62_,
  s_r_98__61_,s_r_98__60_,s_r_98__59_,s_r_98__58_,s_r_98__57_,s_r_98__56_,s_r_98__55_,
  s_r_98__54_,s_r_98__53_,s_r_98__52_,s_r_98__51_,s_r_98__50_,s_r_98__49_,
  s_r_98__48_,s_r_98__47_,s_r_98__46_,s_r_98__45_,s_r_98__44_,s_r_98__43_,s_r_98__42_,
  s_r_98__41_,s_r_98__40_,s_r_98__39_,s_r_98__38_,s_r_98__37_,s_r_98__36_,s_r_98__35_,
  s_r_98__34_,s_r_98__33_,s_r_98__32_,s_r_98__31_,s_r_98__30_,s_r_98__29_,
  s_r_98__28_,s_r_98__27_,s_r_98__26_,s_r_98__25_,s_r_98__24_,s_r_98__23_,s_r_98__22_,
  s_r_98__21_,s_r_98__20_,s_r_98__19_,s_r_98__18_,s_r_98__17_,s_r_98__16_,s_r_98__15_,
  s_r_98__14_,s_r_98__13_,s_r_98__12_,s_r_98__11_,s_r_98__10_,s_r_98__9_,
  s_r_98__8_,s_r_98__7_,s_r_98__6_,s_r_98__5_,s_r_98__4_,s_r_98__3_,s_r_98__2_,s_r_98__1_,
  s_r_98__0_,s_r_97__127_,s_r_97__126_,s_r_97__125_,s_r_97__124_,s_r_97__123_,
  s_r_97__122_,s_r_97__121_,s_r_97__120_,s_r_97__119_,s_r_97__118_,s_r_97__117_,
  s_r_97__116_,s_r_97__115_,s_r_97__114_,s_r_97__113_,s_r_97__112_,s_r_97__111_,
  s_r_97__110_,s_r_97__109_,s_r_97__108_,s_r_97__107_,s_r_97__106_,s_r_97__105_,
  s_r_97__104_,s_r_97__103_,s_r_97__102_,s_r_97__101_,s_r_97__100_,s_r_97__99_,s_r_97__98_,
  s_r_97__97_,s_r_97__96_,s_r_97__95_,s_r_97__94_,s_r_97__93_,s_r_97__92_,
  s_r_97__91_,s_r_97__90_,s_r_97__89_,s_r_97__88_,s_r_97__87_,s_r_97__86_,s_r_97__85_,
  s_r_97__84_,s_r_97__83_,s_r_97__82_,s_r_97__81_,s_r_97__80_,s_r_97__79_,s_r_97__78_,
  s_r_97__77_,s_r_97__76_,s_r_97__75_,s_r_97__74_,s_r_97__73_,s_r_97__72_,
  s_r_97__71_,s_r_97__70_,s_r_97__69_,s_r_97__68_,s_r_97__67_,s_r_97__66_,s_r_97__65_,
  s_r_97__64_,s_r_97__63_,s_r_97__62_,s_r_97__61_,s_r_97__60_,s_r_97__59_,s_r_97__58_,
  s_r_97__57_,s_r_97__56_,s_r_97__55_,s_r_97__54_,s_r_97__53_,s_r_97__52_,
  s_r_97__51_,s_r_97__50_,s_r_97__49_,s_r_97__48_,s_r_97__47_,s_r_97__46_,s_r_97__45_,
  s_r_97__44_,s_r_97__43_,s_r_97__42_,s_r_97__41_,s_r_97__40_,s_r_97__39_,s_r_97__38_,
  s_r_97__37_,s_r_97__36_,s_r_97__35_,s_r_97__34_,s_r_97__33_,s_r_97__32_,
  s_r_97__31_,s_r_97__30_,s_r_97__29_,s_r_97__28_,s_r_97__27_,s_r_97__26_,s_r_97__25_,
  s_r_97__24_,s_r_97__23_,s_r_97__22_,s_r_97__21_,s_r_97__20_,s_r_97__19_,s_r_97__18_,
  s_r_97__17_,s_r_97__16_,s_r_97__15_,s_r_97__14_,s_r_97__13_,s_r_97__12_,
  s_r_97__11_,s_r_97__10_,s_r_97__9_,s_r_97__8_,s_r_97__7_,s_r_97__6_,s_r_97__5_,s_r_97__4_,
  s_r_97__3_,s_r_97__2_,s_r_97__1_,s_r_97__0_,s_r_96__127_,s_r_96__126_,
  s_r_96__125_,s_r_96__124_,s_r_96__123_,s_r_96__122_,s_r_96__121_,s_r_96__120_,
  s_r_96__119_,s_r_96__118_,s_r_96__117_,s_r_96__116_,s_r_96__115_,s_r_96__114_,s_r_96__113_,
  s_r_96__112_,s_r_96__111_,s_r_96__110_,s_r_96__109_,s_r_96__108_,s_r_96__107_,
  s_r_96__106_,s_r_96__105_,s_r_96__104_,s_r_96__103_,s_r_96__102_,s_r_96__101_,
  s_r_96__100_,s_r_96__99_,s_r_96__98_,s_r_96__97_,s_r_96__96_,s_r_96__95_,s_r_96__94_,
  s_r_96__93_,s_r_96__92_,s_r_96__91_,s_r_96__90_,s_r_96__89_,s_r_96__88_,
  s_r_96__87_,s_r_96__86_,s_r_96__85_,s_r_96__84_,s_r_96__83_,s_r_96__82_,s_r_96__81_,
  s_r_96__80_,s_r_96__79_,s_r_96__78_,s_r_96__77_,s_r_96__76_,s_r_96__75_,s_r_96__74_,
  s_r_96__73_,s_r_96__72_,s_r_96__71_,s_r_96__70_,s_r_96__69_,s_r_96__68_,
  s_r_96__67_,s_r_96__66_,s_r_96__65_,s_r_96__64_,s_r_96__63_,s_r_96__62_,s_r_96__61_,
  s_r_96__60_,s_r_96__59_,s_r_96__58_,s_r_96__57_,s_r_96__56_,s_r_96__55_,s_r_96__54_,
  s_r_96__53_,s_r_96__52_,s_r_96__51_,s_r_96__50_,s_r_96__49_,s_r_96__48_,
  s_r_96__47_,s_r_96__46_,s_r_96__45_,s_r_96__44_,s_r_96__43_,s_r_96__42_,s_r_96__41_,
  s_r_96__40_,s_r_96__39_,s_r_96__38_,s_r_96__37_,s_r_96__36_,s_r_96__35_,s_r_96__34_,
  s_r_96__33_,s_r_96__32_,s_r_96__31_,s_r_96__30_,s_r_96__29_,s_r_96__28_,
  s_r_96__27_,s_r_96__26_,s_r_96__25_,s_r_96__24_,s_r_96__23_,s_r_96__22_,s_r_96__21_,
  s_r_96__20_,s_r_96__19_,s_r_96__18_,s_r_96__17_,s_r_96__16_,s_r_96__15_,s_r_96__14_,
  s_r_96__13_,s_r_96__12_,s_r_96__11_,s_r_96__10_,s_r_96__9_,s_r_96__8_,
  s_r_96__7_,s_r_96__6_,s_r_96__5_,s_r_96__4_,s_r_96__3_,s_r_96__2_,s_r_96__1_,s_r_96__0_,
  s_r_95__127_,s_r_95__126_,s_r_95__125_,s_r_95__124_,s_r_95__123_,s_r_95__122_,
  s_r_95__121_,s_r_95__120_,s_r_95__119_,s_r_95__118_,s_r_95__117_,s_r_95__116_,
  s_r_95__115_,s_r_95__114_,s_r_95__113_,s_r_95__112_,s_r_95__111_,s_r_95__110_,
  s_r_95__109_,s_r_95__108_,s_r_95__107_,s_r_95__106_,s_r_95__105_,s_r_95__104_,
  s_r_95__103_,s_r_95__102_,s_r_95__101_,s_r_95__100_,s_r_95__99_,s_r_95__98_,s_r_95__97_,
  s_r_95__96_,s_r_95__95_,s_r_95__94_,s_r_95__93_,s_r_95__92_,s_r_95__91_,
  s_r_95__90_,s_r_95__89_,s_r_95__88_,s_r_95__87_,s_r_95__86_,s_r_95__85_,s_r_95__84_,
  s_r_95__83_,s_r_95__82_,s_r_95__81_,s_r_95__80_,s_r_95__79_,s_r_95__78_,s_r_95__77_,
  s_r_95__76_,s_r_95__75_,s_r_95__74_,s_r_95__73_,s_r_95__72_,s_r_95__71_,
  s_r_95__70_,s_r_95__69_,s_r_95__68_,s_r_95__67_,s_r_95__66_,s_r_95__65_,s_r_95__64_,
  s_r_95__63_,s_r_95__62_,s_r_95__61_,s_r_95__60_,s_r_95__59_,s_r_95__58_,s_r_95__57_,
  s_r_95__56_,s_r_95__55_,s_r_95__54_,s_r_95__53_,s_r_95__52_,s_r_95__51_,
  s_r_95__50_,s_r_95__49_,s_r_95__48_,s_r_95__47_,s_r_95__46_,s_r_95__45_,s_r_95__44_,
  s_r_95__43_,s_r_95__42_,s_r_95__41_,s_r_95__40_,s_r_95__39_,s_r_95__38_,s_r_95__37_,
  s_r_95__36_,s_r_95__35_,s_r_95__34_,s_r_95__33_,s_r_95__32_,s_r_95__31_,
  s_r_95__30_,s_r_95__29_,s_r_95__28_,s_r_95__27_,s_r_95__26_,s_r_95__25_,s_r_95__24_,
  s_r_95__23_,s_r_95__22_,s_r_95__21_,s_r_95__20_,s_r_95__19_,s_r_95__18_,s_r_95__17_,
  s_r_95__16_,s_r_95__15_,s_r_95__14_,s_r_95__13_,s_r_95__12_,s_r_95__11_,
  s_r_95__10_,s_r_95__9_,s_r_95__8_,s_r_95__7_,s_r_95__6_,s_r_95__5_,s_r_95__4_,s_r_95__3_,
  s_r_95__2_,s_r_95__1_,s_r_95__0_,prod_accum_98__99_,prod_accum_98__98_,
  prod_accum_98__97_,prod_accum_98__96_,prod_accum_98__95_,prod_accum_98__94_,
  prod_accum_98__93_,prod_accum_98__92_,prod_accum_98__91_,prod_accum_98__90_,
  prod_accum_98__89_,prod_accum_98__88_,prod_accum_98__87_,prod_accum_98__86_,prod_accum_98__85_,
  prod_accum_98__84_,prod_accum_98__83_,prod_accum_98__82_,prod_accum_98__81_,
  prod_accum_98__80_,prod_accum_98__79_,prod_accum_98__78_,prod_accum_98__77_,
  prod_accum_98__76_,prod_accum_98__75_,prod_accum_98__74_,prod_accum_98__73_,
  prod_accum_98__72_,prod_accum_98__71_,prod_accum_98__70_,prod_accum_98__69_,prod_accum_98__68_,
  prod_accum_98__67_,prod_accum_98__66_,prod_accum_98__65_,prod_accum_98__64_,
  prod_accum_98__63_,prod_accum_98__62_,prod_accum_98__61_,prod_accum_98__60_,
  prod_accum_98__59_,prod_accum_98__58_,prod_accum_98__57_,prod_accum_98__56_,
  prod_accum_98__55_,prod_accum_98__54_,prod_accum_98__53_,prod_accum_98__52_,
  prod_accum_98__51_,prod_accum_98__50_,prod_accum_98__49_,prod_accum_98__48_,prod_accum_98__47_,
  prod_accum_98__46_,prod_accum_98__45_,prod_accum_98__44_,prod_accum_98__43_,
  prod_accum_98__42_,prod_accum_98__41_,prod_accum_98__40_,prod_accum_98__39_,
  prod_accum_98__38_,prod_accum_98__37_,prod_accum_98__36_,prod_accum_98__35_,
  prod_accum_98__34_,prod_accum_98__33_,prod_accum_98__32_,prod_accum_98__31_,
  prod_accum_98__30_,prod_accum_98__29_,prod_accum_98__28_,prod_accum_98__27_,prod_accum_98__26_,
  prod_accum_98__25_,prod_accum_98__24_,prod_accum_98__23_,prod_accum_98__22_,
  prod_accum_98__21_,prod_accum_98__20_,prod_accum_98__19_,prod_accum_98__18_,
  prod_accum_98__17_,prod_accum_98__16_,prod_accum_98__15_,prod_accum_98__14_,
  prod_accum_98__13_,prod_accum_98__12_,prod_accum_98__11_,prod_accum_98__10_,prod_accum_98__9_,
  prod_accum_98__8_,prod_accum_98__7_,prod_accum_98__6_,prod_accum_98__5_,
  prod_accum_98__4_,prod_accum_98__3_,prod_accum_98__2_,prod_accum_98__1_,
  prod_accum_98__0_,prod_accum_97__98_,prod_accum_97__97_,prod_accum_97__96_,prod_accum_97__95_,
  prod_accum_97__94_,prod_accum_97__93_,prod_accum_97__92_,prod_accum_97__91_,
  prod_accum_97__90_,prod_accum_97__89_,prod_accum_97__88_,prod_accum_97__87_,
  prod_accum_97__86_,prod_accum_97__85_,prod_accum_97__84_,prod_accum_97__83_,
  prod_accum_97__82_,prod_accum_97__81_,prod_accum_97__80_,prod_accum_97__79_,
  prod_accum_97__78_,prod_accum_97__77_,prod_accum_97__76_,prod_accum_97__75_,prod_accum_97__74_,
  prod_accum_97__73_,prod_accum_97__72_,prod_accum_97__71_,prod_accum_97__70_,
  prod_accum_97__69_,prod_accum_97__68_,prod_accum_97__67_,prod_accum_97__66_,
  prod_accum_97__65_,prod_accum_97__64_,prod_accum_97__63_,prod_accum_97__62_,
  prod_accum_97__61_,prod_accum_97__60_,prod_accum_97__59_,prod_accum_97__58_,prod_accum_97__57_,
  prod_accum_97__56_,prod_accum_97__55_,prod_accum_97__54_,prod_accum_97__53_,
  prod_accum_97__52_,prod_accum_97__51_,prod_accum_97__50_,prod_accum_97__49_,
  prod_accum_97__48_,prod_accum_97__47_,prod_accum_97__46_,prod_accum_97__45_,
  prod_accum_97__44_,prod_accum_97__43_,prod_accum_97__42_,prod_accum_97__41_,
  prod_accum_97__40_,prod_accum_97__39_,prod_accum_97__38_,prod_accum_97__37_,prod_accum_97__36_,
  prod_accum_97__35_,prod_accum_97__34_,prod_accum_97__33_,prod_accum_97__32_,
  prod_accum_97__31_,prod_accum_97__30_,prod_accum_97__29_,prod_accum_97__28_,
  prod_accum_97__27_,prod_accum_97__26_,prod_accum_97__25_,prod_accum_97__24_,
  prod_accum_97__23_,prod_accum_97__22_,prod_accum_97__21_,prod_accum_97__20_,
  prod_accum_97__19_,prod_accum_97__18_,prod_accum_97__17_,prod_accum_97__16_,prod_accum_97__15_,
  prod_accum_97__14_,prod_accum_97__13_,prod_accum_97__12_,prod_accum_97__11_,
  prod_accum_97__10_,prod_accum_97__9_,prod_accum_97__8_,prod_accum_97__7_,
  prod_accum_97__6_,prod_accum_97__5_,prod_accum_97__4_,prod_accum_97__3_,prod_accum_97__2_,
  prod_accum_97__1_,prod_accum_97__0_,prod_accum_96__97_,prod_accum_96__96_,
  prod_accum_96__95_,prod_accum_96__94_,prod_accum_96__93_,prod_accum_96__92_,
  prod_accum_96__91_,prod_accum_96__90_,prod_accum_96__89_,prod_accum_96__88_,
  prod_accum_96__87_,prod_accum_96__86_,prod_accum_96__85_,prod_accum_96__84_,prod_accum_96__83_,
  prod_accum_96__82_,prod_accum_96__81_,prod_accum_96__80_,prod_accum_96__79_,
  prod_accum_96__78_,prod_accum_96__77_,prod_accum_96__76_,prod_accum_96__75_,
  prod_accum_96__74_,prod_accum_96__73_,prod_accum_96__72_,prod_accum_96__71_,
  prod_accum_96__70_,prod_accum_96__69_,prod_accum_96__68_,prod_accum_96__67_,
  prod_accum_96__66_,prod_accum_96__65_,prod_accum_96__64_,prod_accum_96__63_,prod_accum_96__62_,
  prod_accum_96__61_,prod_accum_96__60_,prod_accum_96__59_,prod_accum_96__58_,
  prod_accum_96__57_,prod_accum_96__56_,prod_accum_96__55_,prod_accum_96__54_,
  prod_accum_96__53_,prod_accum_96__52_,prod_accum_96__51_,prod_accum_96__50_,
  prod_accum_96__49_,prod_accum_96__48_,prod_accum_96__47_,prod_accum_96__46_,prod_accum_96__45_,
  prod_accum_96__44_,prod_accum_96__43_,prod_accum_96__42_,prod_accum_96__41_,
  prod_accum_96__40_,prod_accum_96__39_,prod_accum_96__38_,prod_accum_96__37_,
  prod_accum_96__36_,prod_accum_96__35_,prod_accum_96__34_,prod_accum_96__33_,
  prod_accum_96__32_,prod_accum_96__31_,prod_accum_96__30_,prod_accum_96__29_,
  prod_accum_96__28_,prod_accum_96__27_,prod_accum_96__26_,prod_accum_96__25_,prod_accum_96__24_,
  prod_accum_96__23_,prod_accum_96__22_,prod_accum_96__21_,prod_accum_96__20_,
  prod_accum_96__19_,prod_accum_96__18_,prod_accum_96__17_,prod_accum_96__16_,
  prod_accum_96__15_,prod_accum_96__14_,prod_accum_96__13_,prod_accum_96__12_,
  prod_accum_96__11_,prod_accum_96__10_,prod_accum_96__9_,prod_accum_96__8_,prod_accum_96__7_,
  prod_accum_96__6_,prod_accum_96__5_,prod_accum_96__4_,prod_accum_96__3_,
  prod_accum_96__2_,prod_accum_96__1_,prod_accum_96__0_,prod_accum_95__96_,
  prod_accum_95__95_,prod_accum_95__94_,prod_accum_95__93_,prod_accum_95__92_,prod_accum_95__91_,
  prod_accum_95__90_,prod_accum_95__89_,prod_accum_95__88_,prod_accum_95__87_,
  prod_accum_95__86_,prod_accum_95__85_,prod_accum_95__84_,prod_accum_95__83_,
  prod_accum_95__82_,prod_accum_95__81_,prod_accum_95__80_,prod_accum_95__79_,
  prod_accum_95__78_,prod_accum_95__77_,prod_accum_95__76_,prod_accum_95__75_,
  prod_accum_95__74_,prod_accum_95__73_,prod_accum_95__72_,prod_accum_95__71_,prod_accum_95__70_,
  prod_accum_95__69_,prod_accum_95__68_,prod_accum_95__67_,prod_accum_95__66_,
  prod_accum_95__65_,prod_accum_95__64_,prod_accum_95__63_,prod_accum_95__62_,
  prod_accum_95__61_,prod_accum_95__60_,prod_accum_95__59_,prod_accum_95__58_,
  prod_accum_95__57_,prod_accum_95__56_,prod_accum_95__55_,prod_accum_95__54_,
  prod_accum_95__53_,prod_accum_95__52_,prod_accum_95__51_,prod_accum_95__50_,prod_accum_95__49_,
  prod_accum_95__48_,prod_accum_95__47_,prod_accum_95__46_,prod_accum_95__45_,
  prod_accum_95__44_,prod_accum_95__43_,prod_accum_95__42_,prod_accum_95__41_,
  prod_accum_95__40_,prod_accum_95__39_,prod_accum_95__38_,prod_accum_95__37_,
  prod_accum_95__36_,prod_accum_95__35_,prod_accum_95__34_,prod_accum_95__33_,prod_accum_95__32_,
  prod_accum_95__31_,prod_accum_95__30_,prod_accum_95__29_,prod_accum_95__28_,
  prod_accum_95__27_,prod_accum_95__26_,prod_accum_95__25_,prod_accum_95__24_,
  prod_accum_95__23_,prod_accum_95__22_,prod_accum_95__21_,prod_accum_95__20_,
  prod_accum_95__19_,prod_accum_95__18_,prod_accum_95__17_,prod_accum_95__16_,
  prod_accum_95__15_,prod_accum_95__14_,prod_accum_95__13_,prod_accum_95__12_,prod_accum_95__11_,
  prod_accum_95__10_,prod_accum_95__9_,prod_accum_95__8_,prod_accum_95__7_,
  prod_accum_95__6_,prod_accum_95__5_,prod_accum_95__4_,prod_accum_95__3_,
  prod_accum_95__2_,prod_accum_95__1_,prod_accum_95__0_,s_r_102__127_,s_r_102__126_,s_r_102__125_,
  s_r_102__124_,s_r_102__123_,s_r_102__122_,s_r_102__121_,s_r_102__120_,
  s_r_102__119_,s_r_102__118_,s_r_102__117_,s_r_102__116_,s_r_102__115_,s_r_102__114_,
  s_r_102__113_,s_r_102__112_,s_r_102__111_,s_r_102__110_,s_r_102__109_,s_r_102__108_,
  s_r_102__107_,s_r_102__106_,s_r_102__105_,s_r_102__104_,s_r_102__103_,
  s_r_102__102_,s_r_102__101_,s_r_102__100_,s_r_102__99_,s_r_102__98_,s_r_102__97_,
  s_r_102__96_,s_r_102__95_,s_r_102__94_,s_r_102__93_,s_r_102__92_,s_r_102__91_,s_r_102__90_,
  s_r_102__89_,s_r_102__88_,s_r_102__87_,s_r_102__86_,s_r_102__85_,s_r_102__84_,
  s_r_102__83_,s_r_102__82_,s_r_102__81_,s_r_102__80_,s_r_102__79_,s_r_102__78_,
  s_r_102__77_,s_r_102__76_,s_r_102__75_,s_r_102__74_,s_r_102__73_,s_r_102__72_,
  s_r_102__71_,s_r_102__70_,s_r_102__69_,s_r_102__68_,s_r_102__67_,s_r_102__66_,
  s_r_102__65_,s_r_102__64_,s_r_102__63_,s_r_102__62_,s_r_102__61_,s_r_102__60_,
  s_r_102__59_,s_r_102__58_,s_r_102__57_,s_r_102__56_,s_r_102__55_,s_r_102__54_,
  s_r_102__53_,s_r_102__52_,s_r_102__51_,s_r_102__50_,s_r_102__49_,s_r_102__48_,s_r_102__47_,
  s_r_102__46_,s_r_102__45_,s_r_102__44_,s_r_102__43_,s_r_102__42_,s_r_102__41_,
  s_r_102__40_,s_r_102__39_,s_r_102__38_,s_r_102__37_,s_r_102__36_,s_r_102__35_,
  s_r_102__34_,s_r_102__33_,s_r_102__32_,s_r_102__31_,s_r_102__30_,s_r_102__29_,
  s_r_102__28_,s_r_102__27_,s_r_102__26_,s_r_102__25_,s_r_102__24_,s_r_102__23_,
  s_r_102__22_,s_r_102__21_,s_r_102__20_,s_r_102__19_,s_r_102__18_,s_r_102__17_,
  s_r_102__16_,s_r_102__15_,s_r_102__14_,s_r_102__13_,s_r_102__12_,s_r_102__11_,s_r_102__10_,
  s_r_102__9_,s_r_102__8_,s_r_102__7_,s_r_102__6_,s_r_102__5_,s_r_102__4_,
  s_r_102__3_,s_r_102__2_,s_r_102__1_,s_r_102__0_,s_r_101__127_,s_r_101__126_,
  s_r_101__125_,s_r_101__124_,s_r_101__123_,s_r_101__122_,s_r_101__121_,s_r_101__120_,
  s_r_101__119_,s_r_101__118_,s_r_101__117_,s_r_101__116_,s_r_101__115_,s_r_101__114_,
  s_r_101__113_,s_r_101__112_,s_r_101__111_,s_r_101__110_,s_r_101__109_,s_r_101__108_,
  s_r_101__107_,s_r_101__106_,s_r_101__105_,s_r_101__104_,s_r_101__103_,
  s_r_101__102_,s_r_101__101_,s_r_101__100_,s_r_101__99_,s_r_101__98_,s_r_101__97_,
  s_r_101__96_,s_r_101__95_,s_r_101__94_,s_r_101__93_,s_r_101__92_,s_r_101__91_,
  s_r_101__90_,s_r_101__89_,s_r_101__88_,s_r_101__87_,s_r_101__86_,s_r_101__85_,s_r_101__84_,
  s_r_101__83_,s_r_101__82_,s_r_101__81_,s_r_101__80_,s_r_101__79_,s_r_101__78_,
  s_r_101__77_,s_r_101__76_,s_r_101__75_,s_r_101__74_,s_r_101__73_,s_r_101__72_,
  s_r_101__71_,s_r_101__70_,s_r_101__69_,s_r_101__68_,s_r_101__67_,s_r_101__66_,
  s_r_101__65_,s_r_101__64_,s_r_101__63_,s_r_101__62_,s_r_101__61_,s_r_101__60_,
  s_r_101__59_,s_r_101__58_,s_r_101__57_,s_r_101__56_,s_r_101__55_,s_r_101__54_,
  s_r_101__53_,s_r_101__52_,s_r_101__51_,s_r_101__50_,s_r_101__49_,s_r_101__48_,
  s_r_101__47_,s_r_101__46_,s_r_101__45_,s_r_101__44_,s_r_101__43_,s_r_101__42_,s_r_101__41_,
  s_r_101__40_,s_r_101__39_,s_r_101__38_,s_r_101__37_,s_r_101__36_,s_r_101__35_,
  s_r_101__34_,s_r_101__33_,s_r_101__32_,s_r_101__31_,s_r_101__30_,s_r_101__29_,
  s_r_101__28_,s_r_101__27_,s_r_101__26_,s_r_101__25_,s_r_101__24_,s_r_101__23_,
  s_r_101__22_,s_r_101__21_,s_r_101__20_,s_r_101__19_,s_r_101__18_,s_r_101__17_,
  s_r_101__16_,s_r_101__15_,s_r_101__14_,s_r_101__13_,s_r_101__12_,s_r_101__11_,
  s_r_101__10_,s_r_101__9_,s_r_101__8_,s_r_101__7_,s_r_101__6_,s_r_101__5_,s_r_101__4_,
  s_r_101__3_,s_r_101__2_,s_r_101__1_,s_r_101__0_,s_r_100__127_,s_r_100__126_,
  s_r_100__125_,s_r_100__124_,s_r_100__123_,s_r_100__122_,s_r_100__121_,s_r_100__120_,
  s_r_100__119_,s_r_100__118_,s_r_100__117_,s_r_100__116_,s_r_100__115_,s_r_100__114_,
  s_r_100__113_,s_r_100__112_,s_r_100__111_,s_r_100__110_,s_r_100__109_,
  s_r_100__108_,s_r_100__107_,s_r_100__106_,s_r_100__105_,s_r_100__104_,s_r_100__103_,
  s_r_100__102_,s_r_100__101_,s_r_100__100_,s_r_100__99_,s_r_100__98_,s_r_100__97_,
  s_r_100__96_,s_r_100__95_,s_r_100__94_,s_r_100__93_,s_r_100__92_,s_r_100__91_,
  s_r_100__90_,s_r_100__89_,s_r_100__88_,s_r_100__87_,s_r_100__86_,s_r_100__85_,
  s_r_100__84_,s_r_100__83_,s_r_100__82_,s_r_100__81_,s_r_100__80_,s_r_100__79_,s_r_100__78_,
  s_r_100__77_,s_r_100__76_,s_r_100__75_,s_r_100__74_,s_r_100__73_,s_r_100__72_,
  s_r_100__71_,s_r_100__70_,s_r_100__69_,s_r_100__68_,s_r_100__67_,s_r_100__66_,
  s_r_100__65_,s_r_100__64_,s_r_100__63_,s_r_100__62_,s_r_100__61_,s_r_100__60_,
  s_r_100__59_,s_r_100__58_,s_r_100__57_,s_r_100__56_,s_r_100__55_,s_r_100__54_,
  s_r_100__53_,s_r_100__52_,s_r_100__51_,s_r_100__50_,s_r_100__49_,s_r_100__48_,
  s_r_100__47_,s_r_100__46_,s_r_100__45_,s_r_100__44_,s_r_100__43_,s_r_100__42_,
  s_r_100__41_,s_r_100__40_,s_r_100__39_,s_r_100__38_,s_r_100__37_,s_r_100__36_,s_r_100__35_,
  s_r_100__34_,s_r_100__33_,s_r_100__32_,s_r_100__31_,s_r_100__30_,s_r_100__29_,
  s_r_100__28_,s_r_100__27_,s_r_100__26_,s_r_100__25_,s_r_100__24_,s_r_100__23_,
  s_r_100__22_,s_r_100__21_,s_r_100__20_,s_r_100__19_,s_r_100__18_,s_r_100__17_,
  s_r_100__16_,s_r_100__15_,s_r_100__14_,s_r_100__13_,s_r_100__12_,s_r_100__11_,
  s_r_100__10_,s_r_100__9_,s_r_100__8_,s_r_100__7_,s_r_100__6_,s_r_100__5_,s_r_100__4_,
  s_r_100__3_,s_r_100__2_,s_r_100__1_,s_r_100__0_,s_r_99__127_,s_r_99__126_,
  s_r_99__125_,s_r_99__124_,s_r_99__123_,s_r_99__122_,s_r_99__121_,s_r_99__120_,
  s_r_99__119_,s_r_99__118_,s_r_99__117_,s_r_99__116_,s_r_99__115_,s_r_99__114_,s_r_99__113_,
  s_r_99__112_,s_r_99__111_,s_r_99__110_,s_r_99__109_,s_r_99__108_,s_r_99__107_,
  s_r_99__106_,s_r_99__105_,s_r_99__104_,s_r_99__103_,s_r_99__102_,s_r_99__101_,
  s_r_99__100_,s_r_99__99_,s_r_99__98_,s_r_99__97_,s_r_99__96_,s_r_99__95_,s_r_99__94_,
  s_r_99__93_,s_r_99__92_,s_r_99__91_,s_r_99__90_,s_r_99__89_,s_r_99__88_,
  s_r_99__87_,s_r_99__86_,s_r_99__85_,s_r_99__84_,s_r_99__83_,s_r_99__82_,s_r_99__81_,
  s_r_99__80_,s_r_99__79_,s_r_99__78_,s_r_99__77_,s_r_99__76_,s_r_99__75_,s_r_99__74_,
  s_r_99__73_,s_r_99__72_,s_r_99__71_,s_r_99__70_,s_r_99__69_,s_r_99__68_,
  s_r_99__67_,s_r_99__66_,s_r_99__65_,s_r_99__64_,s_r_99__63_,s_r_99__62_,s_r_99__61_,
  s_r_99__60_,s_r_99__59_,s_r_99__58_,s_r_99__57_,s_r_99__56_,s_r_99__55_,s_r_99__54_,
  s_r_99__53_,s_r_99__52_,s_r_99__51_,s_r_99__50_,s_r_99__49_,s_r_99__48_,
  s_r_99__47_,s_r_99__46_,s_r_99__45_,s_r_99__44_,s_r_99__43_,s_r_99__42_,s_r_99__41_,
  s_r_99__40_,s_r_99__39_,s_r_99__38_,s_r_99__37_,s_r_99__36_,s_r_99__35_,s_r_99__34_,
  s_r_99__33_,s_r_99__32_,s_r_99__31_,s_r_99__30_,s_r_99__29_,s_r_99__28_,
  s_r_99__27_,s_r_99__26_,s_r_99__25_,s_r_99__24_,s_r_99__23_,s_r_99__22_,s_r_99__21_,
  s_r_99__20_,s_r_99__19_,s_r_99__18_,s_r_99__17_,s_r_99__16_,s_r_99__15_,s_r_99__14_,
  s_r_99__13_,s_r_99__12_,s_r_99__11_,s_r_99__10_,s_r_99__9_,s_r_99__8_,
  s_r_99__7_,s_r_99__6_,s_r_99__5_,s_r_99__4_,s_r_99__3_,s_r_99__2_,s_r_99__1_,s_r_99__0_,
  prod_accum_102__103_,prod_accum_102__102_,prod_accum_102__101_,
  prod_accum_102__100_,prod_accum_102__99_,prod_accum_102__98_,prod_accum_102__97_,
  prod_accum_102__96_,prod_accum_102__95_,prod_accum_102__94_,prod_accum_102__93_,
  prod_accum_102__92_,prod_accum_102__91_,prod_accum_102__90_,prod_accum_102__89_,
  prod_accum_102__88_,prod_accum_102__87_,prod_accum_102__86_,prod_accum_102__85_,
  prod_accum_102__84_,prod_accum_102__83_,prod_accum_102__82_,prod_accum_102__81_,
  prod_accum_102__80_,prod_accum_102__79_,prod_accum_102__78_,prod_accum_102__77_,
  prod_accum_102__76_,prod_accum_102__75_,prod_accum_102__74_,prod_accum_102__73_,
  prod_accum_102__72_,prod_accum_102__71_,prod_accum_102__70_,prod_accum_102__69_,
  prod_accum_102__68_,prod_accum_102__67_,prod_accum_102__66_,prod_accum_102__65_,
  prod_accum_102__64_,prod_accum_102__63_,prod_accum_102__62_,prod_accum_102__61_,
  prod_accum_102__60_,prod_accum_102__59_,prod_accum_102__58_,prod_accum_102__57_,
  prod_accum_102__56_,prod_accum_102__55_,prod_accum_102__54_,prod_accum_102__53_,
  prod_accum_102__52_,prod_accum_102__51_,prod_accum_102__50_,prod_accum_102__49_,
  prod_accum_102__48_,prod_accum_102__47_,prod_accum_102__46_,prod_accum_102__45_,
  prod_accum_102__44_,prod_accum_102__43_,prod_accum_102__42_,prod_accum_102__41_,
  prod_accum_102__40_,prod_accum_102__39_,prod_accum_102__38_,prod_accum_102__37_,
  prod_accum_102__36_,prod_accum_102__35_,prod_accum_102__34_,prod_accum_102__33_,
  prod_accum_102__32_,prod_accum_102__31_,prod_accum_102__30_,prod_accum_102__29_,
  prod_accum_102__28_,prod_accum_102__27_,prod_accum_102__26_,prod_accum_102__25_,
  prod_accum_102__24_,prod_accum_102__23_,prod_accum_102__22_,prod_accum_102__21_,
  prod_accum_102__20_,prod_accum_102__19_,prod_accum_102__18_,prod_accum_102__17_,
  prod_accum_102__16_,prod_accum_102__15_,prod_accum_102__14_,prod_accum_102__13_,
  prod_accum_102__12_,prod_accum_102__11_,prod_accum_102__10_,prod_accum_102__9_,prod_accum_102__8_,
  prod_accum_102__7_,prod_accum_102__6_,prod_accum_102__5_,prod_accum_102__4_,
  prod_accum_102__3_,prod_accum_102__2_,prod_accum_102__1_,prod_accum_102__0_,
  prod_accum_101__102_,prod_accum_101__101_,prod_accum_101__100_,prod_accum_101__99_,
  prod_accum_101__98_,prod_accum_101__97_,prod_accum_101__96_,prod_accum_101__95_,
  prod_accum_101__94_,prod_accum_101__93_,prod_accum_101__92_,prod_accum_101__91_,
  prod_accum_101__90_,prod_accum_101__89_,prod_accum_101__88_,prod_accum_101__87_,
  prod_accum_101__86_,prod_accum_101__85_,prod_accum_101__84_,prod_accum_101__83_,
  prod_accum_101__82_,prod_accum_101__81_,prod_accum_101__80_,prod_accum_101__79_,
  prod_accum_101__78_,prod_accum_101__77_,prod_accum_101__76_,prod_accum_101__75_,
  prod_accum_101__74_,prod_accum_101__73_,prod_accum_101__72_,prod_accum_101__71_,
  prod_accum_101__70_,prod_accum_101__69_,prod_accum_101__68_,prod_accum_101__67_,
  prod_accum_101__66_,prod_accum_101__65_,prod_accum_101__64_,prod_accum_101__63_,
  prod_accum_101__62_,prod_accum_101__61_,prod_accum_101__60_,prod_accum_101__59_,
  prod_accum_101__58_,prod_accum_101__57_,prod_accum_101__56_,prod_accum_101__55_,
  prod_accum_101__54_,prod_accum_101__53_,prod_accum_101__52_,prod_accum_101__51_,
  prod_accum_101__50_,prod_accum_101__49_,prod_accum_101__48_,prod_accum_101__47_,
  prod_accum_101__46_,prod_accum_101__45_,prod_accum_101__44_,prod_accum_101__43_,
  prod_accum_101__42_,prod_accum_101__41_,prod_accum_101__40_,prod_accum_101__39_,
  prod_accum_101__38_,prod_accum_101__37_,prod_accum_101__36_,prod_accum_101__35_,
  prod_accum_101__34_,prod_accum_101__33_,prod_accum_101__32_,prod_accum_101__31_,
  prod_accum_101__30_,prod_accum_101__29_,prod_accum_101__28_,prod_accum_101__27_,
  prod_accum_101__26_,prod_accum_101__25_,prod_accum_101__24_,prod_accum_101__23_,
  prod_accum_101__22_,prod_accum_101__21_,prod_accum_101__20_,prod_accum_101__19_,
  prod_accum_101__18_,prod_accum_101__17_,prod_accum_101__16_,prod_accum_101__15_,
  prod_accum_101__14_,prod_accum_101__13_,prod_accum_101__12_,prod_accum_101__11_,
  prod_accum_101__10_,prod_accum_101__9_,prod_accum_101__8_,prod_accum_101__7_,
  prod_accum_101__6_,prod_accum_101__5_,prod_accum_101__4_,prod_accum_101__3_,
  prod_accum_101__2_,prod_accum_101__1_,prod_accum_101__0_,prod_accum_100__101_,
  prod_accum_100__100_,prod_accum_100__99_,prod_accum_100__98_,prod_accum_100__97_,
  prod_accum_100__96_,prod_accum_100__95_,prod_accum_100__94_,prod_accum_100__93_,
  prod_accum_100__92_,prod_accum_100__91_,prod_accum_100__90_,prod_accum_100__89_,
  prod_accum_100__88_,prod_accum_100__87_,prod_accum_100__86_,prod_accum_100__85_,
  prod_accum_100__84_,prod_accum_100__83_,prod_accum_100__82_,prod_accum_100__81_,
  prod_accum_100__80_,prod_accum_100__79_,prod_accum_100__78_,prod_accum_100__77_,
  prod_accum_100__76_,prod_accum_100__75_,prod_accum_100__74_,prod_accum_100__73_,
  prod_accum_100__72_,prod_accum_100__71_,prod_accum_100__70_,prod_accum_100__69_,
  prod_accum_100__68_,prod_accum_100__67_,prod_accum_100__66_,prod_accum_100__65_,
  prod_accum_100__64_,prod_accum_100__63_,prod_accum_100__62_,prod_accum_100__61_,
  prod_accum_100__60_,prod_accum_100__59_,prod_accum_100__58_,prod_accum_100__57_,
  prod_accum_100__56_,prod_accum_100__55_,prod_accum_100__54_,prod_accum_100__53_,
  prod_accum_100__52_,prod_accum_100__51_,prod_accum_100__50_,prod_accum_100__49_,
  prod_accum_100__48_,prod_accum_100__47_,prod_accum_100__46_,prod_accum_100__45_,
  prod_accum_100__44_,prod_accum_100__43_,prod_accum_100__42_,prod_accum_100__41_,
  prod_accum_100__40_,prod_accum_100__39_,prod_accum_100__38_,prod_accum_100__37_,
  prod_accum_100__36_,prod_accum_100__35_,prod_accum_100__34_,prod_accum_100__33_,
  prod_accum_100__32_,prod_accum_100__31_,prod_accum_100__30_,prod_accum_100__29_,
  prod_accum_100__28_,prod_accum_100__27_,prod_accum_100__26_,prod_accum_100__25_,
  prod_accum_100__24_,prod_accum_100__23_,prod_accum_100__22_,prod_accum_100__21_,
  prod_accum_100__20_,prod_accum_100__19_,prod_accum_100__18_,prod_accum_100__17_,
  prod_accum_100__16_,prod_accum_100__15_,prod_accum_100__14_,prod_accum_100__13_,
  prod_accum_100__12_,prod_accum_100__11_,prod_accum_100__10_,prod_accum_100__9_,
  prod_accum_100__8_,prod_accum_100__7_,prod_accum_100__6_,prod_accum_100__5_,
  prod_accum_100__4_,prod_accum_100__3_,prod_accum_100__2_,prod_accum_100__1_,prod_accum_100__0_,
  prod_accum_99__100_,prod_accum_99__99_,prod_accum_99__98_,prod_accum_99__97_,
  prod_accum_99__96_,prod_accum_99__95_,prod_accum_99__94_,prod_accum_99__93_,
  prod_accum_99__92_,prod_accum_99__91_,prod_accum_99__90_,prod_accum_99__89_,
  prod_accum_99__88_,prod_accum_99__87_,prod_accum_99__86_,prod_accum_99__85_,
  prod_accum_99__84_,prod_accum_99__83_,prod_accum_99__82_,prod_accum_99__81_,prod_accum_99__80_,
  prod_accum_99__79_,prod_accum_99__78_,prod_accum_99__77_,prod_accum_99__76_,
  prod_accum_99__75_,prod_accum_99__74_,prod_accum_99__73_,prod_accum_99__72_,
  prod_accum_99__71_,prod_accum_99__70_,prod_accum_99__69_,prod_accum_99__68_,
  prod_accum_99__67_,prod_accum_99__66_,prod_accum_99__65_,prod_accum_99__64_,prod_accum_99__63_,
  prod_accum_99__62_,prod_accum_99__61_,prod_accum_99__60_,prod_accum_99__59_,
  prod_accum_99__58_,prod_accum_99__57_,prod_accum_99__56_,prod_accum_99__55_,
  prod_accum_99__54_,prod_accum_99__53_,prod_accum_99__52_,prod_accum_99__51_,
  prod_accum_99__50_,prod_accum_99__49_,prod_accum_99__48_,prod_accum_99__47_,
  prod_accum_99__46_,prod_accum_99__45_,prod_accum_99__44_,prod_accum_99__43_,prod_accum_99__42_,
  prod_accum_99__41_,prod_accum_99__40_,prod_accum_99__39_,prod_accum_99__38_,
  prod_accum_99__37_,prod_accum_99__36_,prod_accum_99__35_,prod_accum_99__34_,
  prod_accum_99__33_,prod_accum_99__32_,prod_accum_99__31_,prod_accum_99__30_,
  prod_accum_99__29_,prod_accum_99__28_,prod_accum_99__27_,prod_accum_99__26_,
  prod_accum_99__25_,prod_accum_99__24_,prod_accum_99__23_,prod_accum_99__22_,prod_accum_99__21_,
  prod_accum_99__20_,prod_accum_99__19_,prod_accum_99__18_,prod_accum_99__17_,
  prod_accum_99__16_,prod_accum_99__15_,prod_accum_99__14_,prod_accum_99__13_,
  prod_accum_99__12_,prod_accum_99__11_,prod_accum_99__10_,prod_accum_99__9_,
  prod_accum_99__8_,prod_accum_99__7_,prod_accum_99__6_,prod_accum_99__5_,prod_accum_99__4_,
  prod_accum_99__3_,prod_accum_99__2_,prod_accum_99__1_,prod_accum_99__0_,
  s_r_106__127_,s_r_106__126_,s_r_106__125_,s_r_106__124_,s_r_106__123_,s_r_106__122_,
  s_r_106__121_,s_r_106__120_,s_r_106__119_,s_r_106__118_,s_r_106__117_,s_r_106__116_,
  s_r_106__115_,s_r_106__114_,s_r_106__113_,s_r_106__112_,s_r_106__111_,s_r_106__110_,
  s_r_106__109_,s_r_106__108_,s_r_106__107_,s_r_106__106_,s_r_106__105_,
  s_r_106__104_,s_r_106__103_,s_r_106__102_,s_r_106__101_,s_r_106__100_,s_r_106__99_,
  s_r_106__98_,s_r_106__97_,s_r_106__96_,s_r_106__95_,s_r_106__94_,s_r_106__93_,
  s_r_106__92_,s_r_106__91_,s_r_106__90_,s_r_106__89_,s_r_106__88_,s_r_106__87_,
  s_r_106__86_,s_r_106__85_,s_r_106__84_,s_r_106__83_,s_r_106__82_,s_r_106__81_,s_r_106__80_,
  s_r_106__79_,s_r_106__78_,s_r_106__77_,s_r_106__76_,s_r_106__75_,s_r_106__74_,
  s_r_106__73_,s_r_106__72_,s_r_106__71_,s_r_106__70_,s_r_106__69_,s_r_106__68_,
  s_r_106__67_,s_r_106__66_,s_r_106__65_,s_r_106__64_,s_r_106__63_,s_r_106__62_,
  s_r_106__61_,s_r_106__60_,s_r_106__59_,s_r_106__58_,s_r_106__57_,s_r_106__56_,
  s_r_106__55_,s_r_106__54_,s_r_106__53_,s_r_106__52_,s_r_106__51_,s_r_106__50_,
  s_r_106__49_,s_r_106__48_,s_r_106__47_,s_r_106__46_,s_r_106__45_,s_r_106__44_,s_r_106__43_,
  s_r_106__42_,s_r_106__41_,s_r_106__40_,s_r_106__39_,s_r_106__38_,s_r_106__37_,
  s_r_106__36_,s_r_106__35_,s_r_106__34_,s_r_106__33_,s_r_106__32_,s_r_106__31_,
  s_r_106__30_,s_r_106__29_,s_r_106__28_,s_r_106__27_,s_r_106__26_,s_r_106__25_,
  s_r_106__24_,s_r_106__23_,s_r_106__22_,s_r_106__21_,s_r_106__20_,s_r_106__19_,
  s_r_106__18_,s_r_106__17_,s_r_106__16_,s_r_106__15_,s_r_106__14_,s_r_106__13_,
  s_r_106__12_,s_r_106__11_,s_r_106__10_,s_r_106__9_,s_r_106__8_,s_r_106__7_,s_r_106__6_,
  s_r_106__5_,s_r_106__4_,s_r_106__3_,s_r_106__2_,s_r_106__1_,s_r_106__0_,
  s_r_105__127_,s_r_105__126_,s_r_105__125_,s_r_105__124_,s_r_105__123_,s_r_105__122_,
  s_r_105__121_,s_r_105__120_,s_r_105__119_,s_r_105__118_,s_r_105__117_,s_r_105__116_,
  s_r_105__115_,s_r_105__114_,s_r_105__113_,s_r_105__112_,s_r_105__111_,
  s_r_105__110_,s_r_105__109_,s_r_105__108_,s_r_105__107_,s_r_105__106_,s_r_105__105_,
  s_r_105__104_,s_r_105__103_,s_r_105__102_,s_r_105__101_,s_r_105__100_,s_r_105__99_,
  s_r_105__98_,s_r_105__97_,s_r_105__96_,s_r_105__95_,s_r_105__94_,s_r_105__93_,
  s_r_105__92_,s_r_105__91_,s_r_105__90_,s_r_105__89_,s_r_105__88_,s_r_105__87_,
  s_r_105__86_,s_r_105__85_,s_r_105__84_,s_r_105__83_,s_r_105__82_,s_r_105__81_,
  s_r_105__80_,s_r_105__79_,s_r_105__78_,s_r_105__77_,s_r_105__76_,s_r_105__75_,s_r_105__74_,
  s_r_105__73_,s_r_105__72_,s_r_105__71_,s_r_105__70_,s_r_105__69_,s_r_105__68_,
  s_r_105__67_,s_r_105__66_,s_r_105__65_,s_r_105__64_,s_r_105__63_,s_r_105__62_,
  s_r_105__61_,s_r_105__60_,s_r_105__59_,s_r_105__58_,s_r_105__57_,s_r_105__56_,
  s_r_105__55_,s_r_105__54_,s_r_105__53_,s_r_105__52_,s_r_105__51_,s_r_105__50_,
  s_r_105__49_,s_r_105__48_,s_r_105__47_,s_r_105__46_,s_r_105__45_,s_r_105__44_,
  s_r_105__43_,s_r_105__42_,s_r_105__41_,s_r_105__40_,s_r_105__39_,s_r_105__38_,s_r_105__37_,
  s_r_105__36_,s_r_105__35_,s_r_105__34_,s_r_105__33_,s_r_105__32_,s_r_105__31_,
  s_r_105__30_,s_r_105__29_,s_r_105__28_,s_r_105__27_,s_r_105__26_,s_r_105__25_,
  s_r_105__24_,s_r_105__23_,s_r_105__22_,s_r_105__21_,s_r_105__20_,s_r_105__19_,
  s_r_105__18_,s_r_105__17_,s_r_105__16_,s_r_105__15_,s_r_105__14_,s_r_105__13_,
  s_r_105__12_,s_r_105__11_,s_r_105__10_,s_r_105__9_,s_r_105__8_,s_r_105__7_,s_r_105__6_,
  s_r_105__5_,s_r_105__4_,s_r_105__3_,s_r_105__2_,s_r_105__1_,s_r_105__0_,
  s_r_104__127_,s_r_104__126_,s_r_104__125_,s_r_104__124_,s_r_104__123_,s_r_104__122_,
  s_r_104__121_,s_r_104__120_,s_r_104__119_,s_r_104__118_,s_r_104__117_,s_r_104__116_,
  s_r_104__115_,s_r_104__114_,s_r_104__113_,s_r_104__112_,s_r_104__111_,
  s_r_104__110_,s_r_104__109_,s_r_104__108_,s_r_104__107_,s_r_104__106_,s_r_104__105_,
  s_r_104__104_,s_r_104__103_,s_r_104__102_,s_r_104__101_,s_r_104__100_,s_r_104__99_,
  s_r_104__98_,s_r_104__97_,s_r_104__96_,s_r_104__95_,s_r_104__94_,s_r_104__93_,
  s_r_104__92_,s_r_104__91_,s_r_104__90_,s_r_104__89_,s_r_104__88_,s_r_104__87_,
  s_r_104__86_,s_r_104__85_,s_r_104__84_,s_r_104__83_,s_r_104__82_,s_r_104__81_,
  s_r_104__80_,s_r_104__79_,s_r_104__78_,s_r_104__77_,s_r_104__76_,s_r_104__75_,
  s_r_104__74_,s_r_104__73_,s_r_104__72_,s_r_104__71_,s_r_104__70_,s_r_104__69_,s_r_104__68_,
  s_r_104__67_,s_r_104__66_,s_r_104__65_,s_r_104__64_,s_r_104__63_,s_r_104__62_,
  s_r_104__61_,s_r_104__60_,s_r_104__59_,s_r_104__58_,s_r_104__57_,s_r_104__56_,
  s_r_104__55_,s_r_104__54_,s_r_104__53_,s_r_104__52_,s_r_104__51_,s_r_104__50_,
  s_r_104__49_,s_r_104__48_,s_r_104__47_,s_r_104__46_,s_r_104__45_,s_r_104__44_,
  s_r_104__43_,s_r_104__42_,s_r_104__41_,s_r_104__40_,s_r_104__39_,s_r_104__38_,
  s_r_104__37_,s_r_104__36_,s_r_104__35_,s_r_104__34_,s_r_104__33_,s_r_104__32_,s_r_104__31_,
  s_r_104__30_,s_r_104__29_,s_r_104__28_,s_r_104__27_,s_r_104__26_,s_r_104__25_,
  s_r_104__24_,s_r_104__23_,s_r_104__22_,s_r_104__21_,s_r_104__20_,s_r_104__19_,
  s_r_104__18_,s_r_104__17_,s_r_104__16_,s_r_104__15_,s_r_104__14_,s_r_104__13_,
  s_r_104__12_,s_r_104__11_,s_r_104__10_,s_r_104__9_,s_r_104__8_,s_r_104__7_,
  s_r_104__6_,s_r_104__5_,s_r_104__4_,s_r_104__3_,s_r_104__2_,s_r_104__1_,s_r_104__0_,
  s_r_103__127_,s_r_103__126_,s_r_103__125_,s_r_103__124_,s_r_103__123_,s_r_103__122_,
  s_r_103__121_,s_r_103__120_,s_r_103__119_,s_r_103__118_,s_r_103__117_,
  s_r_103__116_,s_r_103__115_,s_r_103__114_,s_r_103__113_,s_r_103__112_,s_r_103__111_,
  s_r_103__110_,s_r_103__109_,s_r_103__108_,s_r_103__107_,s_r_103__106_,s_r_103__105_,
  s_r_103__104_,s_r_103__103_,s_r_103__102_,s_r_103__101_,s_r_103__100_,s_r_103__99_,
  s_r_103__98_,s_r_103__97_,s_r_103__96_,s_r_103__95_,s_r_103__94_,s_r_103__93_,
  s_r_103__92_,s_r_103__91_,s_r_103__90_,s_r_103__89_,s_r_103__88_,s_r_103__87_,
  s_r_103__86_,s_r_103__85_,s_r_103__84_,s_r_103__83_,s_r_103__82_,s_r_103__81_,
  s_r_103__80_,s_r_103__79_,s_r_103__78_,s_r_103__77_,s_r_103__76_,s_r_103__75_,
  s_r_103__74_,s_r_103__73_,s_r_103__72_,s_r_103__71_,s_r_103__70_,s_r_103__69_,
  s_r_103__68_,s_r_103__67_,s_r_103__66_,s_r_103__65_,s_r_103__64_,s_r_103__63_,s_r_103__62_,
  s_r_103__61_,s_r_103__60_,s_r_103__59_,s_r_103__58_,s_r_103__57_,s_r_103__56_,
  s_r_103__55_,s_r_103__54_,s_r_103__53_,s_r_103__52_,s_r_103__51_,s_r_103__50_,
  s_r_103__49_,s_r_103__48_,s_r_103__47_,s_r_103__46_,s_r_103__45_,s_r_103__44_,
  s_r_103__43_,s_r_103__42_,s_r_103__41_,s_r_103__40_,s_r_103__39_,s_r_103__38_,
  s_r_103__37_,s_r_103__36_,s_r_103__35_,s_r_103__34_,s_r_103__33_,s_r_103__32_,
  s_r_103__31_,s_r_103__30_,s_r_103__29_,s_r_103__28_,s_r_103__27_,s_r_103__26_,s_r_103__25_,
  s_r_103__24_,s_r_103__23_,s_r_103__22_,s_r_103__21_,s_r_103__20_,s_r_103__19_,
  s_r_103__18_,s_r_103__17_,s_r_103__16_,s_r_103__15_,s_r_103__14_,s_r_103__13_,
  s_r_103__12_,s_r_103__11_,s_r_103__10_,s_r_103__9_,s_r_103__8_,s_r_103__7_,
  s_r_103__6_,s_r_103__5_,s_r_103__4_,s_r_103__3_,s_r_103__2_,s_r_103__1_,s_r_103__0_,
  prod_accum_106__107_,prod_accum_106__106_,prod_accum_106__105_,prod_accum_106__104_,
  prod_accum_106__103_,prod_accum_106__102_,prod_accum_106__101_,
  prod_accum_106__100_,prod_accum_106__99_,prod_accum_106__98_,prod_accum_106__97_,
  prod_accum_106__96_,prod_accum_106__95_,prod_accum_106__94_,prod_accum_106__93_,
  prod_accum_106__92_,prod_accum_106__91_,prod_accum_106__90_,prod_accum_106__89_,
  prod_accum_106__88_,prod_accum_106__87_,prod_accum_106__86_,prod_accum_106__85_,
  prod_accum_106__84_,prod_accum_106__83_,prod_accum_106__82_,prod_accum_106__81_,
  prod_accum_106__80_,prod_accum_106__79_,prod_accum_106__78_,prod_accum_106__77_,
  prod_accum_106__76_,prod_accum_106__75_,prod_accum_106__74_,prod_accum_106__73_,
  prod_accum_106__72_,prod_accum_106__71_,prod_accum_106__70_,prod_accum_106__69_,
  prod_accum_106__68_,prod_accum_106__67_,prod_accum_106__66_,prod_accum_106__65_,
  prod_accum_106__64_,prod_accum_106__63_,prod_accum_106__62_,prod_accum_106__61_,
  prod_accum_106__60_,prod_accum_106__59_,prod_accum_106__58_,prod_accum_106__57_,
  prod_accum_106__56_,prod_accum_106__55_,prod_accum_106__54_,prod_accum_106__53_,
  prod_accum_106__52_,prod_accum_106__51_,prod_accum_106__50_,prod_accum_106__49_,
  prod_accum_106__48_,prod_accum_106__47_,prod_accum_106__46_,prod_accum_106__45_,
  prod_accum_106__44_,prod_accum_106__43_,prod_accum_106__42_,prod_accum_106__41_,
  prod_accum_106__40_,prod_accum_106__39_,prod_accum_106__38_,prod_accum_106__37_,
  prod_accum_106__36_,prod_accum_106__35_,prod_accum_106__34_,prod_accum_106__33_,
  prod_accum_106__32_,prod_accum_106__31_,prod_accum_106__30_,prod_accum_106__29_,
  prod_accum_106__28_,prod_accum_106__27_,prod_accum_106__26_,prod_accum_106__25_,
  prod_accum_106__24_,prod_accum_106__23_,prod_accum_106__22_,prod_accum_106__21_,
  prod_accum_106__20_,prod_accum_106__19_,prod_accum_106__18_,prod_accum_106__17_,
  prod_accum_106__16_,prod_accum_106__15_,prod_accum_106__14_,prod_accum_106__13_,
  prod_accum_106__12_,prod_accum_106__11_,prod_accum_106__10_,prod_accum_106__9_,
  prod_accum_106__8_,prod_accum_106__7_,prod_accum_106__6_,prod_accum_106__5_,prod_accum_106__4_,
  prod_accum_106__3_,prod_accum_106__2_,prod_accum_106__1_,prod_accum_106__0_,
  prod_accum_105__106_,prod_accum_105__105_,prod_accum_105__104_,prod_accum_105__103_,
  prod_accum_105__102_,prod_accum_105__101_,prod_accum_105__100_,prod_accum_105__99_,
  prod_accum_105__98_,prod_accum_105__97_,prod_accum_105__96_,prod_accum_105__95_,
  prod_accum_105__94_,prod_accum_105__93_,prod_accum_105__92_,prod_accum_105__91_,
  prod_accum_105__90_,prod_accum_105__89_,prod_accum_105__88_,prod_accum_105__87_,
  prod_accum_105__86_,prod_accum_105__85_,prod_accum_105__84_,prod_accum_105__83_,
  prod_accum_105__82_,prod_accum_105__81_,prod_accum_105__80_,prod_accum_105__79_,
  prod_accum_105__78_,prod_accum_105__77_,prod_accum_105__76_,prod_accum_105__75_,
  prod_accum_105__74_,prod_accum_105__73_,prod_accum_105__72_,prod_accum_105__71_,
  prod_accum_105__70_,prod_accum_105__69_,prod_accum_105__68_,prod_accum_105__67_,
  prod_accum_105__66_,prod_accum_105__65_,prod_accum_105__64_,prod_accum_105__63_,
  prod_accum_105__62_,prod_accum_105__61_,prod_accum_105__60_,prod_accum_105__59_,
  prod_accum_105__58_,prod_accum_105__57_,prod_accum_105__56_,prod_accum_105__55_,
  prod_accum_105__54_,prod_accum_105__53_,prod_accum_105__52_,prod_accum_105__51_,
  prod_accum_105__50_,prod_accum_105__49_,prod_accum_105__48_,prod_accum_105__47_,
  prod_accum_105__46_,prod_accum_105__45_,prod_accum_105__44_,prod_accum_105__43_,
  prod_accum_105__42_,prod_accum_105__41_,prod_accum_105__40_,prod_accum_105__39_,
  prod_accum_105__38_,prod_accum_105__37_,prod_accum_105__36_,prod_accum_105__35_,
  prod_accum_105__34_,prod_accum_105__33_,prod_accum_105__32_,prod_accum_105__31_,
  prod_accum_105__30_,prod_accum_105__29_,prod_accum_105__28_,prod_accum_105__27_,
  prod_accum_105__26_,prod_accum_105__25_,prod_accum_105__24_,prod_accum_105__23_,
  prod_accum_105__22_,prod_accum_105__21_,prod_accum_105__20_,prod_accum_105__19_,
  prod_accum_105__18_,prod_accum_105__17_,prod_accum_105__16_,prod_accum_105__15_,
  prod_accum_105__14_,prod_accum_105__13_,prod_accum_105__12_,prod_accum_105__11_,
  prod_accum_105__10_,prod_accum_105__9_,prod_accum_105__8_,prod_accum_105__7_,
  prod_accum_105__6_,prod_accum_105__5_,prod_accum_105__4_,prod_accum_105__3_,
  prod_accum_105__2_,prod_accum_105__1_,prod_accum_105__0_,prod_accum_104__105_,
  prod_accum_104__104_,prod_accum_104__103_,prod_accum_104__102_,prod_accum_104__101_,
  prod_accum_104__100_,prod_accum_104__99_,prod_accum_104__98_,prod_accum_104__97_,
  prod_accum_104__96_,prod_accum_104__95_,prod_accum_104__94_,prod_accum_104__93_,
  prod_accum_104__92_,prod_accum_104__91_,prod_accum_104__90_,prod_accum_104__89_,
  prod_accum_104__88_,prod_accum_104__87_,prod_accum_104__86_,prod_accum_104__85_,
  prod_accum_104__84_,prod_accum_104__83_,prod_accum_104__82_,prod_accum_104__81_,
  prod_accum_104__80_,prod_accum_104__79_,prod_accum_104__78_,prod_accum_104__77_,
  prod_accum_104__76_,prod_accum_104__75_,prod_accum_104__74_,prod_accum_104__73_,
  prod_accum_104__72_,prod_accum_104__71_,prod_accum_104__70_,prod_accum_104__69_,
  prod_accum_104__68_,prod_accum_104__67_,prod_accum_104__66_,prod_accum_104__65_,
  prod_accum_104__64_,prod_accum_104__63_,prod_accum_104__62_,prod_accum_104__61_,
  prod_accum_104__60_,prod_accum_104__59_,prod_accum_104__58_,prod_accum_104__57_,
  prod_accum_104__56_,prod_accum_104__55_,prod_accum_104__54_,prod_accum_104__53_,
  prod_accum_104__52_,prod_accum_104__51_,prod_accum_104__50_,prod_accum_104__49_,
  prod_accum_104__48_,prod_accum_104__47_,prod_accum_104__46_,prod_accum_104__45_,
  prod_accum_104__44_,prod_accum_104__43_,prod_accum_104__42_,prod_accum_104__41_,
  prod_accum_104__40_,prod_accum_104__39_,prod_accum_104__38_,prod_accum_104__37_,
  prod_accum_104__36_,prod_accum_104__35_,prod_accum_104__34_,prod_accum_104__33_,
  prod_accum_104__32_,prod_accum_104__31_,prod_accum_104__30_,prod_accum_104__29_,
  prod_accum_104__28_,prod_accum_104__27_,prod_accum_104__26_,prod_accum_104__25_,
  prod_accum_104__24_,prod_accum_104__23_,prod_accum_104__22_,prod_accum_104__21_,
  prod_accum_104__20_,prod_accum_104__19_,prod_accum_104__18_,prod_accum_104__17_,
  prod_accum_104__16_,prod_accum_104__15_,prod_accum_104__14_,prod_accum_104__13_,
  prod_accum_104__12_,prod_accum_104__11_,prod_accum_104__10_,prod_accum_104__9_,
  prod_accum_104__8_,prod_accum_104__7_,prod_accum_104__6_,prod_accum_104__5_,
  prod_accum_104__4_,prod_accum_104__3_,prod_accum_104__2_,prod_accum_104__1_,
  prod_accum_104__0_,prod_accum_103__104_,prod_accum_103__103_,prod_accum_103__102_,
  prod_accum_103__101_,prod_accum_103__100_,prod_accum_103__99_,prod_accum_103__98_,
  prod_accum_103__97_,prod_accum_103__96_,prod_accum_103__95_,prod_accum_103__94_,
  prod_accum_103__93_,prod_accum_103__92_,prod_accum_103__91_,prod_accum_103__90_,
  prod_accum_103__89_,prod_accum_103__88_,prod_accum_103__87_,prod_accum_103__86_,
  prod_accum_103__85_,prod_accum_103__84_,prod_accum_103__83_,prod_accum_103__82_,
  prod_accum_103__81_,prod_accum_103__80_,prod_accum_103__79_,prod_accum_103__78_,
  prod_accum_103__77_,prod_accum_103__76_,prod_accum_103__75_,prod_accum_103__74_,
  prod_accum_103__73_,prod_accum_103__72_,prod_accum_103__71_,prod_accum_103__70_,
  prod_accum_103__69_,prod_accum_103__68_,prod_accum_103__67_,prod_accum_103__66_,
  prod_accum_103__65_,prod_accum_103__64_,prod_accum_103__63_,prod_accum_103__62_,
  prod_accum_103__61_,prod_accum_103__60_,prod_accum_103__59_,prod_accum_103__58_,
  prod_accum_103__57_,prod_accum_103__56_,prod_accum_103__55_,prod_accum_103__54_,
  prod_accum_103__53_,prod_accum_103__52_,prod_accum_103__51_,prod_accum_103__50_,
  prod_accum_103__49_,prod_accum_103__48_,prod_accum_103__47_,prod_accum_103__46_,
  prod_accum_103__45_,prod_accum_103__44_,prod_accum_103__43_,prod_accum_103__42_,
  prod_accum_103__41_,prod_accum_103__40_,prod_accum_103__39_,prod_accum_103__38_,
  prod_accum_103__37_,prod_accum_103__36_,prod_accum_103__35_,prod_accum_103__34_,
  prod_accum_103__33_,prod_accum_103__32_,prod_accum_103__31_,prod_accum_103__30_,
  prod_accum_103__29_,prod_accum_103__28_,prod_accum_103__27_,prod_accum_103__26_,
  prod_accum_103__25_,prod_accum_103__24_,prod_accum_103__23_,prod_accum_103__22_,
  prod_accum_103__21_,prod_accum_103__20_,prod_accum_103__19_,prod_accum_103__18_,
  prod_accum_103__17_,prod_accum_103__16_,prod_accum_103__15_,prod_accum_103__14_,
  prod_accum_103__13_,prod_accum_103__12_,prod_accum_103__11_,prod_accum_103__10_,
  prod_accum_103__9_,prod_accum_103__8_,prod_accum_103__7_,prod_accum_103__6_,
  prod_accum_103__5_,prod_accum_103__4_,prod_accum_103__3_,prod_accum_103__2_,
  prod_accum_103__1_,prod_accum_103__0_,s_r_110__127_,s_r_110__126_,s_r_110__125_,s_r_110__124_,
  s_r_110__123_,s_r_110__122_,s_r_110__121_,s_r_110__120_,s_r_110__119_,
  s_r_110__118_,s_r_110__117_,s_r_110__116_,s_r_110__115_,s_r_110__114_,s_r_110__113_,
  s_r_110__112_,s_r_110__111_,s_r_110__110_,s_r_110__109_,s_r_110__108_,s_r_110__107_,
  s_r_110__106_,s_r_110__105_,s_r_110__104_,s_r_110__103_,s_r_110__102_,s_r_110__101_,
  s_r_110__100_,s_r_110__99_,s_r_110__98_,s_r_110__97_,s_r_110__96_,s_r_110__95_,
  s_r_110__94_,s_r_110__93_,s_r_110__92_,s_r_110__91_,s_r_110__90_,s_r_110__89_,
  s_r_110__88_,s_r_110__87_,s_r_110__86_,s_r_110__85_,s_r_110__84_,s_r_110__83_,
  s_r_110__82_,s_r_110__81_,s_r_110__80_,s_r_110__79_,s_r_110__78_,s_r_110__77_,
  s_r_110__76_,s_r_110__75_,s_r_110__74_,s_r_110__73_,s_r_110__72_,s_r_110__71_,
  s_r_110__70_,s_r_110__69_,s_r_110__68_,s_r_110__67_,s_r_110__66_,s_r_110__65_,
  s_r_110__64_,s_r_110__63_,s_r_110__62_,s_r_110__61_,s_r_110__60_,s_r_110__59_,s_r_110__58_,
  s_r_110__57_,s_r_110__56_,s_r_110__55_,s_r_110__54_,s_r_110__53_,s_r_110__52_,
  s_r_110__51_,s_r_110__50_,s_r_110__49_,s_r_110__48_,s_r_110__47_,s_r_110__46_,
  s_r_110__45_,s_r_110__44_,s_r_110__43_,s_r_110__42_,s_r_110__41_,s_r_110__40_,
  s_r_110__39_,s_r_110__38_,s_r_110__37_,s_r_110__36_,s_r_110__35_,s_r_110__34_,
  s_r_110__33_,s_r_110__32_,s_r_110__31_,s_r_110__30_,s_r_110__29_,s_r_110__28_,
  s_r_110__27_,s_r_110__26_,s_r_110__25_,s_r_110__24_,s_r_110__23_,s_r_110__22_,s_r_110__21_,
  s_r_110__20_,s_r_110__19_,s_r_110__18_,s_r_110__17_,s_r_110__16_,s_r_110__15_,
  s_r_110__14_,s_r_110__13_,s_r_110__12_,s_r_110__11_,s_r_110__10_,s_r_110__9_,
  s_r_110__8_,s_r_110__7_,s_r_110__6_,s_r_110__5_,s_r_110__4_,s_r_110__3_,s_r_110__2_,
  s_r_110__1_,s_r_110__0_,s_r_109__127_,s_r_109__126_,s_r_109__125_,s_r_109__124_,
  s_r_109__123_,s_r_109__122_,s_r_109__121_,s_r_109__120_,s_r_109__119_,
  s_r_109__118_,s_r_109__117_,s_r_109__116_,s_r_109__115_,s_r_109__114_,s_r_109__113_,
  s_r_109__112_,s_r_109__111_,s_r_109__110_,s_r_109__109_,s_r_109__108_,s_r_109__107_,
  s_r_109__106_,s_r_109__105_,s_r_109__104_,s_r_109__103_,s_r_109__102_,
  s_r_109__101_,s_r_109__100_,s_r_109__99_,s_r_109__98_,s_r_109__97_,s_r_109__96_,s_r_109__95_,
  s_r_109__94_,s_r_109__93_,s_r_109__92_,s_r_109__91_,s_r_109__90_,s_r_109__89_,
  s_r_109__88_,s_r_109__87_,s_r_109__86_,s_r_109__85_,s_r_109__84_,s_r_109__83_,
  s_r_109__82_,s_r_109__81_,s_r_109__80_,s_r_109__79_,s_r_109__78_,s_r_109__77_,
  s_r_109__76_,s_r_109__75_,s_r_109__74_,s_r_109__73_,s_r_109__72_,s_r_109__71_,
  s_r_109__70_,s_r_109__69_,s_r_109__68_,s_r_109__67_,s_r_109__66_,s_r_109__65_,
  s_r_109__64_,s_r_109__63_,s_r_109__62_,s_r_109__61_,s_r_109__60_,s_r_109__59_,
  s_r_109__58_,s_r_109__57_,s_r_109__56_,s_r_109__55_,s_r_109__54_,s_r_109__53_,s_r_109__52_,
  s_r_109__51_,s_r_109__50_,s_r_109__49_,s_r_109__48_,s_r_109__47_,s_r_109__46_,
  s_r_109__45_,s_r_109__44_,s_r_109__43_,s_r_109__42_,s_r_109__41_,s_r_109__40_,
  s_r_109__39_,s_r_109__38_,s_r_109__37_,s_r_109__36_,s_r_109__35_,s_r_109__34_,
  s_r_109__33_,s_r_109__32_,s_r_109__31_,s_r_109__30_,s_r_109__29_,s_r_109__28_,
  s_r_109__27_,s_r_109__26_,s_r_109__25_,s_r_109__24_,s_r_109__23_,s_r_109__22_,
  s_r_109__21_,s_r_109__20_,s_r_109__19_,s_r_109__18_,s_r_109__17_,s_r_109__16_,s_r_109__15_,
  s_r_109__14_,s_r_109__13_,s_r_109__12_,s_r_109__11_,s_r_109__10_,s_r_109__9_,
  s_r_109__8_,s_r_109__7_,s_r_109__6_,s_r_109__5_,s_r_109__4_,s_r_109__3_,
  s_r_109__2_,s_r_109__1_,s_r_109__0_,s_r_108__127_,s_r_108__126_,s_r_108__125_,
  s_r_108__124_,s_r_108__123_,s_r_108__122_,s_r_108__121_,s_r_108__120_,s_r_108__119_,
  s_r_108__118_,s_r_108__117_,s_r_108__116_,s_r_108__115_,s_r_108__114_,s_r_108__113_,
  s_r_108__112_,s_r_108__111_,s_r_108__110_,s_r_108__109_,s_r_108__108_,s_r_108__107_,
  s_r_108__106_,s_r_108__105_,s_r_108__104_,s_r_108__103_,s_r_108__102_,
  s_r_108__101_,s_r_108__100_,s_r_108__99_,s_r_108__98_,s_r_108__97_,s_r_108__96_,
  s_r_108__95_,s_r_108__94_,s_r_108__93_,s_r_108__92_,s_r_108__91_,s_r_108__90_,s_r_108__89_,
  s_r_108__88_,s_r_108__87_,s_r_108__86_,s_r_108__85_,s_r_108__84_,s_r_108__83_,
  s_r_108__82_,s_r_108__81_,s_r_108__80_,s_r_108__79_,s_r_108__78_,s_r_108__77_,
  s_r_108__76_,s_r_108__75_,s_r_108__74_,s_r_108__73_,s_r_108__72_,s_r_108__71_,
  s_r_108__70_,s_r_108__69_,s_r_108__68_,s_r_108__67_,s_r_108__66_,s_r_108__65_,
  s_r_108__64_,s_r_108__63_,s_r_108__62_,s_r_108__61_,s_r_108__60_,s_r_108__59_,
  s_r_108__58_,s_r_108__57_,s_r_108__56_,s_r_108__55_,s_r_108__54_,s_r_108__53_,
  s_r_108__52_,s_r_108__51_,s_r_108__50_,s_r_108__49_,s_r_108__48_,s_r_108__47_,s_r_108__46_,
  s_r_108__45_,s_r_108__44_,s_r_108__43_,s_r_108__42_,s_r_108__41_,s_r_108__40_,
  s_r_108__39_,s_r_108__38_,s_r_108__37_,s_r_108__36_,s_r_108__35_,s_r_108__34_,
  s_r_108__33_,s_r_108__32_,s_r_108__31_,s_r_108__30_,s_r_108__29_,s_r_108__28_,
  s_r_108__27_,s_r_108__26_,s_r_108__25_,s_r_108__24_,s_r_108__23_,s_r_108__22_,
  s_r_108__21_,s_r_108__20_,s_r_108__19_,s_r_108__18_,s_r_108__17_,s_r_108__16_,
  s_r_108__15_,s_r_108__14_,s_r_108__13_,s_r_108__12_,s_r_108__11_,s_r_108__10_,s_r_108__9_,
  s_r_108__8_,s_r_108__7_,s_r_108__6_,s_r_108__5_,s_r_108__4_,s_r_108__3_,
  s_r_108__2_,s_r_108__1_,s_r_108__0_,s_r_107__127_,s_r_107__126_,s_r_107__125_,
  s_r_107__124_,s_r_107__123_,s_r_107__122_,s_r_107__121_,s_r_107__120_,s_r_107__119_,
  s_r_107__118_,s_r_107__117_,s_r_107__116_,s_r_107__115_,s_r_107__114_,s_r_107__113_,
  s_r_107__112_,s_r_107__111_,s_r_107__110_,s_r_107__109_,s_r_107__108_,
  s_r_107__107_,s_r_107__106_,s_r_107__105_,s_r_107__104_,s_r_107__103_,s_r_107__102_,
  s_r_107__101_,s_r_107__100_,s_r_107__99_,s_r_107__98_,s_r_107__97_,s_r_107__96_,
  s_r_107__95_,s_r_107__94_,s_r_107__93_,s_r_107__92_,s_r_107__91_,s_r_107__90_,
  s_r_107__89_,s_r_107__88_,s_r_107__87_,s_r_107__86_,s_r_107__85_,s_r_107__84_,s_r_107__83_,
  s_r_107__82_,s_r_107__81_,s_r_107__80_,s_r_107__79_,s_r_107__78_,s_r_107__77_,
  s_r_107__76_,s_r_107__75_,s_r_107__74_,s_r_107__73_,s_r_107__72_,s_r_107__71_,
  s_r_107__70_,s_r_107__69_,s_r_107__68_,s_r_107__67_,s_r_107__66_,s_r_107__65_,
  s_r_107__64_,s_r_107__63_,s_r_107__62_,s_r_107__61_,s_r_107__60_,s_r_107__59_,
  s_r_107__58_,s_r_107__57_,s_r_107__56_,s_r_107__55_,s_r_107__54_,s_r_107__53_,
  s_r_107__52_,s_r_107__51_,s_r_107__50_,s_r_107__49_,s_r_107__48_,s_r_107__47_,
  s_r_107__46_,s_r_107__45_,s_r_107__44_,s_r_107__43_,s_r_107__42_,s_r_107__41_,s_r_107__40_,
  s_r_107__39_,s_r_107__38_,s_r_107__37_,s_r_107__36_,s_r_107__35_,s_r_107__34_,
  s_r_107__33_,s_r_107__32_,s_r_107__31_,s_r_107__30_,s_r_107__29_,s_r_107__28_,
  s_r_107__27_,s_r_107__26_,s_r_107__25_,s_r_107__24_,s_r_107__23_,s_r_107__22_,
  s_r_107__21_,s_r_107__20_,s_r_107__19_,s_r_107__18_,s_r_107__17_,s_r_107__16_,
  s_r_107__15_,s_r_107__14_,s_r_107__13_,s_r_107__12_,s_r_107__11_,s_r_107__10_,
  s_r_107__9_,s_r_107__8_,s_r_107__7_,s_r_107__6_,s_r_107__5_,s_r_107__4_,s_r_107__3_,
  s_r_107__2_,s_r_107__1_,s_r_107__0_,prod_accum_110__111_,prod_accum_110__110_,
  prod_accum_110__109_,prod_accum_110__108_,prod_accum_110__107_,prod_accum_110__106_,
  prod_accum_110__105_,prod_accum_110__104_,prod_accum_110__103_,prod_accum_110__102_,
  prod_accum_110__101_,prod_accum_110__100_,prod_accum_110__99_,
  prod_accum_110__98_,prod_accum_110__97_,prod_accum_110__96_,prod_accum_110__95_,
  prod_accum_110__94_,prod_accum_110__93_,prod_accum_110__92_,prod_accum_110__91_,
  prod_accum_110__90_,prod_accum_110__89_,prod_accum_110__88_,prod_accum_110__87_,
  prod_accum_110__86_,prod_accum_110__85_,prod_accum_110__84_,prod_accum_110__83_,
  prod_accum_110__82_,prod_accum_110__81_,prod_accum_110__80_,prod_accum_110__79_,
  prod_accum_110__78_,prod_accum_110__77_,prod_accum_110__76_,prod_accum_110__75_,
  prod_accum_110__74_,prod_accum_110__73_,prod_accum_110__72_,prod_accum_110__71_,
  prod_accum_110__70_,prod_accum_110__69_,prod_accum_110__68_,prod_accum_110__67_,
  prod_accum_110__66_,prod_accum_110__65_,prod_accum_110__64_,prod_accum_110__63_,
  prod_accum_110__62_,prod_accum_110__61_,prod_accum_110__60_,prod_accum_110__59_,
  prod_accum_110__58_,prod_accum_110__57_,prod_accum_110__56_,prod_accum_110__55_,
  prod_accum_110__54_,prod_accum_110__53_,prod_accum_110__52_,prod_accum_110__51_,
  prod_accum_110__50_,prod_accum_110__49_,prod_accum_110__48_,prod_accum_110__47_,
  prod_accum_110__46_,prod_accum_110__45_,prod_accum_110__44_,prod_accum_110__43_,
  prod_accum_110__42_,prod_accum_110__41_,prod_accum_110__40_,prod_accum_110__39_,
  prod_accum_110__38_,prod_accum_110__37_,prod_accum_110__36_,prod_accum_110__35_,
  prod_accum_110__34_,prod_accum_110__33_,prod_accum_110__32_,prod_accum_110__31_,
  prod_accum_110__30_,prod_accum_110__29_,prod_accum_110__28_,prod_accum_110__27_,
  prod_accum_110__26_,prod_accum_110__25_,prod_accum_110__24_,prod_accum_110__23_,
  prod_accum_110__22_,prod_accum_110__21_,prod_accum_110__20_,prod_accum_110__19_,
  prod_accum_110__18_,prod_accum_110__17_,prod_accum_110__16_,prod_accum_110__15_,
  prod_accum_110__14_,prod_accum_110__13_,prod_accum_110__12_,prod_accum_110__11_,
  prod_accum_110__10_,prod_accum_110__9_,prod_accum_110__8_,prod_accum_110__7_,prod_accum_110__6_,
  prod_accum_110__5_,prod_accum_110__4_,prod_accum_110__3_,prod_accum_110__2_,
  prod_accum_110__1_,prod_accum_110__0_,prod_accum_109__110_,prod_accum_109__109_,
  prod_accum_109__108_,prod_accum_109__107_,prod_accum_109__106_,prod_accum_109__105_,
  prod_accum_109__104_,prod_accum_109__103_,prod_accum_109__102_,
  prod_accum_109__101_,prod_accum_109__100_,prod_accum_109__99_,prod_accum_109__98_,
  prod_accum_109__97_,prod_accum_109__96_,prod_accum_109__95_,prod_accum_109__94_,
  prod_accum_109__93_,prod_accum_109__92_,prod_accum_109__91_,prod_accum_109__90_,
  prod_accum_109__89_,prod_accum_109__88_,prod_accum_109__87_,prod_accum_109__86_,
  prod_accum_109__85_,prod_accum_109__84_,prod_accum_109__83_,prod_accum_109__82_,
  prod_accum_109__81_,prod_accum_109__80_,prod_accum_109__79_,prod_accum_109__78_,
  prod_accum_109__77_,prod_accum_109__76_,prod_accum_109__75_,prod_accum_109__74_,
  prod_accum_109__73_,prod_accum_109__72_,prod_accum_109__71_,prod_accum_109__70_,
  prod_accum_109__69_,prod_accum_109__68_,prod_accum_109__67_,prod_accum_109__66_,
  prod_accum_109__65_,prod_accum_109__64_,prod_accum_109__63_,prod_accum_109__62_,
  prod_accum_109__61_,prod_accum_109__60_,prod_accum_109__59_,prod_accum_109__58_,
  prod_accum_109__57_,prod_accum_109__56_,prod_accum_109__55_,prod_accum_109__54_,
  prod_accum_109__53_,prod_accum_109__52_,prod_accum_109__51_,prod_accum_109__50_,
  prod_accum_109__49_,prod_accum_109__48_,prod_accum_109__47_,prod_accum_109__46_,
  prod_accum_109__45_,prod_accum_109__44_,prod_accum_109__43_,prod_accum_109__42_,
  prod_accum_109__41_,prod_accum_109__40_,prod_accum_109__39_,prod_accum_109__38_,
  prod_accum_109__37_,prod_accum_109__36_,prod_accum_109__35_,prod_accum_109__34_,
  prod_accum_109__33_,prod_accum_109__32_,prod_accum_109__31_,prod_accum_109__30_,
  prod_accum_109__29_,prod_accum_109__28_,prod_accum_109__27_,prod_accum_109__26_,
  prod_accum_109__25_,prod_accum_109__24_,prod_accum_109__23_,prod_accum_109__22_,
  prod_accum_109__21_,prod_accum_109__20_,prod_accum_109__19_,prod_accum_109__18_,
  prod_accum_109__17_,prod_accum_109__16_,prod_accum_109__15_,prod_accum_109__14_,
  prod_accum_109__13_,prod_accum_109__12_,prod_accum_109__11_,prod_accum_109__10_,
  prod_accum_109__9_,prod_accum_109__8_,prod_accum_109__7_,prod_accum_109__6_,prod_accum_109__5_,
  prod_accum_109__4_,prod_accum_109__3_,prod_accum_109__2_,prod_accum_109__1_,
  prod_accum_109__0_,prod_accum_108__109_,prod_accum_108__108_,prod_accum_108__107_,
  prod_accum_108__106_,prod_accum_108__105_,prod_accum_108__104_,prod_accum_108__103_,
  prod_accum_108__102_,prod_accum_108__101_,prod_accum_108__100_,
  prod_accum_108__99_,prod_accum_108__98_,prod_accum_108__97_,prod_accum_108__96_,
  prod_accum_108__95_,prod_accum_108__94_,prod_accum_108__93_,prod_accum_108__92_,
  prod_accum_108__91_,prod_accum_108__90_,prod_accum_108__89_,prod_accum_108__88_,
  prod_accum_108__87_,prod_accum_108__86_,prod_accum_108__85_,prod_accum_108__84_,
  prod_accum_108__83_,prod_accum_108__82_,prod_accum_108__81_,prod_accum_108__80_,
  prod_accum_108__79_,prod_accum_108__78_,prod_accum_108__77_,prod_accum_108__76_,
  prod_accum_108__75_,prod_accum_108__74_,prod_accum_108__73_,prod_accum_108__72_,
  prod_accum_108__71_,prod_accum_108__70_,prod_accum_108__69_,prod_accum_108__68_,
  prod_accum_108__67_,prod_accum_108__66_,prod_accum_108__65_,prod_accum_108__64_,
  prod_accum_108__63_,prod_accum_108__62_,prod_accum_108__61_,prod_accum_108__60_,
  prod_accum_108__59_,prod_accum_108__58_,prod_accum_108__57_,prod_accum_108__56_,
  prod_accum_108__55_,prod_accum_108__54_,prod_accum_108__53_,prod_accum_108__52_,
  prod_accum_108__51_,prod_accum_108__50_,prod_accum_108__49_,prod_accum_108__48_,
  prod_accum_108__47_,prod_accum_108__46_,prod_accum_108__45_,prod_accum_108__44_,
  prod_accum_108__43_,prod_accum_108__42_,prod_accum_108__41_,prod_accum_108__40_,
  prod_accum_108__39_,prod_accum_108__38_,prod_accum_108__37_,prod_accum_108__36_,
  prod_accum_108__35_,prod_accum_108__34_,prod_accum_108__33_,prod_accum_108__32_,
  prod_accum_108__31_,prod_accum_108__30_,prod_accum_108__29_,prod_accum_108__28_,
  prod_accum_108__27_,prod_accum_108__26_,prod_accum_108__25_,prod_accum_108__24_,
  prod_accum_108__23_,prod_accum_108__22_,prod_accum_108__21_,prod_accum_108__20_,
  prod_accum_108__19_,prod_accum_108__18_,prod_accum_108__17_,prod_accum_108__16_,
  prod_accum_108__15_,prod_accum_108__14_,prod_accum_108__13_,prod_accum_108__12_,
  prod_accum_108__11_,prod_accum_108__10_,prod_accum_108__9_,prod_accum_108__8_,prod_accum_108__7_,
  prod_accum_108__6_,prod_accum_108__5_,prod_accum_108__4_,prod_accum_108__3_,
  prod_accum_108__2_,prod_accum_108__1_,prod_accum_108__0_,prod_accum_107__108_,
  prod_accum_107__107_,prod_accum_107__106_,prod_accum_107__105_,prod_accum_107__104_,
  prod_accum_107__103_,prod_accum_107__102_,prod_accum_107__101_,
  prod_accum_107__100_,prod_accum_107__99_,prod_accum_107__98_,prod_accum_107__97_,
  prod_accum_107__96_,prod_accum_107__95_,prod_accum_107__94_,prod_accum_107__93_,
  prod_accum_107__92_,prod_accum_107__91_,prod_accum_107__90_,prod_accum_107__89_,
  prod_accum_107__88_,prod_accum_107__87_,prod_accum_107__86_,prod_accum_107__85_,
  prod_accum_107__84_,prod_accum_107__83_,prod_accum_107__82_,prod_accum_107__81_,
  prod_accum_107__80_,prod_accum_107__79_,prod_accum_107__78_,prod_accum_107__77_,
  prod_accum_107__76_,prod_accum_107__75_,prod_accum_107__74_,prod_accum_107__73_,
  prod_accum_107__72_,prod_accum_107__71_,prod_accum_107__70_,prod_accum_107__69_,
  prod_accum_107__68_,prod_accum_107__67_,prod_accum_107__66_,prod_accum_107__65_,
  prod_accum_107__64_,prod_accum_107__63_,prod_accum_107__62_,prod_accum_107__61_,
  prod_accum_107__60_,prod_accum_107__59_,prod_accum_107__58_,prod_accum_107__57_,
  prod_accum_107__56_,prod_accum_107__55_,prod_accum_107__54_,prod_accum_107__53_,
  prod_accum_107__52_,prod_accum_107__51_,prod_accum_107__50_,prod_accum_107__49_,
  prod_accum_107__48_,prod_accum_107__47_,prod_accum_107__46_,prod_accum_107__45_,
  prod_accum_107__44_,prod_accum_107__43_,prod_accum_107__42_,prod_accum_107__41_,
  prod_accum_107__40_,prod_accum_107__39_,prod_accum_107__38_,prod_accum_107__37_,
  prod_accum_107__36_,prod_accum_107__35_,prod_accum_107__34_,prod_accum_107__33_,
  prod_accum_107__32_,prod_accum_107__31_,prod_accum_107__30_,prod_accum_107__29_,
  prod_accum_107__28_,prod_accum_107__27_,prod_accum_107__26_,prod_accum_107__25_,
  prod_accum_107__24_,prod_accum_107__23_,prod_accum_107__22_,prod_accum_107__21_,
  prod_accum_107__20_,prod_accum_107__19_,prod_accum_107__18_,prod_accum_107__17_,
  prod_accum_107__16_,prod_accum_107__15_,prod_accum_107__14_,prod_accum_107__13_,
  prod_accum_107__12_,prod_accum_107__11_,prod_accum_107__10_,prod_accum_107__9_,prod_accum_107__8_,
  prod_accum_107__7_,prod_accum_107__6_,prod_accum_107__5_,prod_accum_107__4_,
  prod_accum_107__3_,prod_accum_107__2_,prod_accum_107__1_,prod_accum_107__0_,
  s_r_114__127_,s_r_114__126_,s_r_114__125_,s_r_114__124_,s_r_114__123_,s_r_114__122_,
  s_r_114__121_,s_r_114__120_,s_r_114__119_,s_r_114__118_,s_r_114__117_,s_r_114__116_,
  s_r_114__115_,s_r_114__114_,s_r_114__113_,s_r_114__112_,s_r_114__111_,
  s_r_114__110_,s_r_114__109_,s_r_114__108_,s_r_114__107_,s_r_114__106_,s_r_114__105_,
  s_r_114__104_,s_r_114__103_,s_r_114__102_,s_r_114__101_,s_r_114__100_,s_r_114__99_,
  s_r_114__98_,s_r_114__97_,s_r_114__96_,s_r_114__95_,s_r_114__94_,s_r_114__93_,
  s_r_114__92_,s_r_114__91_,s_r_114__90_,s_r_114__89_,s_r_114__88_,s_r_114__87_,
  s_r_114__86_,s_r_114__85_,s_r_114__84_,s_r_114__83_,s_r_114__82_,s_r_114__81_,
  s_r_114__80_,s_r_114__79_,s_r_114__78_,s_r_114__77_,s_r_114__76_,s_r_114__75_,
  s_r_114__74_,s_r_114__73_,s_r_114__72_,s_r_114__71_,s_r_114__70_,s_r_114__69_,s_r_114__68_,
  s_r_114__67_,s_r_114__66_,s_r_114__65_,s_r_114__64_,s_r_114__63_,s_r_114__62_,
  s_r_114__61_,s_r_114__60_,s_r_114__59_,s_r_114__58_,s_r_114__57_,s_r_114__56_,
  s_r_114__55_,s_r_114__54_,s_r_114__53_,s_r_114__52_,s_r_114__51_,s_r_114__50_,
  s_r_114__49_,s_r_114__48_,s_r_114__47_,s_r_114__46_,s_r_114__45_,s_r_114__44_,
  s_r_114__43_,s_r_114__42_,s_r_114__41_,s_r_114__40_,s_r_114__39_,s_r_114__38_,
  s_r_114__37_,s_r_114__36_,s_r_114__35_,s_r_114__34_,s_r_114__33_,s_r_114__32_,s_r_114__31_,
  s_r_114__30_,s_r_114__29_,s_r_114__28_,s_r_114__27_,s_r_114__26_,s_r_114__25_,
  s_r_114__24_,s_r_114__23_,s_r_114__22_,s_r_114__21_,s_r_114__20_,s_r_114__19_,
  s_r_114__18_,s_r_114__17_,s_r_114__16_,s_r_114__15_,s_r_114__14_,s_r_114__13_,
  s_r_114__12_,s_r_114__11_,s_r_114__10_,s_r_114__9_,s_r_114__8_,s_r_114__7_,
  s_r_114__6_,s_r_114__5_,s_r_114__4_,s_r_114__3_,s_r_114__2_,s_r_114__1_,s_r_114__0_,
  s_r_113__127_,s_r_113__126_,s_r_113__125_,s_r_113__124_,s_r_113__123_,s_r_113__122_,
  s_r_113__121_,s_r_113__120_,s_r_113__119_,s_r_113__118_,s_r_113__117_,
  s_r_113__116_,s_r_113__115_,s_r_113__114_,s_r_113__113_,s_r_113__112_,s_r_113__111_,
  s_r_113__110_,s_r_113__109_,s_r_113__108_,s_r_113__107_,s_r_113__106_,s_r_113__105_,
  s_r_113__104_,s_r_113__103_,s_r_113__102_,s_r_113__101_,s_r_113__100_,s_r_113__99_,
  s_r_113__98_,s_r_113__97_,s_r_113__96_,s_r_113__95_,s_r_113__94_,s_r_113__93_,
  s_r_113__92_,s_r_113__91_,s_r_113__90_,s_r_113__89_,s_r_113__88_,s_r_113__87_,
  s_r_113__86_,s_r_113__85_,s_r_113__84_,s_r_113__83_,s_r_113__82_,s_r_113__81_,
  s_r_113__80_,s_r_113__79_,s_r_113__78_,s_r_113__77_,s_r_113__76_,s_r_113__75_,
  s_r_113__74_,s_r_113__73_,s_r_113__72_,s_r_113__71_,s_r_113__70_,s_r_113__69_,
  s_r_113__68_,s_r_113__67_,s_r_113__66_,s_r_113__65_,s_r_113__64_,s_r_113__63_,s_r_113__62_,
  s_r_113__61_,s_r_113__60_,s_r_113__59_,s_r_113__58_,s_r_113__57_,s_r_113__56_,
  s_r_113__55_,s_r_113__54_,s_r_113__53_,s_r_113__52_,s_r_113__51_,s_r_113__50_,
  s_r_113__49_,s_r_113__48_,s_r_113__47_,s_r_113__46_,s_r_113__45_,s_r_113__44_,
  s_r_113__43_,s_r_113__42_,s_r_113__41_,s_r_113__40_,s_r_113__39_,s_r_113__38_,
  s_r_113__37_,s_r_113__36_,s_r_113__35_,s_r_113__34_,s_r_113__33_,s_r_113__32_,
  s_r_113__31_,s_r_113__30_,s_r_113__29_,s_r_113__28_,s_r_113__27_,s_r_113__26_,s_r_113__25_,
  s_r_113__24_,s_r_113__23_,s_r_113__22_,s_r_113__21_,s_r_113__20_,s_r_113__19_,
  s_r_113__18_,s_r_113__17_,s_r_113__16_,s_r_113__15_,s_r_113__14_,s_r_113__13_,
  s_r_113__12_,s_r_113__11_,s_r_113__10_,s_r_113__9_,s_r_113__8_,s_r_113__7_,
  s_r_113__6_,s_r_113__5_,s_r_113__4_,s_r_113__3_,s_r_113__2_,s_r_113__1_,s_r_113__0_,
  s_r_112__127_,s_r_112__126_,s_r_112__125_,s_r_112__124_,s_r_112__123_,s_r_112__122_,
  s_r_112__121_,s_r_112__120_,s_r_112__119_,s_r_112__118_,s_r_112__117_,
  s_r_112__116_,s_r_112__115_,s_r_112__114_,s_r_112__113_,s_r_112__112_,s_r_112__111_,
  s_r_112__110_,s_r_112__109_,s_r_112__108_,s_r_112__107_,s_r_112__106_,s_r_112__105_,
  s_r_112__104_,s_r_112__103_,s_r_112__102_,s_r_112__101_,s_r_112__100_,s_r_112__99_,
  s_r_112__98_,s_r_112__97_,s_r_112__96_,s_r_112__95_,s_r_112__94_,s_r_112__93_,
  s_r_112__92_,s_r_112__91_,s_r_112__90_,s_r_112__89_,s_r_112__88_,s_r_112__87_,
  s_r_112__86_,s_r_112__85_,s_r_112__84_,s_r_112__83_,s_r_112__82_,s_r_112__81_,
  s_r_112__80_,s_r_112__79_,s_r_112__78_,s_r_112__77_,s_r_112__76_,s_r_112__75_,
  s_r_112__74_,s_r_112__73_,s_r_112__72_,s_r_112__71_,s_r_112__70_,s_r_112__69_,
  s_r_112__68_,s_r_112__67_,s_r_112__66_,s_r_112__65_,s_r_112__64_,s_r_112__63_,
  s_r_112__62_,s_r_112__61_,s_r_112__60_,s_r_112__59_,s_r_112__58_,s_r_112__57_,s_r_112__56_,
  s_r_112__55_,s_r_112__54_,s_r_112__53_,s_r_112__52_,s_r_112__51_,s_r_112__50_,
  s_r_112__49_,s_r_112__48_,s_r_112__47_,s_r_112__46_,s_r_112__45_,s_r_112__44_,
  s_r_112__43_,s_r_112__42_,s_r_112__41_,s_r_112__40_,s_r_112__39_,s_r_112__38_,
  s_r_112__37_,s_r_112__36_,s_r_112__35_,s_r_112__34_,s_r_112__33_,s_r_112__32_,
  s_r_112__31_,s_r_112__30_,s_r_112__29_,s_r_112__28_,s_r_112__27_,s_r_112__26_,
  s_r_112__25_,s_r_112__24_,s_r_112__23_,s_r_112__22_,s_r_112__21_,s_r_112__20_,s_r_112__19_,
  s_r_112__18_,s_r_112__17_,s_r_112__16_,s_r_112__15_,s_r_112__14_,s_r_112__13_,
  s_r_112__12_,s_r_112__11_,s_r_112__10_,s_r_112__9_,s_r_112__8_,s_r_112__7_,
  s_r_112__6_,s_r_112__5_,s_r_112__4_,s_r_112__3_,s_r_112__2_,s_r_112__1_,s_r_112__0_,
  s_r_111__127_,s_r_111__126_,s_r_111__125_,s_r_111__124_,s_r_111__123_,
  s_r_111__122_,s_r_111__121_,s_r_111__120_,s_r_111__119_,s_r_111__118_,s_r_111__117_,
  s_r_111__116_,s_r_111__115_,s_r_111__114_,s_r_111__113_,s_r_111__112_,s_r_111__111_,
  s_r_111__110_,s_r_111__109_,s_r_111__108_,s_r_111__107_,s_r_111__106_,s_r_111__105_,
  s_r_111__104_,s_r_111__103_,s_r_111__102_,s_r_111__101_,s_r_111__100_,
  s_r_111__99_,s_r_111__98_,s_r_111__97_,s_r_111__96_,s_r_111__95_,s_r_111__94_,s_r_111__93_,
  s_r_111__92_,s_r_111__91_,s_r_111__90_,s_r_111__89_,s_r_111__88_,s_r_111__87_,
  s_r_111__86_,s_r_111__85_,s_r_111__84_,s_r_111__83_,s_r_111__82_,s_r_111__81_,
  s_r_111__80_,s_r_111__79_,s_r_111__78_,s_r_111__77_,s_r_111__76_,s_r_111__75_,
  s_r_111__74_,s_r_111__73_,s_r_111__72_,s_r_111__71_,s_r_111__70_,s_r_111__69_,
  s_r_111__68_,s_r_111__67_,s_r_111__66_,s_r_111__65_,s_r_111__64_,s_r_111__63_,
  s_r_111__62_,s_r_111__61_,s_r_111__60_,s_r_111__59_,s_r_111__58_,s_r_111__57_,
  s_r_111__56_,s_r_111__55_,s_r_111__54_,s_r_111__53_,s_r_111__52_,s_r_111__51_,s_r_111__50_,
  s_r_111__49_,s_r_111__48_,s_r_111__47_,s_r_111__46_,s_r_111__45_,s_r_111__44_,
  s_r_111__43_,s_r_111__42_,s_r_111__41_,s_r_111__40_,s_r_111__39_,s_r_111__38_,
  s_r_111__37_,s_r_111__36_,s_r_111__35_,s_r_111__34_,s_r_111__33_,s_r_111__32_,
  s_r_111__31_,s_r_111__30_,s_r_111__29_,s_r_111__28_,s_r_111__27_,s_r_111__26_,
  s_r_111__25_,s_r_111__24_,s_r_111__23_,s_r_111__22_,s_r_111__21_,s_r_111__20_,
  s_r_111__19_,s_r_111__18_,s_r_111__17_,s_r_111__16_,s_r_111__15_,s_r_111__14_,s_r_111__13_,
  s_r_111__12_,s_r_111__11_,s_r_111__10_,s_r_111__9_,s_r_111__8_,s_r_111__7_,
  s_r_111__6_,s_r_111__5_,s_r_111__4_,s_r_111__3_,s_r_111__2_,s_r_111__1_,s_r_111__0_,
  prod_accum_114__115_,prod_accum_114__114_,prod_accum_114__113_,
  prod_accum_114__112_,prod_accum_114__111_,prod_accum_114__110_,prod_accum_114__109_,
  prod_accum_114__108_,prod_accum_114__107_,prod_accum_114__106_,prod_accum_114__105_,
  prod_accum_114__104_,prod_accum_114__103_,prod_accum_114__102_,prod_accum_114__101_,
  prod_accum_114__100_,prod_accum_114__99_,prod_accum_114__98_,prod_accum_114__97_,
  prod_accum_114__96_,prod_accum_114__95_,prod_accum_114__94_,prod_accum_114__93_,
  prod_accum_114__92_,prod_accum_114__91_,prod_accum_114__90_,prod_accum_114__89_,
  prod_accum_114__88_,prod_accum_114__87_,prod_accum_114__86_,prod_accum_114__85_,
  prod_accum_114__84_,prod_accum_114__83_,prod_accum_114__82_,prod_accum_114__81_,
  prod_accum_114__80_,prod_accum_114__79_,prod_accum_114__78_,prod_accum_114__77_,
  prod_accum_114__76_,prod_accum_114__75_,prod_accum_114__74_,prod_accum_114__73_,
  prod_accum_114__72_,prod_accum_114__71_,prod_accum_114__70_,prod_accum_114__69_,
  prod_accum_114__68_,prod_accum_114__67_,prod_accum_114__66_,prod_accum_114__65_,
  prod_accum_114__64_,prod_accum_114__63_,prod_accum_114__62_,prod_accum_114__61_,
  prod_accum_114__60_,prod_accum_114__59_,prod_accum_114__58_,prod_accum_114__57_,
  prod_accum_114__56_,prod_accum_114__55_,prod_accum_114__54_,prod_accum_114__53_,
  prod_accum_114__52_,prod_accum_114__51_,prod_accum_114__50_,prod_accum_114__49_,
  prod_accum_114__48_,prod_accum_114__47_,prod_accum_114__46_,prod_accum_114__45_,
  prod_accum_114__44_,prod_accum_114__43_,prod_accum_114__42_,prod_accum_114__41_,
  prod_accum_114__40_,prod_accum_114__39_,prod_accum_114__38_,prod_accum_114__37_,
  prod_accum_114__36_,prod_accum_114__35_,prod_accum_114__34_,prod_accum_114__33_,
  prod_accum_114__32_,prod_accum_114__31_,prod_accum_114__30_,prod_accum_114__29_,
  prod_accum_114__28_,prod_accum_114__27_,prod_accum_114__26_,prod_accum_114__25_,
  prod_accum_114__24_,prod_accum_114__23_,prod_accum_114__22_,prod_accum_114__21_,
  prod_accum_114__20_,prod_accum_114__19_,prod_accum_114__18_,prod_accum_114__17_,
  prod_accum_114__16_,prod_accum_114__15_,prod_accum_114__14_,prod_accum_114__13_,
  prod_accum_114__12_,prod_accum_114__11_,prod_accum_114__10_,prod_accum_114__9_,
  prod_accum_114__8_,prod_accum_114__7_,prod_accum_114__6_,prod_accum_114__5_,
  prod_accum_114__4_,prod_accum_114__3_,prod_accum_114__2_,prod_accum_114__1_,
  prod_accum_114__0_,prod_accum_113__114_,prod_accum_113__113_,prod_accum_113__112_,
  prod_accum_113__111_,prod_accum_113__110_,prod_accum_113__109_,prod_accum_113__108_,
  prod_accum_113__107_,prod_accum_113__106_,prod_accum_113__105_,prod_accum_113__104_,
  prod_accum_113__103_,prod_accum_113__102_,prod_accum_113__101_,prod_accum_113__100_,
  prod_accum_113__99_,prod_accum_113__98_,prod_accum_113__97_,prod_accum_113__96_,
  prod_accum_113__95_,prod_accum_113__94_,prod_accum_113__93_,prod_accum_113__92_,
  prod_accum_113__91_,prod_accum_113__90_,prod_accum_113__89_,prod_accum_113__88_,
  prod_accum_113__87_,prod_accum_113__86_,prod_accum_113__85_,prod_accum_113__84_,
  prod_accum_113__83_,prod_accum_113__82_,prod_accum_113__81_,prod_accum_113__80_,
  prod_accum_113__79_,prod_accum_113__78_,prod_accum_113__77_,prod_accum_113__76_,
  prod_accum_113__75_,prod_accum_113__74_,prod_accum_113__73_,prod_accum_113__72_,
  prod_accum_113__71_,prod_accum_113__70_,prod_accum_113__69_,prod_accum_113__68_,
  prod_accum_113__67_,prod_accum_113__66_,prod_accum_113__65_,prod_accum_113__64_,
  prod_accum_113__63_,prod_accum_113__62_,prod_accum_113__61_,prod_accum_113__60_,
  prod_accum_113__59_,prod_accum_113__58_,prod_accum_113__57_,prod_accum_113__56_,
  prod_accum_113__55_,prod_accum_113__54_,prod_accum_113__53_,prod_accum_113__52_,
  prod_accum_113__51_,prod_accum_113__50_,prod_accum_113__49_,prod_accum_113__48_,
  prod_accum_113__47_,prod_accum_113__46_,prod_accum_113__45_,prod_accum_113__44_,
  prod_accum_113__43_,prod_accum_113__42_,prod_accum_113__41_,prod_accum_113__40_,
  prod_accum_113__39_,prod_accum_113__38_,prod_accum_113__37_,prod_accum_113__36_,
  prod_accum_113__35_,prod_accum_113__34_,prod_accum_113__33_,prod_accum_113__32_,
  prod_accum_113__31_,prod_accum_113__30_,prod_accum_113__29_,prod_accum_113__28_,
  prod_accum_113__27_,prod_accum_113__26_,prod_accum_113__25_,prod_accum_113__24_,
  prod_accum_113__23_,prod_accum_113__22_,prod_accum_113__21_,prod_accum_113__20_,
  prod_accum_113__19_,prod_accum_113__18_,prod_accum_113__17_,prod_accum_113__16_,
  prod_accum_113__15_,prod_accum_113__14_,prod_accum_113__13_,prod_accum_113__12_,
  prod_accum_113__11_,prod_accum_113__10_,prod_accum_113__9_,prod_accum_113__8_,
  prod_accum_113__7_,prod_accum_113__6_,prod_accum_113__5_,prod_accum_113__4_,
  prod_accum_113__3_,prod_accum_113__2_,prod_accum_113__1_,prod_accum_113__0_,
  prod_accum_112__113_,prod_accum_112__112_,prod_accum_112__111_,prod_accum_112__110_,
  prod_accum_112__109_,prod_accum_112__108_,prod_accum_112__107_,prod_accum_112__106_,
  prod_accum_112__105_,prod_accum_112__104_,prod_accum_112__103_,
  prod_accum_112__102_,prod_accum_112__101_,prod_accum_112__100_,prod_accum_112__99_,
  prod_accum_112__98_,prod_accum_112__97_,prod_accum_112__96_,prod_accum_112__95_,
  prod_accum_112__94_,prod_accum_112__93_,prod_accum_112__92_,prod_accum_112__91_,
  prod_accum_112__90_,prod_accum_112__89_,prod_accum_112__88_,prod_accum_112__87_,
  prod_accum_112__86_,prod_accum_112__85_,prod_accum_112__84_,prod_accum_112__83_,
  prod_accum_112__82_,prod_accum_112__81_,prod_accum_112__80_,prod_accum_112__79_,
  prod_accum_112__78_,prod_accum_112__77_,prod_accum_112__76_,prod_accum_112__75_,
  prod_accum_112__74_,prod_accum_112__73_,prod_accum_112__72_,prod_accum_112__71_,
  prod_accum_112__70_,prod_accum_112__69_,prod_accum_112__68_,prod_accum_112__67_,
  prod_accum_112__66_,prod_accum_112__65_,prod_accum_112__64_,prod_accum_112__63_,
  prod_accum_112__62_,prod_accum_112__61_,prod_accum_112__60_,prod_accum_112__59_,
  prod_accum_112__58_,prod_accum_112__57_,prod_accum_112__56_,prod_accum_112__55_,
  prod_accum_112__54_,prod_accum_112__53_,prod_accum_112__52_,prod_accum_112__51_,
  prod_accum_112__50_,prod_accum_112__49_,prod_accum_112__48_,prod_accum_112__47_,
  prod_accum_112__46_,prod_accum_112__45_,prod_accum_112__44_,prod_accum_112__43_,
  prod_accum_112__42_,prod_accum_112__41_,prod_accum_112__40_,prod_accum_112__39_,
  prod_accum_112__38_,prod_accum_112__37_,prod_accum_112__36_,prod_accum_112__35_,
  prod_accum_112__34_,prod_accum_112__33_,prod_accum_112__32_,prod_accum_112__31_,
  prod_accum_112__30_,prod_accum_112__29_,prod_accum_112__28_,prod_accum_112__27_,
  prod_accum_112__26_,prod_accum_112__25_,prod_accum_112__24_,prod_accum_112__23_,
  prod_accum_112__22_,prod_accum_112__21_,prod_accum_112__20_,prod_accum_112__19_,
  prod_accum_112__18_,prod_accum_112__17_,prod_accum_112__16_,prod_accum_112__15_,
  prod_accum_112__14_,prod_accum_112__13_,prod_accum_112__12_,prod_accum_112__11_,
  prod_accum_112__10_,prod_accum_112__9_,prod_accum_112__8_,prod_accum_112__7_,prod_accum_112__6_,
  prod_accum_112__5_,prod_accum_112__4_,prod_accum_112__3_,prod_accum_112__2_,
  prod_accum_112__1_,prod_accum_112__0_,prod_accum_111__112_,prod_accum_111__111_,
  prod_accum_111__110_,prod_accum_111__109_,prod_accum_111__108_,prod_accum_111__107_,
  prod_accum_111__106_,prod_accum_111__105_,prod_accum_111__104_,
  prod_accum_111__103_,prod_accum_111__102_,prod_accum_111__101_,prod_accum_111__100_,
  prod_accum_111__99_,prod_accum_111__98_,prod_accum_111__97_,prod_accum_111__96_,
  prod_accum_111__95_,prod_accum_111__94_,prod_accum_111__93_,prod_accum_111__92_,
  prod_accum_111__91_,prod_accum_111__90_,prod_accum_111__89_,prod_accum_111__88_,
  prod_accum_111__87_,prod_accum_111__86_,prod_accum_111__85_,prod_accum_111__84_,
  prod_accum_111__83_,prod_accum_111__82_,prod_accum_111__81_,prod_accum_111__80_,
  prod_accum_111__79_,prod_accum_111__78_,prod_accum_111__77_,prod_accum_111__76_,
  prod_accum_111__75_,prod_accum_111__74_,prod_accum_111__73_,prod_accum_111__72_,
  prod_accum_111__71_,prod_accum_111__70_,prod_accum_111__69_,prod_accum_111__68_,
  prod_accum_111__67_,prod_accum_111__66_,prod_accum_111__65_,prod_accum_111__64_,
  prod_accum_111__63_,prod_accum_111__62_,prod_accum_111__61_,prod_accum_111__60_,
  prod_accum_111__59_,prod_accum_111__58_,prod_accum_111__57_,prod_accum_111__56_,
  prod_accum_111__55_,prod_accum_111__54_,prod_accum_111__53_,prod_accum_111__52_,
  prod_accum_111__51_,prod_accum_111__50_,prod_accum_111__49_,prod_accum_111__48_,
  prod_accum_111__47_,prod_accum_111__46_,prod_accum_111__45_,prod_accum_111__44_,
  prod_accum_111__43_,prod_accum_111__42_,prod_accum_111__41_,prod_accum_111__40_,
  prod_accum_111__39_,prod_accum_111__38_,prod_accum_111__37_,prod_accum_111__36_,
  prod_accum_111__35_,prod_accum_111__34_,prod_accum_111__33_,prod_accum_111__32_,
  prod_accum_111__31_,prod_accum_111__30_,prod_accum_111__29_,prod_accum_111__28_,
  prod_accum_111__27_,prod_accum_111__26_,prod_accum_111__25_,prod_accum_111__24_,
  prod_accum_111__23_,prod_accum_111__22_,prod_accum_111__21_,prod_accum_111__20_,
  prod_accum_111__19_,prod_accum_111__18_,prod_accum_111__17_,prod_accum_111__16_,
  prod_accum_111__15_,prod_accum_111__14_,prod_accum_111__13_,prod_accum_111__12_,
  prod_accum_111__11_,prod_accum_111__10_,prod_accum_111__9_,prod_accum_111__8_,
  prod_accum_111__7_,prod_accum_111__6_,prod_accum_111__5_,prod_accum_111__4_,prod_accum_111__3_,
  prod_accum_111__2_,prod_accum_111__1_,prod_accum_111__0_,s_r_118__127_,
  s_r_118__126_,s_r_118__125_,s_r_118__124_,s_r_118__123_,s_r_118__122_,s_r_118__121_,
  s_r_118__120_,s_r_118__119_,s_r_118__118_,s_r_118__117_,s_r_118__116_,s_r_118__115_,
  s_r_118__114_,s_r_118__113_,s_r_118__112_,s_r_118__111_,s_r_118__110_,
  s_r_118__109_,s_r_118__108_,s_r_118__107_,s_r_118__106_,s_r_118__105_,s_r_118__104_,
  s_r_118__103_,s_r_118__102_,s_r_118__101_,s_r_118__100_,s_r_118__99_,s_r_118__98_,
  s_r_118__97_,s_r_118__96_,s_r_118__95_,s_r_118__94_,s_r_118__93_,s_r_118__92_,
  s_r_118__91_,s_r_118__90_,s_r_118__89_,s_r_118__88_,s_r_118__87_,s_r_118__86_,
  s_r_118__85_,s_r_118__84_,s_r_118__83_,s_r_118__82_,s_r_118__81_,s_r_118__80_,
  s_r_118__79_,s_r_118__78_,s_r_118__77_,s_r_118__76_,s_r_118__75_,s_r_118__74_,s_r_118__73_,
  s_r_118__72_,s_r_118__71_,s_r_118__70_,s_r_118__69_,s_r_118__68_,s_r_118__67_,
  s_r_118__66_,s_r_118__65_,s_r_118__64_,s_r_118__63_,s_r_118__62_,s_r_118__61_,
  s_r_118__60_,s_r_118__59_,s_r_118__58_,s_r_118__57_,s_r_118__56_,s_r_118__55_,
  s_r_118__54_,s_r_118__53_,s_r_118__52_,s_r_118__51_,s_r_118__50_,s_r_118__49_,
  s_r_118__48_,s_r_118__47_,s_r_118__46_,s_r_118__45_,s_r_118__44_,s_r_118__43_,
  s_r_118__42_,s_r_118__41_,s_r_118__40_,s_r_118__39_,s_r_118__38_,s_r_118__37_,
  s_r_118__36_,s_r_118__35_,s_r_118__34_,s_r_118__33_,s_r_118__32_,s_r_118__31_,s_r_118__30_,
  s_r_118__29_,s_r_118__28_,s_r_118__27_,s_r_118__26_,s_r_118__25_,s_r_118__24_,
  s_r_118__23_,s_r_118__22_,s_r_118__21_,s_r_118__20_,s_r_118__19_,s_r_118__18_,
  s_r_118__17_,s_r_118__16_,s_r_118__15_,s_r_118__14_,s_r_118__13_,s_r_118__12_,
  s_r_118__11_,s_r_118__10_,s_r_118__9_,s_r_118__8_,s_r_118__7_,s_r_118__6_,s_r_118__5_,
  s_r_118__4_,s_r_118__3_,s_r_118__2_,s_r_118__1_,s_r_118__0_,s_r_117__127_,
  s_r_117__126_,s_r_117__125_,s_r_117__124_,s_r_117__123_,s_r_117__122_,s_r_117__121_,
  s_r_117__120_,s_r_117__119_,s_r_117__118_,s_r_117__117_,s_r_117__116_,
  s_r_117__115_,s_r_117__114_,s_r_117__113_,s_r_117__112_,s_r_117__111_,s_r_117__110_,
  s_r_117__109_,s_r_117__108_,s_r_117__107_,s_r_117__106_,s_r_117__105_,s_r_117__104_,
  s_r_117__103_,s_r_117__102_,s_r_117__101_,s_r_117__100_,s_r_117__99_,s_r_117__98_,
  s_r_117__97_,s_r_117__96_,s_r_117__95_,s_r_117__94_,s_r_117__93_,s_r_117__92_,
  s_r_117__91_,s_r_117__90_,s_r_117__89_,s_r_117__88_,s_r_117__87_,s_r_117__86_,
  s_r_117__85_,s_r_117__84_,s_r_117__83_,s_r_117__82_,s_r_117__81_,s_r_117__80_,
  s_r_117__79_,s_r_117__78_,s_r_117__77_,s_r_117__76_,s_r_117__75_,s_r_117__74_,
  s_r_117__73_,s_r_117__72_,s_r_117__71_,s_r_117__70_,s_r_117__69_,s_r_117__68_,s_r_117__67_,
  s_r_117__66_,s_r_117__65_,s_r_117__64_,s_r_117__63_,s_r_117__62_,s_r_117__61_,
  s_r_117__60_,s_r_117__59_,s_r_117__58_,s_r_117__57_,s_r_117__56_,s_r_117__55_,
  s_r_117__54_,s_r_117__53_,s_r_117__52_,s_r_117__51_,s_r_117__50_,s_r_117__49_,
  s_r_117__48_,s_r_117__47_,s_r_117__46_,s_r_117__45_,s_r_117__44_,s_r_117__43_,
  s_r_117__42_,s_r_117__41_,s_r_117__40_,s_r_117__39_,s_r_117__38_,s_r_117__37_,
  s_r_117__36_,s_r_117__35_,s_r_117__34_,s_r_117__33_,s_r_117__32_,s_r_117__31_,
  s_r_117__30_,s_r_117__29_,s_r_117__28_,s_r_117__27_,s_r_117__26_,s_r_117__25_,s_r_117__24_,
  s_r_117__23_,s_r_117__22_,s_r_117__21_,s_r_117__20_,s_r_117__19_,s_r_117__18_,
  s_r_117__17_,s_r_117__16_,s_r_117__15_,s_r_117__14_,s_r_117__13_,s_r_117__12_,
  s_r_117__11_,s_r_117__10_,s_r_117__9_,s_r_117__8_,s_r_117__7_,s_r_117__6_,
  s_r_117__5_,s_r_117__4_,s_r_117__3_,s_r_117__2_,s_r_117__1_,s_r_117__0_,s_r_116__127_,
  s_r_116__126_,s_r_116__125_,s_r_116__124_,s_r_116__123_,s_r_116__122_,s_r_116__121_,
  s_r_116__120_,s_r_116__119_,s_r_116__118_,s_r_116__117_,s_r_116__116_,
  s_r_116__115_,s_r_116__114_,s_r_116__113_,s_r_116__112_,s_r_116__111_,s_r_116__110_,
  s_r_116__109_,s_r_116__108_,s_r_116__107_,s_r_116__106_,s_r_116__105_,s_r_116__104_,
  s_r_116__103_,s_r_116__102_,s_r_116__101_,s_r_116__100_,s_r_116__99_,s_r_116__98_,
  s_r_116__97_,s_r_116__96_,s_r_116__95_,s_r_116__94_,s_r_116__93_,s_r_116__92_,
  s_r_116__91_,s_r_116__90_,s_r_116__89_,s_r_116__88_,s_r_116__87_,s_r_116__86_,
  s_r_116__85_,s_r_116__84_,s_r_116__83_,s_r_116__82_,s_r_116__81_,s_r_116__80_,
  s_r_116__79_,s_r_116__78_,s_r_116__77_,s_r_116__76_,s_r_116__75_,s_r_116__74_,
  s_r_116__73_,s_r_116__72_,s_r_116__71_,s_r_116__70_,s_r_116__69_,s_r_116__68_,
  s_r_116__67_,s_r_116__66_,s_r_116__65_,s_r_116__64_,s_r_116__63_,s_r_116__62_,s_r_116__61_,
  s_r_116__60_,s_r_116__59_,s_r_116__58_,s_r_116__57_,s_r_116__56_,s_r_116__55_,
  s_r_116__54_,s_r_116__53_,s_r_116__52_,s_r_116__51_,s_r_116__50_,s_r_116__49_,
  s_r_116__48_,s_r_116__47_,s_r_116__46_,s_r_116__45_,s_r_116__44_,s_r_116__43_,
  s_r_116__42_,s_r_116__41_,s_r_116__40_,s_r_116__39_,s_r_116__38_,s_r_116__37_,
  s_r_116__36_,s_r_116__35_,s_r_116__34_,s_r_116__33_,s_r_116__32_,s_r_116__31_,
  s_r_116__30_,s_r_116__29_,s_r_116__28_,s_r_116__27_,s_r_116__26_,s_r_116__25_,
  s_r_116__24_,s_r_116__23_,s_r_116__22_,s_r_116__21_,s_r_116__20_,s_r_116__19_,s_r_116__18_,
  s_r_116__17_,s_r_116__16_,s_r_116__15_,s_r_116__14_,s_r_116__13_,s_r_116__12_,
  s_r_116__11_,s_r_116__10_,s_r_116__9_,s_r_116__8_,s_r_116__7_,s_r_116__6_,
  s_r_116__5_,s_r_116__4_,s_r_116__3_,s_r_116__2_,s_r_116__1_,s_r_116__0_,s_r_115__127_,
  s_r_115__126_,s_r_115__125_,s_r_115__124_,s_r_115__123_,s_r_115__122_,
  s_r_115__121_,s_r_115__120_,s_r_115__119_,s_r_115__118_,s_r_115__117_,s_r_115__116_,
  s_r_115__115_,s_r_115__114_,s_r_115__113_,s_r_115__112_,s_r_115__111_,s_r_115__110_,
  s_r_115__109_,s_r_115__108_,s_r_115__107_,s_r_115__106_,s_r_115__105_,s_r_115__104_,
  s_r_115__103_,s_r_115__102_,s_r_115__101_,s_r_115__100_,s_r_115__99_,
  s_r_115__98_,s_r_115__97_,s_r_115__96_,s_r_115__95_,s_r_115__94_,s_r_115__93_,s_r_115__92_,
  s_r_115__91_,s_r_115__90_,s_r_115__89_,s_r_115__88_,s_r_115__87_,s_r_115__86_,
  s_r_115__85_,s_r_115__84_,s_r_115__83_,s_r_115__82_,s_r_115__81_,s_r_115__80_,
  s_r_115__79_,s_r_115__78_,s_r_115__77_,s_r_115__76_,s_r_115__75_,s_r_115__74_,
  s_r_115__73_,s_r_115__72_,s_r_115__71_,s_r_115__70_,s_r_115__69_,s_r_115__68_,
  s_r_115__67_,s_r_115__66_,s_r_115__65_,s_r_115__64_,s_r_115__63_,s_r_115__62_,
  s_r_115__61_,s_r_115__60_,s_r_115__59_,s_r_115__58_,s_r_115__57_,s_r_115__56_,s_r_115__55_,
  s_r_115__54_,s_r_115__53_,s_r_115__52_,s_r_115__51_,s_r_115__50_,s_r_115__49_,
  s_r_115__48_,s_r_115__47_,s_r_115__46_,s_r_115__45_,s_r_115__44_,s_r_115__43_,
  s_r_115__42_,s_r_115__41_,s_r_115__40_,s_r_115__39_,s_r_115__38_,s_r_115__37_,
  s_r_115__36_,s_r_115__35_,s_r_115__34_,s_r_115__33_,s_r_115__32_,s_r_115__31_,
  s_r_115__30_,s_r_115__29_,s_r_115__28_,s_r_115__27_,s_r_115__26_,s_r_115__25_,
  s_r_115__24_,s_r_115__23_,s_r_115__22_,s_r_115__21_,s_r_115__20_,s_r_115__19_,
  s_r_115__18_,s_r_115__17_,s_r_115__16_,s_r_115__15_,s_r_115__14_,s_r_115__13_,s_r_115__12_,
  s_r_115__11_,s_r_115__10_,s_r_115__9_,s_r_115__8_,s_r_115__7_,s_r_115__6_,
  s_r_115__5_,s_r_115__4_,s_r_115__3_,s_r_115__2_,s_r_115__1_,s_r_115__0_,
  prod_accum_118__119_,prod_accum_118__118_,prod_accum_118__117_,prod_accum_118__116_,
  prod_accum_118__115_,prod_accum_118__114_,prod_accum_118__113_,prod_accum_118__112_,
  prod_accum_118__111_,prod_accum_118__110_,prod_accum_118__109_,prod_accum_118__108_,
  prod_accum_118__107_,prod_accum_118__106_,prod_accum_118__105_,
  prod_accum_118__104_,prod_accum_118__103_,prod_accum_118__102_,prod_accum_118__101_,
  prod_accum_118__100_,prod_accum_118__99_,prod_accum_118__98_,prod_accum_118__97_,
  prod_accum_118__96_,prod_accum_118__95_,prod_accum_118__94_,prod_accum_118__93_,
  prod_accum_118__92_,prod_accum_118__91_,prod_accum_118__90_,prod_accum_118__89_,
  prod_accum_118__88_,prod_accum_118__87_,prod_accum_118__86_,prod_accum_118__85_,
  prod_accum_118__84_,prod_accum_118__83_,prod_accum_118__82_,prod_accum_118__81_,
  prod_accum_118__80_,prod_accum_118__79_,prod_accum_118__78_,prod_accum_118__77_,
  prod_accum_118__76_,prod_accum_118__75_,prod_accum_118__74_,prod_accum_118__73_,
  prod_accum_118__72_,prod_accum_118__71_,prod_accum_118__70_,prod_accum_118__69_,
  prod_accum_118__68_,prod_accum_118__67_,prod_accum_118__66_,prod_accum_118__65_,
  prod_accum_118__64_,prod_accum_118__63_,prod_accum_118__62_,prod_accum_118__61_,
  prod_accum_118__60_,prod_accum_118__59_,prod_accum_118__58_,prod_accum_118__57_,
  prod_accum_118__56_,prod_accum_118__55_,prod_accum_118__54_,prod_accum_118__53_,
  prod_accum_118__52_,prod_accum_118__51_,prod_accum_118__50_,prod_accum_118__49_,
  prod_accum_118__48_,prod_accum_118__47_,prod_accum_118__46_,prod_accum_118__45_,
  prod_accum_118__44_,prod_accum_118__43_,prod_accum_118__42_,prod_accum_118__41_,
  prod_accum_118__40_,prod_accum_118__39_,prod_accum_118__38_,prod_accum_118__37_,
  prod_accum_118__36_,prod_accum_118__35_,prod_accum_118__34_,prod_accum_118__33_,
  prod_accum_118__32_,prod_accum_118__31_,prod_accum_118__30_,prod_accum_118__29_,
  prod_accum_118__28_,prod_accum_118__27_,prod_accum_118__26_,prod_accum_118__25_,
  prod_accum_118__24_,prod_accum_118__23_,prod_accum_118__22_,prod_accum_118__21_,
  prod_accum_118__20_,prod_accum_118__19_,prod_accum_118__18_,prod_accum_118__17_,
  prod_accum_118__16_,prod_accum_118__15_,prod_accum_118__14_,prod_accum_118__13_,
  prod_accum_118__12_,prod_accum_118__11_,prod_accum_118__10_,prod_accum_118__9_,
  prod_accum_118__8_,prod_accum_118__7_,prod_accum_118__6_,prod_accum_118__5_,prod_accum_118__4_,
  prod_accum_118__3_,prod_accum_118__2_,prod_accum_118__1_,prod_accum_118__0_,
  prod_accum_117__118_,prod_accum_117__117_,prod_accum_117__116_,prod_accum_117__115_,
  prod_accum_117__114_,prod_accum_117__113_,prod_accum_117__112_,
  prod_accum_117__111_,prod_accum_117__110_,prod_accum_117__109_,prod_accum_117__108_,
  prod_accum_117__107_,prod_accum_117__106_,prod_accum_117__105_,prod_accum_117__104_,
  prod_accum_117__103_,prod_accum_117__102_,prod_accum_117__101_,prod_accum_117__100_,
  prod_accum_117__99_,prod_accum_117__98_,prod_accum_117__97_,prod_accum_117__96_,
  prod_accum_117__95_,prod_accum_117__94_,prod_accum_117__93_,prod_accum_117__92_,
  prod_accum_117__91_,prod_accum_117__90_,prod_accum_117__89_,prod_accum_117__88_,
  prod_accum_117__87_,prod_accum_117__86_,prod_accum_117__85_,prod_accum_117__84_,
  prod_accum_117__83_,prod_accum_117__82_,prod_accum_117__81_,prod_accum_117__80_,
  prod_accum_117__79_,prod_accum_117__78_,prod_accum_117__77_,prod_accum_117__76_,
  prod_accum_117__75_,prod_accum_117__74_,prod_accum_117__73_,prod_accum_117__72_,
  prod_accum_117__71_,prod_accum_117__70_,prod_accum_117__69_,prod_accum_117__68_,
  prod_accum_117__67_,prod_accum_117__66_,prod_accum_117__65_,prod_accum_117__64_,
  prod_accum_117__63_,prod_accum_117__62_,prod_accum_117__61_,prod_accum_117__60_,
  prod_accum_117__59_,prod_accum_117__58_,prod_accum_117__57_,prod_accum_117__56_,
  prod_accum_117__55_,prod_accum_117__54_,prod_accum_117__53_,prod_accum_117__52_,
  prod_accum_117__51_,prod_accum_117__50_,prod_accum_117__49_,prod_accum_117__48_,
  prod_accum_117__47_,prod_accum_117__46_,prod_accum_117__45_,prod_accum_117__44_,
  prod_accum_117__43_,prod_accum_117__42_,prod_accum_117__41_,prod_accum_117__40_,
  prod_accum_117__39_,prod_accum_117__38_,prod_accum_117__37_,prod_accum_117__36_,
  prod_accum_117__35_,prod_accum_117__34_,prod_accum_117__33_,prod_accum_117__32_,
  prod_accum_117__31_,prod_accum_117__30_,prod_accum_117__29_,prod_accum_117__28_,
  prod_accum_117__27_,prod_accum_117__26_,prod_accum_117__25_,prod_accum_117__24_,
  prod_accum_117__23_,prod_accum_117__22_,prod_accum_117__21_,prod_accum_117__20_,
  prod_accum_117__19_,prod_accum_117__18_,prod_accum_117__17_,prod_accum_117__16_,
  prod_accum_117__15_,prod_accum_117__14_,prod_accum_117__13_,prod_accum_117__12_,
  prod_accum_117__11_,prod_accum_117__10_,prod_accum_117__9_,prod_accum_117__8_,
  prod_accum_117__7_,prod_accum_117__6_,prod_accum_117__5_,prod_accum_117__4_,
  prod_accum_117__3_,prod_accum_117__2_,prod_accum_117__1_,prod_accum_117__0_,
  prod_accum_116__117_,prod_accum_116__116_,prod_accum_116__115_,prod_accum_116__114_,
  prod_accum_116__113_,prod_accum_116__112_,prod_accum_116__111_,prod_accum_116__110_,
  prod_accum_116__109_,prod_accum_116__108_,prod_accum_116__107_,prod_accum_116__106_,
  prod_accum_116__105_,prod_accum_116__104_,prod_accum_116__103_,prod_accum_116__102_,
  prod_accum_116__101_,prod_accum_116__100_,prod_accum_116__99_,
  prod_accum_116__98_,prod_accum_116__97_,prod_accum_116__96_,prod_accum_116__95_,
  prod_accum_116__94_,prod_accum_116__93_,prod_accum_116__92_,prod_accum_116__91_,
  prod_accum_116__90_,prod_accum_116__89_,prod_accum_116__88_,prod_accum_116__87_,
  prod_accum_116__86_,prod_accum_116__85_,prod_accum_116__84_,prod_accum_116__83_,
  prod_accum_116__82_,prod_accum_116__81_,prod_accum_116__80_,prod_accum_116__79_,
  prod_accum_116__78_,prod_accum_116__77_,prod_accum_116__76_,prod_accum_116__75_,
  prod_accum_116__74_,prod_accum_116__73_,prod_accum_116__72_,prod_accum_116__71_,
  prod_accum_116__70_,prod_accum_116__69_,prod_accum_116__68_,prod_accum_116__67_,
  prod_accum_116__66_,prod_accum_116__65_,prod_accum_116__64_,prod_accum_116__63_,
  prod_accum_116__62_,prod_accum_116__61_,prod_accum_116__60_,prod_accum_116__59_,
  prod_accum_116__58_,prod_accum_116__57_,prod_accum_116__56_,prod_accum_116__55_,
  prod_accum_116__54_,prod_accum_116__53_,prod_accum_116__52_,prod_accum_116__51_,
  prod_accum_116__50_,prod_accum_116__49_,prod_accum_116__48_,prod_accum_116__47_,
  prod_accum_116__46_,prod_accum_116__45_,prod_accum_116__44_,prod_accum_116__43_,
  prod_accum_116__42_,prod_accum_116__41_,prod_accum_116__40_,prod_accum_116__39_,
  prod_accum_116__38_,prod_accum_116__37_,prod_accum_116__36_,prod_accum_116__35_,
  prod_accum_116__34_,prod_accum_116__33_,prod_accum_116__32_,prod_accum_116__31_,
  prod_accum_116__30_,prod_accum_116__29_,prod_accum_116__28_,prod_accum_116__27_,
  prod_accum_116__26_,prod_accum_116__25_,prod_accum_116__24_,prod_accum_116__23_,
  prod_accum_116__22_,prod_accum_116__21_,prod_accum_116__20_,prod_accum_116__19_,
  prod_accum_116__18_,prod_accum_116__17_,prod_accum_116__16_,prod_accum_116__15_,
  prod_accum_116__14_,prod_accum_116__13_,prod_accum_116__12_,prod_accum_116__11_,
  prod_accum_116__10_,prod_accum_116__9_,prod_accum_116__8_,prod_accum_116__7_,prod_accum_116__6_,
  prod_accum_116__5_,prod_accum_116__4_,prod_accum_116__3_,prod_accum_116__2_,
  prod_accum_116__1_,prod_accum_116__0_,prod_accum_115__116_,prod_accum_115__115_,
  prod_accum_115__114_,prod_accum_115__113_,prod_accum_115__112_,prod_accum_115__111_,
  prod_accum_115__110_,prod_accum_115__109_,prod_accum_115__108_,
  prod_accum_115__107_,prod_accum_115__106_,prod_accum_115__105_,prod_accum_115__104_,
  prod_accum_115__103_,prod_accum_115__102_,prod_accum_115__101_,prod_accum_115__100_,
  prod_accum_115__99_,prod_accum_115__98_,prod_accum_115__97_,prod_accum_115__96_,
  prod_accum_115__95_,prod_accum_115__94_,prod_accum_115__93_,prod_accum_115__92_,
  prod_accum_115__91_,prod_accum_115__90_,prod_accum_115__89_,prod_accum_115__88_,
  prod_accum_115__87_,prod_accum_115__86_,prod_accum_115__85_,prod_accum_115__84_,
  prod_accum_115__83_,prod_accum_115__82_,prod_accum_115__81_,prod_accum_115__80_,
  prod_accum_115__79_,prod_accum_115__78_,prod_accum_115__77_,prod_accum_115__76_,
  prod_accum_115__75_,prod_accum_115__74_,prod_accum_115__73_,prod_accum_115__72_,
  prod_accum_115__71_,prod_accum_115__70_,prod_accum_115__69_,prod_accum_115__68_,
  prod_accum_115__67_,prod_accum_115__66_,prod_accum_115__65_,prod_accum_115__64_,
  prod_accum_115__63_,prod_accum_115__62_,prod_accum_115__61_,prod_accum_115__60_,
  prod_accum_115__59_,prod_accum_115__58_,prod_accum_115__57_,prod_accum_115__56_,
  prod_accum_115__55_,prod_accum_115__54_,prod_accum_115__53_,prod_accum_115__52_,
  prod_accum_115__51_,prod_accum_115__50_,prod_accum_115__49_,prod_accum_115__48_,
  prod_accum_115__47_,prod_accum_115__46_,prod_accum_115__45_,prod_accum_115__44_,
  prod_accum_115__43_,prod_accum_115__42_,prod_accum_115__41_,prod_accum_115__40_,
  prod_accum_115__39_,prod_accum_115__38_,prod_accum_115__37_,prod_accum_115__36_,
  prod_accum_115__35_,prod_accum_115__34_,prod_accum_115__33_,prod_accum_115__32_,
  prod_accum_115__31_,prod_accum_115__30_,prod_accum_115__29_,prod_accum_115__28_,
  prod_accum_115__27_,prod_accum_115__26_,prod_accum_115__25_,prod_accum_115__24_,
  prod_accum_115__23_,prod_accum_115__22_,prod_accum_115__21_,prod_accum_115__20_,
  prod_accum_115__19_,prod_accum_115__18_,prod_accum_115__17_,prod_accum_115__16_,
  prod_accum_115__15_,prod_accum_115__14_,prod_accum_115__13_,prod_accum_115__12_,
  prod_accum_115__11_,prod_accum_115__10_,prod_accum_115__9_,prod_accum_115__8_,
  prod_accum_115__7_,prod_accum_115__6_,prod_accum_115__5_,prod_accum_115__4_,
  prod_accum_115__3_,prod_accum_115__2_,prod_accum_115__1_,prod_accum_115__0_,s_r_122__127_,
  s_r_122__126_,s_r_122__125_,s_r_122__124_,s_r_122__123_,s_r_122__122_,s_r_122__121_,
  s_r_122__120_,s_r_122__119_,s_r_122__118_,s_r_122__117_,s_r_122__116_,
  s_r_122__115_,s_r_122__114_,s_r_122__113_,s_r_122__112_,s_r_122__111_,s_r_122__110_,
  s_r_122__109_,s_r_122__108_,s_r_122__107_,s_r_122__106_,s_r_122__105_,s_r_122__104_,
  s_r_122__103_,s_r_122__102_,s_r_122__101_,s_r_122__100_,s_r_122__99_,s_r_122__98_,
  s_r_122__97_,s_r_122__96_,s_r_122__95_,s_r_122__94_,s_r_122__93_,s_r_122__92_,
  s_r_122__91_,s_r_122__90_,s_r_122__89_,s_r_122__88_,s_r_122__87_,s_r_122__86_,
  s_r_122__85_,s_r_122__84_,s_r_122__83_,s_r_122__82_,s_r_122__81_,s_r_122__80_,
  s_r_122__79_,s_r_122__78_,s_r_122__77_,s_r_122__76_,s_r_122__75_,s_r_122__74_,
  s_r_122__73_,s_r_122__72_,s_r_122__71_,s_r_122__70_,s_r_122__69_,s_r_122__68_,s_r_122__67_,
  s_r_122__66_,s_r_122__65_,s_r_122__64_,s_r_122__63_,s_r_122__62_,s_r_122__61_,
  s_r_122__60_,s_r_122__59_,s_r_122__58_,s_r_122__57_,s_r_122__56_,s_r_122__55_,
  s_r_122__54_,s_r_122__53_,s_r_122__52_,s_r_122__51_,s_r_122__50_,s_r_122__49_,
  s_r_122__48_,s_r_122__47_,s_r_122__46_,s_r_122__45_,s_r_122__44_,s_r_122__43_,
  s_r_122__42_,s_r_122__41_,s_r_122__40_,s_r_122__39_,s_r_122__38_,s_r_122__37_,
  s_r_122__36_,s_r_122__35_,s_r_122__34_,s_r_122__33_,s_r_122__32_,s_r_122__31_,
  s_r_122__30_,s_r_122__29_,s_r_122__28_,s_r_122__27_,s_r_122__26_,s_r_122__25_,s_r_122__24_,
  s_r_122__23_,s_r_122__22_,s_r_122__21_,s_r_122__20_,s_r_122__19_,s_r_122__18_,
  s_r_122__17_,s_r_122__16_,s_r_122__15_,s_r_122__14_,s_r_122__13_,s_r_122__12_,
  s_r_122__11_,s_r_122__10_,s_r_122__9_,s_r_122__8_,s_r_122__7_,s_r_122__6_,
  s_r_122__5_,s_r_122__4_,s_r_122__3_,s_r_122__2_,s_r_122__1_,s_r_122__0_,s_r_121__127_,
  s_r_121__126_,s_r_121__125_,s_r_121__124_,s_r_121__123_,s_r_121__122_,s_r_121__121_,
  s_r_121__120_,s_r_121__119_,s_r_121__118_,s_r_121__117_,s_r_121__116_,
  s_r_121__115_,s_r_121__114_,s_r_121__113_,s_r_121__112_,s_r_121__111_,s_r_121__110_,
  s_r_121__109_,s_r_121__108_,s_r_121__107_,s_r_121__106_,s_r_121__105_,s_r_121__104_,
  s_r_121__103_,s_r_121__102_,s_r_121__101_,s_r_121__100_,s_r_121__99_,s_r_121__98_,
  s_r_121__97_,s_r_121__96_,s_r_121__95_,s_r_121__94_,s_r_121__93_,s_r_121__92_,
  s_r_121__91_,s_r_121__90_,s_r_121__89_,s_r_121__88_,s_r_121__87_,s_r_121__86_,
  s_r_121__85_,s_r_121__84_,s_r_121__83_,s_r_121__82_,s_r_121__81_,s_r_121__80_,
  s_r_121__79_,s_r_121__78_,s_r_121__77_,s_r_121__76_,s_r_121__75_,s_r_121__74_,
  s_r_121__73_,s_r_121__72_,s_r_121__71_,s_r_121__70_,s_r_121__69_,s_r_121__68_,
  s_r_121__67_,s_r_121__66_,s_r_121__65_,s_r_121__64_,s_r_121__63_,s_r_121__62_,s_r_121__61_,
  s_r_121__60_,s_r_121__59_,s_r_121__58_,s_r_121__57_,s_r_121__56_,s_r_121__55_,
  s_r_121__54_,s_r_121__53_,s_r_121__52_,s_r_121__51_,s_r_121__50_,s_r_121__49_,
  s_r_121__48_,s_r_121__47_,s_r_121__46_,s_r_121__45_,s_r_121__44_,s_r_121__43_,
  s_r_121__42_,s_r_121__41_,s_r_121__40_,s_r_121__39_,s_r_121__38_,s_r_121__37_,
  s_r_121__36_,s_r_121__35_,s_r_121__34_,s_r_121__33_,s_r_121__32_,s_r_121__31_,
  s_r_121__30_,s_r_121__29_,s_r_121__28_,s_r_121__27_,s_r_121__26_,s_r_121__25_,
  s_r_121__24_,s_r_121__23_,s_r_121__22_,s_r_121__21_,s_r_121__20_,s_r_121__19_,s_r_121__18_,
  s_r_121__17_,s_r_121__16_,s_r_121__15_,s_r_121__14_,s_r_121__13_,s_r_121__12_,
  s_r_121__11_,s_r_121__10_,s_r_121__9_,s_r_121__8_,s_r_121__7_,s_r_121__6_,
  s_r_121__5_,s_r_121__4_,s_r_121__3_,s_r_121__2_,s_r_121__1_,s_r_121__0_,s_r_120__127_,
  s_r_120__126_,s_r_120__125_,s_r_120__124_,s_r_120__123_,s_r_120__122_,
  s_r_120__121_,s_r_120__120_,s_r_120__119_,s_r_120__118_,s_r_120__117_,s_r_120__116_,
  s_r_120__115_,s_r_120__114_,s_r_120__113_,s_r_120__112_,s_r_120__111_,s_r_120__110_,
  s_r_120__109_,s_r_120__108_,s_r_120__107_,s_r_120__106_,s_r_120__105_,s_r_120__104_,
  s_r_120__103_,s_r_120__102_,s_r_120__101_,s_r_120__100_,s_r_120__99_,
  s_r_120__98_,s_r_120__97_,s_r_120__96_,s_r_120__95_,s_r_120__94_,s_r_120__93_,s_r_120__92_,
  s_r_120__91_,s_r_120__90_,s_r_120__89_,s_r_120__88_,s_r_120__87_,s_r_120__86_,
  s_r_120__85_,s_r_120__84_,s_r_120__83_,s_r_120__82_,s_r_120__81_,s_r_120__80_,
  s_r_120__79_,s_r_120__78_,s_r_120__77_,s_r_120__76_,s_r_120__75_,s_r_120__74_,
  s_r_120__73_,s_r_120__72_,s_r_120__71_,s_r_120__70_,s_r_120__69_,s_r_120__68_,
  s_r_120__67_,s_r_120__66_,s_r_120__65_,s_r_120__64_,s_r_120__63_,s_r_120__62_,
  s_r_120__61_,s_r_120__60_,s_r_120__59_,s_r_120__58_,s_r_120__57_,s_r_120__56_,s_r_120__55_,
  s_r_120__54_,s_r_120__53_,s_r_120__52_,s_r_120__51_,s_r_120__50_,s_r_120__49_,
  s_r_120__48_,s_r_120__47_,s_r_120__46_,s_r_120__45_,s_r_120__44_,s_r_120__43_,
  s_r_120__42_,s_r_120__41_,s_r_120__40_,s_r_120__39_,s_r_120__38_,s_r_120__37_,
  s_r_120__36_,s_r_120__35_,s_r_120__34_,s_r_120__33_,s_r_120__32_,s_r_120__31_,
  s_r_120__30_,s_r_120__29_,s_r_120__28_,s_r_120__27_,s_r_120__26_,s_r_120__25_,
  s_r_120__24_,s_r_120__23_,s_r_120__22_,s_r_120__21_,s_r_120__20_,s_r_120__19_,
  s_r_120__18_,s_r_120__17_,s_r_120__16_,s_r_120__15_,s_r_120__14_,s_r_120__13_,s_r_120__12_,
  s_r_120__11_,s_r_120__10_,s_r_120__9_,s_r_120__8_,s_r_120__7_,s_r_120__6_,
  s_r_120__5_,s_r_120__4_,s_r_120__3_,s_r_120__2_,s_r_120__1_,s_r_120__0_,s_r_119__127_,
  s_r_119__126_,s_r_119__125_,s_r_119__124_,s_r_119__123_,s_r_119__122_,
  s_r_119__121_,s_r_119__120_,s_r_119__119_,s_r_119__118_,s_r_119__117_,s_r_119__116_,
  s_r_119__115_,s_r_119__114_,s_r_119__113_,s_r_119__112_,s_r_119__111_,s_r_119__110_,
  s_r_119__109_,s_r_119__108_,s_r_119__107_,s_r_119__106_,s_r_119__105_,
  s_r_119__104_,s_r_119__103_,s_r_119__102_,s_r_119__101_,s_r_119__100_,s_r_119__99_,
  s_r_119__98_,s_r_119__97_,s_r_119__96_,s_r_119__95_,s_r_119__94_,s_r_119__93_,
  s_r_119__92_,s_r_119__91_,s_r_119__90_,s_r_119__89_,s_r_119__88_,s_r_119__87_,s_r_119__86_,
  s_r_119__85_,s_r_119__84_,s_r_119__83_,s_r_119__82_,s_r_119__81_,s_r_119__80_,
  s_r_119__79_,s_r_119__78_,s_r_119__77_,s_r_119__76_,s_r_119__75_,s_r_119__74_,
  s_r_119__73_,s_r_119__72_,s_r_119__71_,s_r_119__70_,s_r_119__69_,s_r_119__68_,
  s_r_119__67_,s_r_119__66_,s_r_119__65_,s_r_119__64_,s_r_119__63_,s_r_119__62_,
  s_r_119__61_,s_r_119__60_,s_r_119__59_,s_r_119__58_,s_r_119__57_,s_r_119__56_,
  s_r_119__55_,s_r_119__54_,s_r_119__53_,s_r_119__52_,s_r_119__51_,s_r_119__50_,s_r_119__49_,
  s_r_119__48_,s_r_119__47_,s_r_119__46_,s_r_119__45_,s_r_119__44_,s_r_119__43_,
  s_r_119__42_,s_r_119__41_,s_r_119__40_,s_r_119__39_,s_r_119__38_,s_r_119__37_,
  s_r_119__36_,s_r_119__35_,s_r_119__34_,s_r_119__33_,s_r_119__32_,s_r_119__31_,
  s_r_119__30_,s_r_119__29_,s_r_119__28_,s_r_119__27_,s_r_119__26_,s_r_119__25_,
  s_r_119__24_,s_r_119__23_,s_r_119__22_,s_r_119__21_,s_r_119__20_,s_r_119__19_,
  s_r_119__18_,s_r_119__17_,s_r_119__16_,s_r_119__15_,s_r_119__14_,s_r_119__13_,
  s_r_119__12_,s_r_119__11_,s_r_119__10_,s_r_119__9_,s_r_119__8_,s_r_119__7_,s_r_119__6_,
  s_r_119__5_,s_r_119__4_,s_r_119__3_,s_r_119__2_,s_r_119__1_,s_r_119__0_,
  prod_accum_122__123_,prod_accum_122__122_,prod_accum_122__121_,prod_accum_122__120_,
  prod_accum_122__119_,prod_accum_122__118_,prod_accum_122__117_,prod_accum_122__116_,
  prod_accum_122__115_,prod_accum_122__114_,prod_accum_122__113_,prod_accum_122__112_,
  prod_accum_122__111_,prod_accum_122__110_,prod_accum_122__109_,
  prod_accum_122__108_,prod_accum_122__107_,prod_accum_122__106_,prod_accum_122__105_,
  prod_accum_122__104_,prod_accum_122__103_,prod_accum_122__102_,prod_accum_122__101_,
  prod_accum_122__100_,prod_accum_122__99_,prod_accum_122__98_,prod_accum_122__97_,
  prod_accum_122__96_,prod_accum_122__95_,prod_accum_122__94_,prod_accum_122__93_,
  prod_accum_122__92_,prod_accum_122__91_,prod_accum_122__90_,prod_accum_122__89_,
  prod_accum_122__88_,prod_accum_122__87_,prod_accum_122__86_,prod_accum_122__85_,
  prod_accum_122__84_,prod_accum_122__83_,prod_accum_122__82_,prod_accum_122__81_,
  prod_accum_122__80_,prod_accum_122__79_,prod_accum_122__78_,prod_accum_122__77_,
  prod_accum_122__76_,prod_accum_122__75_,prod_accum_122__74_,prod_accum_122__73_,
  prod_accum_122__72_,prod_accum_122__71_,prod_accum_122__70_,prod_accum_122__69_,
  prod_accum_122__68_,prod_accum_122__67_,prod_accum_122__66_,prod_accum_122__65_,
  prod_accum_122__64_,prod_accum_122__63_,prod_accum_122__62_,prod_accum_122__61_,
  prod_accum_122__60_,prod_accum_122__59_,prod_accum_122__58_,prod_accum_122__57_,
  prod_accum_122__56_,prod_accum_122__55_,prod_accum_122__54_,prod_accum_122__53_,
  prod_accum_122__52_,prod_accum_122__51_,prod_accum_122__50_,prod_accum_122__49_,
  prod_accum_122__48_,prod_accum_122__47_,prod_accum_122__46_,prod_accum_122__45_,
  prod_accum_122__44_,prod_accum_122__43_,prod_accum_122__42_,prod_accum_122__41_,
  prod_accum_122__40_,prod_accum_122__39_,prod_accum_122__38_,prod_accum_122__37_,
  prod_accum_122__36_,prod_accum_122__35_,prod_accum_122__34_,prod_accum_122__33_,
  prod_accum_122__32_,prod_accum_122__31_,prod_accum_122__30_,prod_accum_122__29_,
  prod_accum_122__28_,prod_accum_122__27_,prod_accum_122__26_,prod_accum_122__25_,
  prod_accum_122__24_,prod_accum_122__23_,prod_accum_122__22_,prod_accum_122__21_,
  prod_accum_122__20_,prod_accum_122__19_,prod_accum_122__18_,prod_accum_122__17_,
  prod_accum_122__16_,prod_accum_122__15_,prod_accum_122__14_,prod_accum_122__13_,
  prod_accum_122__12_,prod_accum_122__11_,prod_accum_122__10_,prod_accum_122__9_,
  prod_accum_122__8_,prod_accum_122__7_,prod_accum_122__6_,prod_accum_122__5_,
  prod_accum_122__4_,prod_accum_122__3_,prod_accum_122__2_,prod_accum_122__1_,
  prod_accum_122__0_,prod_accum_121__122_,prod_accum_121__121_,prod_accum_121__120_,
  prod_accum_121__119_,prod_accum_121__118_,prod_accum_121__117_,prod_accum_121__116_,
  prod_accum_121__115_,prod_accum_121__114_,prod_accum_121__113_,prod_accum_121__112_,
  prod_accum_121__111_,prod_accum_121__110_,prod_accum_121__109_,prod_accum_121__108_,
  prod_accum_121__107_,prod_accum_121__106_,prod_accum_121__105_,prod_accum_121__104_,
  prod_accum_121__103_,prod_accum_121__102_,prod_accum_121__101_,
  prod_accum_121__100_,prod_accum_121__99_,prod_accum_121__98_,prod_accum_121__97_,
  prod_accum_121__96_,prod_accum_121__95_,prod_accum_121__94_,prod_accum_121__93_,
  prod_accum_121__92_,prod_accum_121__91_,prod_accum_121__90_,prod_accum_121__89_,
  prod_accum_121__88_,prod_accum_121__87_,prod_accum_121__86_,prod_accum_121__85_,
  prod_accum_121__84_,prod_accum_121__83_,prod_accum_121__82_,prod_accum_121__81_,
  prod_accum_121__80_,prod_accum_121__79_,prod_accum_121__78_,prod_accum_121__77_,
  prod_accum_121__76_,prod_accum_121__75_,prod_accum_121__74_,prod_accum_121__73_,
  prod_accum_121__72_,prod_accum_121__71_,prod_accum_121__70_,prod_accum_121__69_,
  prod_accum_121__68_,prod_accum_121__67_,prod_accum_121__66_,prod_accum_121__65_,
  prod_accum_121__64_,prod_accum_121__63_,prod_accum_121__62_,prod_accum_121__61_,
  prod_accum_121__60_,prod_accum_121__59_,prod_accum_121__58_,prod_accum_121__57_,
  prod_accum_121__56_,prod_accum_121__55_,prod_accum_121__54_,prod_accum_121__53_,
  prod_accum_121__52_,prod_accum_121__51_,prod_accum_121__50_,prod_accum_121__49_,
  prod_accum_121__48_,prod_accum_121__47_,prod_accum_121__46_,prod_accum_121__45_,
  prod_accum_121__44_,prod_accum_121__43_,prod_accum_121__42_,prod_accum_121__41_,
  prod_accum_121__40_,prod_accum_121__39_,prod_accum_121__38_,prod_accum_121__37_,
  prod_accum_121__36_,prod_accum_121__35_,prod_accum_121__34_,prod_accum_121__33_,
  prod_accum_121__32_,prod_accum_121__31_,prod_accum_121__30_,prod_accum_121__29_,
  prod_accum_121__28_,prod_accum_121__27_,prod_accum_121__26_,prod_accum_121__25_,
  prod_accum_121__24_,prod_accum_121__23_,prod_accum_121__22_,prod_accum_121__21_,
  prod_accum_121__20_,prod_accum_121__19_,prod_accum_121__18_,prod_accum_121__17_,
  prod_accum_121__16_,prod_accum_121__15_,prod_accum_121__14_,prod_accum_121__13_,
  prod_accum_121__12_,prod_accum_121__11_,prod_accum_121__10_,prod_accum_121__9_,
  prod_accum_121__8_,prod_accum_121__7_,prod_accum_121__6_,prod_accum_121__5_,prod_accum_121__4_,
  prod_accum_121__3_,prod_accum_121__2_,prod_accum_121__1_,prod_accum_121__0_,
  prod_accum_120__121_,prod_accum_120__120_,prod_accum_120__119_,prod_accum_120__118_,
  prod_accum_120__117_,prod_accum_120__116_,prod_accum_120__115_,
  prod_accum_120__114_,prod_accum_120__113_,prod_accum_120__112_,prod_accum_120__111_,
  prod_accum_120__110_,prod_accum_120__109_,prod_accum_120__108_,prod_accum_120__107_,
  prod_accum_120__106_,prod_accum_120__105_,prod_accum_120__104_,prod_accum_120__103_,
  prod_accum_120__102_,prod_accum_120__101_,prod_accum_120__100_,prod_accum_120__99_,
  prod_accum_120__98_,prod_accum_120__97_,prod_accum_120__96_,prod_accum_120__95_,
  prod_accum_120__94_,prod_accum_120__93_,prod_accum_120__92_,prod_accum_120__91_,
  prod_accum_120__90_,prod_accum_120__89_,prod_accum_120__88_,prod_accum_120__87_,
  prod_accum_120__86_,prod_accum_120__85_,prod_accum_120__84_,prod_accum_120__83_,
  prod_accum_120__82_,prod_accum_120__81_,prod_accum_120__80_,prod_accum_120__79_,
  prod_accum_120__78_,prod_accum_120__77_,prod_accum_120__76_,prod_accum_120__75_,
  prod_accum_120__74_,prod_accum_120__73_,prod_accum_120__72_,prod_accum_120__71_,
  prod_accum_120__70_,prod_accum_120__69_,prod_accum_120__68_,prod_accum_120__67_,
  prod_accum_120__66_,prod_accum_120__65_,prod_accum_120__64_,prod_accum_120__63_,
  prod_accum_120__62_,prod_accum_120__61_,prod_accum_120__60_,prod_accum_120__59_,
  prod_accum_120__58_,prod_accum_120__57_,prod_accum_120__56_,prod_accum_120__55_,
  prod_accum_120__54_,prod_accum_120__53_,prod_accum_120__52_,prod_accum_120__51_,
  prod_accum_120__50_,prod_accum_120__49_,prod_accum_120__48_,prod_accum_120__47_,
  prod_accum_120__46_,prod_accum_120__45_,prod_accum_120__44_,prod_accum_120__43_,
  prod_accum_120__42_,prod_accum_120__41_,prod_accum_120__40_,prod_accum_120__39_,
  prod_accum_120__38_,prod_accum_120__37_,prod_accum_120__36_,prod_accum_120__35_,
  prod_accum_120__34_,prod_accum_120__33_,prod_accum_120__32_,prod_accum_120__31_,
  prod_accum_120__30_,prod_accum_120__29_,prod_accum_120__28_,prod_accum_120__27_,
  prod_accum_120__26_,prod_accum_120__25_,prod_accum_120__24_,prod_accum_120__23_,
  prod_accum_120__22_,prod_accum_120__21_,prod_accum_120__20_,prod_accum_120__19_,
  prod_accum_120__18_,prod_accum_120__17_,prod_accum_120__16_,prod_accum_120__15_,
  prod_accum_120__14_,prod_accum_120__13_,prod_accum_120__12_,prod_accum_120__11_,
  prod_accum_120__10_,prod_accum_120__9_,prod_accum_120__8_,prod_accum_120__7_,
  prod_accum_120__6_,prod_accum_120__5_,prod_accum_120__4_,prod_accum_120__3_,
  prod_accum_120__2_,prod_accum_120__1_,prod_accum_120__0_,prod_accum_119__120_,
  prod_accum_119__119_,prod_accum_119__118_,prod_accum_119__117_,prod_accum_119__116_,
  prod_accum_119__115_,prod_accum_119__114_,prod_accum_119__113_,prod_accum_119__112_,
  prod_accum_119__111_,prod_accum_119__110_,prod_accum_119__109_,prod_accum_119__108_,
  prod_accum_119__107_,prod_accum_119__106_,prod_accum_119__105_,
  prod_accum_119__104_,prod_accum_119__103_,prod_accum_119__102_,prod_accum_119__101_,
  prod_accum_119__100_,prod_accum_119__99_,prod_accum_119__98_,prod_accum_119__97_,
  prod_accum_119__96_,prod_accum_119__95_,prod_accum_119__94_,prod_accum_119__93_,
  prod_accum_119__92_,prod_accum_119__91_,prod_accum_119__90_,prod_accum_119__89_,
  prod_accum_119__88_,prod_accum_119__87_,prod_accum_119__86_,prod_accum_119__85_,
  prod_accum_119__84_,prod_accum_119__83_,prod_accum_119__82_,prod_accum_119__81_,
  prod_accum_119__80_,prod_accum_119__79_,prod_accum_119__78_,prod_accum_119__77_,
  prod_accum_119__76_,prod_accum_119__75_,prod_accum_119__74_,prod_accum_119__73_,
  prod_accum_119__72_,prod_accum_119__71_,prod_accum_119__70_,prod_accum_119__69_,
  prod_accum_119__68_,prod_accum_119__67_,prod_accum_119__66_,prod_accum_119__65_,
  prod_accum_119__64_,prod_accum_119__63_,prod_accum_119__62_,prod_accum_119__61_,
  prod_accum_119__60_,prod_accum_119__59_,prod_accum_119__58_,prod_accum_119__57_,
  prod_accum_119__56_,prod_accum_119__55_,prod_accum_119__54_,prod_accum_119__53_,
  prod_accum_119__52_,prod_accum_119__51_,prod_accum_119__50_,prod_accum_119__49_,
  prod_accum_119__48_,prod_accum_119__47_,prod_accum_119__46_,prod_accum_119__45_,
  prod_accum_119__44_,prod_accum_119__43_,prod_accum_119__42_,prod_accum_119__41_,
  prod_accum_119__40_,prod_accum_119__39_,prod_accum_119__38_,prod_accum_119__37_,
  prod_accum_119__36_,prod_accum_119__35_,prod_accum_119__34_,prod_accum_119__33_,
  prod_accum_119__32_,prod_accum_119__31_,prod_accum_119__30_,prod_accum_119__29_,
  prod_accum_119__28_,prod_accum_119__27_,prod_accum_119__26_,prod_accum_119__25_,
  prod_accum_119__24_,prod_accum_119__23_,prod_accum_119__22_,prod_accum_119__21_,
  prod_accum_119__20_,prod_accum_119__19_,prod_accum_119__18_,prod_accum_119__17_,
  prod_accum_119__16_,prod_accum_119__15_,prod_accum_119__14_,prod_accum_119__13_,
  prod_accum_119__12_,prod_accum_119__11_,prod_accum_119__10_,prod_accum_119__9_,
  prod_accum_119__8_,prod_accum_119__7_,prod_accum_119__6_,prod_accum_119__5_,
  prod_accum_119__4_,prod_accum_119__3_,prod_accum_119__2_,prod_accum_119__1_,prod_accum_119__0_,
  s_r_125__127_,s_r_125__126_,s_r_125__125_,s_r_125__124_,s_r_125__123_,
  s_r_125__122_,s_r_125__121_,s_r_125__120_,s_r_125__119_,s_r_125__118_,s_r_125__117_,
  s_r_125__116_,s_r_125__115_,s_r_125__114_,s_r_125__113_,s_r_125__112_,s_r_125__111_,
  s_r_125__110_,s_r_125__109_,s_r_125__108_,s_r_125__107_,s_r_125__106_,s_r_125__105_,
  s_r_125__104_,s_r_125__103_,s_r_125__102_,s_r_125__101_,s_r_125__100_,
  s_r_125__99_,s_r_125__98_,s_r_125__97_,s_r_125__96_,s_r_125__95_,s_r_125__94_,s_r_125__93_,
  s_r_125__92_,s_r_125__91_,s_r_125__90_,s_r_125__89_,s_r_125__88_,s_r_125__87_,
  s_r_125__86_,s_r_125__85_,s_r_125__84_,s_r_125__83_,s_r_125__82_,s_r_125__81_,
  s_r_125__80_,s_r_125__79_,s_r_125__78_,s_r_125__77_,s_r_125__76_,s_r_125__75_,
  s_r_125__74_,s_r_125__73_,s_r_125__72_,s_r_125__71_,s_r_125__70_,s_r_125__69_,
  s_r_125__68_,s_r_125__67_,s_r_125__66_,s_r_125__65_,s_r_125__64_,s_r_125__63_,
  s_r_125__62_,s_r_125__61_,s_r_125__60_,s_r_125__59_,s_r_125__58_,s_r_125__57_,
  s_r_125__56_,s_r_125__55_,s_r_125__54_,s_r_125__53_,s_r_125__52_,s_r_125__51_,s_r_125__50_,
  s_r_125__49_,s_r_125__48_,s_r_125__47_,s_r_125__46_,s_r_125__45_,s_r_125__44_,
  s_r_125__43_,s_r_125__42_,s_r_125__41_,s_r_125__40_,s_r_125__39_,s_r_125__38_,
  s_r_125__37_,s_r_125__36_,s_r_125__35_,s_r_125__34_,s_r_125__33_,s_r_125__32_,
  s_r_125__31_,s_r_125__30_,s_r_125__29_,s_r_125__28_,s_r_125__27_,s_r_125__26_,
  s_r_125__25_,s_r_125__24_,s_r_125__23_,s_r_125__22_,s_r_125__21_,s_r_125__20_,
  s_r_125__19_,s_r_125__18_,s_r_125__17_,s_r_125__16_,s_r_125__15_,s_r_125__14_,s_r_125__13_,
  s_r_125__12_,s_r_125__11_,s_r_125__10_,s_r_125__9_,s_r_125__8_,s_r_125__7_,
  s_r_125__6_,s_r_125__5_,s_r_125__4_,s_r_125__3_,s_r_125__2_,s_r_125__1_,s_r_125__0_,
  s_r_124__127_,s_r_124__126_,s_r_124__125_,s_r_124__124_,s_r_124__123_,
  s_r_124__122_,s_r_124__121_,s_r_124__120_,s_r_124__119_,s_r_124__118_,s_r_124__117_,
  s_r_124__116_,s_r_124__115_,s_r_124__114_,s_r_124__113_,s_r_124__112_,s_r_124__111_,
  s_r_124__110_,s_r_124__109_,s_r_124__108_,s_r_124__107_,s_r_124__106_,
  s_r_124__105_,s_r_124__104_,s_r_124__103_,s_r_124__102_,s_r_124__101_,s_r_124__100_,
  s_r_124__99_,s_r_124__98_,s_r_124__97_,s_r_124__96_,s_r_124__95_,s_r_124__94_,
  s_r_124__93_,s_r_124__92_,s_r_124__91_,s_r_124__90_,s_r_124__89_,s_r_124__88_,s_r_124__87_,
  s_r_124__86_,s_r_124__85_,s_r_124__84_,s_r_124__83_,s_r_124__82_,s_r_124__81_,
  s_r_124__80_,s_r_124__79_,s_r_124__78_,s_r_124__77_,s_r_124__76_,s_r_124__75_,
  s_r_124__74_,s_r_124__73_,s_r_124__72_,s_r_124__71_,s_r_124__70_,s_r_124__69_,
  s_r_124__68_,s_r_124__67_,s_r_124__66_,s_r_124__65_,s_r_124__64_,s_r_124__63_,
  s_r_124__62_,s_r_124__61_,s_r_124__60_,s_r_124__59_,s_r_124__58_,s_r_124__57_,
  s_r_124__56_,s_r_124__55_,s_r_124__54_,s_r_124__53_,s_r_124__52_,s_r_124__51_,
  s_r_124__50_,s_r_124__49_,s_r_124__48_,s_r_124__47_,s_r_124__46_,s_r_124__45_,s_r_124__44_,
  s_r_124__43_,s_r_124__42_,s_r_124__41_,s_r_124__40_,s_r_124__39_,s_r_124__38_,
  s_r_124__37_,s_r_124__36_,s_r_124__35_,s_r_124__34_,s_r_124__33_,s_r_124__32_,
  s_r_124__31_,s_r_124__30_,s_r_124__29_,s_r_124__28_,s_r_124__27_,s_r_124__26_,
  s_r_124__25_,s_r_124__24_,s_r_124__23_,s_r_124__22_,s_r_124__21_,s_r_124__20_,
  s_r_124__19_,s_r_124__18_,s_r_124__17_,s_r_124__16_,s_r_124__15_,s_r_124__14_,
  s_r_124__13_,s_r_124__12_,s_r_124__11_,s_r_124__10_,s_r_124__9_,s_r_124__8_,s_r_124__7_,
  s_r_124__6_,s_r_124__5_,s_r_124__4_,s_r_124__3_,s_r_124__2_,s_r_124__1_,
  s_r_124__0_,s_r_123__127_,s_r_123__126_,s_r_123__125_,s_r_123__124_,s_r_123__123_,
  s_r_123__122_,s_r_123__121_,s_r_123__120_,s_r_123__119_,s_r_123__118_,s_r_123__117_,
  s_r_123__116_,s_r_123__115_,s_r_123__114_,s_r_123__113_,s_r_123__112_,s_r_123__111_,
  s_r_123__110_,s_r_123__109_,s_r_123__108_,s_r_123__107_,s_r_123__106_,
  s_r_123__105_,s_r_123__104_,s_r_123__103_,s_r_123__102_,s_r_123__101_,s_r_123__100_,
  s_r_123__99_,s_r_123__98_,s_r_123__97_,s_r_123__96_,s_r_123__95_,s_r_123__94_,
  s_r_123__93_,s_r_123__92_,s_r_123__91_,s_r_123__90_,s_r_123__89_,s_r_123__88_,
  s_r_123__87_,s_r_123__86_,s_r_123__85_,s_r_123__84_,s_r_123__83_,s_r_123__82_,s_r_123__81_,
  s_r_123__80_,s_r_123__79_,s_r_123__78_,s_r_123__77_,s_r_123__76_,s_r_123__75_,
  s_r_123__74_,s_r_123__73_,s_r_123__72_,s_r_123__71_,s_r_123__70_,s_r_123__69_,
  s_r_123__68_,s_r_123__67_,s_r_123__66_,s_r_123__65_,s_r_123__64_,s_r_123__63_,
  s_r_123__62_,s_r_123__61_,s_r_123__60_,s_r_123__59_,s_r_123__58_,s_r_123__57_,
  s_r_123__56_,s_r_123__55_,s_r_123__54_,s_r_123__53_,s_r_123__52_,s_r_123__51_,
  s_r_123__50_,s_r_123__49_,s_r_123__48_,s_r_123__47_,s_r_123__46_,s_r_123__45_,
  s_r_123__44_,s_r_123__43_,s_r_123__42_,s_r_123__41_,s_r_123__40_,s_r_123__39_,s_r_123__38_,
  s_r_123__37_,s_r_123__36_,s_r_123__35_,s_r_123__34_,s_r_123__33_,s_r_123__32_,
  s_r_123__31_,s_r_123__30_,s_r_123__29_,s_r_123__28_,s_r_123__27_,s_r_123__26_,
  s_r_123__25_,s_r_123__24_,s_r_123__23_,s_r_123__22_,s_r_123__21_,s_r_123__20_,
  s_r_123__19_,s_r_123__18_,s_r_123__17_,s_r_123__16_,s_r_123__15_,s_r_123__14_,
  s_r_123__13_,s_r_123__12_,s_r_123__11_,s_r_123__10_,s_r_123__9_,s_r_123__8_,s_r_123__7_,
  s_r_123__6_,s_r_123__5_,s_r_123__4_,s_r_123__3_,s_r_123__2_,s_r_123__1_,
  s_r_123__0_,prod_accum_126__127_,prod_accum_125__126_,prod_accum_125__125_,
  prod_accum_125__124_,prod_accum_125__123_,prod_accum_125__122_,prod_accum_125__121_,
  prod_accum_125__120_,prod_accum_125__119_,prod_accum_125__118_,prod_accum_125__117_,
  prod_accum_125__116_,prod_accum_125__115_,prod_accum_125__114_,prod_accum_125__113_,
  prod_accum_125__112_,prod_accum_125__111_,prod_accum_125__110_,
  prod_accum_125__109_,prod_accum_125__108_,prod_accum_125__107_,prod_accum_125__106_,
  prod_accum_125__105_,prod_accum_125__104_,prod_accum_125__103_,prod_accum_125__102_,
  prod_accum_125__101_,prod_accum_125__100_,prod_accum_125__99_,prod_accum_125__98_,
  prod_accum_125__97_,prod_accum_125__96_,prod_accum_125__95_,prod_accum_125__94_,
  prod_accum_125__93_,prod_accum_125__92_,prod_accum_125__91_,prod_accum_125__90_,
  prod_accum_125__89_,prod_accum_125__88_,prod_accum_125__87_,prod_accum_125__86_,
  prod_accum_125__85_,prod_accum_125__84_,prod_accum_125__83_,prod_accum_125__82_,
  prod_accum_125__81_,prod_accum_125__80_,prod_accum_125__79_,prod_accum_125__78_,
  prod_accum_125__77_,prod_accum_125__76_,prod_accum_125__75_,prod_accum_125__74_,
  prod_accum_125__73_,prod_accum_125__72_,prod_accum_125__71_,prod_accum_125__70_,
  prod_accum_125__69_,prod_accum_125__68_,prod_accum_125__67_,prod_accum_125__66_,
  prod_accum_125__65_,prod_accum_125__64_,prod_accum_125__63_,prod_accum_125__62_,
  prod_accum_125__61_,prod_accum_125__60_,prod_accum_125__59_,prod_accum_125__58_,
  prod_accum_125__57_,prod_accum_125__56_,prod_accum_125__55_,prod_accum_125__54_,
  prod_accum_125__53_,prod_accum_125__52_,prod_accum_125__51_,prod_accum_125__50_,
  prod_accum_125__49_,prod_accum_125__48_,prod_accum_125__47_,prod_accum_125__46_,
  prod_accum_125__45_,prod_accum_125__44_,prod_accum_125__43_,prod_accum_125__42_,
  prod_accum_125__41_,prod_accum_125__40_,prod_accum_125__39_,prod_accum_125__38_,
  prod_accum_125__37_,prod_accum_125__36_,prod_accum_125__35_,prod_accum_125__34_,
  prod_accum_125__33_,prod_accum_125__32_,prod_accum_125__31_,prod_accum_125__30_,
  prod_accum_125__29_,prod_accum_125__28_,prod_accum_125__27_,prod_accum_125__26_,
  prod_accum_125__25_,prod_accum_125__24_,prod_accum_125__23_,prod_accum_125__22_,
  prod_accum_125__21_,prod_accum_125__20_,prod_accum_125__19_,prod_accum_125__18_,
  prod_accum_125__17_,prod_accum_125__16_,prod_accum_125__15_,prod_accum_125__14_,
  prod_accum_125__13_,prod_accum_125__12_,prod_accum_125__11_,prod_accum_125__10_,
  prod_accum_125__9_,prod_accum_125__8_,prod_accum_125__7_,prod_accum_125__6_,
  prod_accum_125__5_,prod_accum_125__4_,prod_accum_125__3_,prod_accum_125__2_,
  prod_accum_125__1_,prod_accum_125__0_,prod_accum_124__125_,prod_accum_124__124_,
  prod_accum_124__123_,prod_accum_124__122_,prod_accum_124__121_,prod_accum_124__120_,
  prod_accum_124__119_,prod_accum_124__118_,prod_accum_124__117_,prod_accum_124__116_,
  prod_accum_124__115_,prod_accum_124__114_,prod_accum_124__113_,prod_accum_124__112_,
  prod_accum_124__111_,prod_accum_124__110_,prod_accum_124__109_,prod_accum_124__108_,
  prod_accum_124__107_,prod_accum_124__106_,prod_accum_124__105_,
  prod_accum_124__104_,prod_accum_124__103_,prod_accum_124__102_,prod_accum_124__101_,
  prod_accum_124__100_,prod_accum_124__99_,prod_accum_124__98_,prod_accum_124__97_,
  prod_accum_124__96_,prod_accum_124__95_,prod_accum_124__94_,prod_accum_124__93_,
  prod_accum_124__92_,prod_accum_124__91_,prod_accum_124__90_,prod_accum_124__89_,
  prod_accum_124__88_,prod_accum_124__87_,prod_accum_124__86_,prod_accum_124__85_,
  prod_accum_124__84_,prod_accum_124__83_,prod_accum_124__82_,prod_accum_124__81_,
  prod_accum_124__80_,prod_accum_124__79_,prod_accum_124__78_,prod_accum_124__77_,
  prod_accum_124__76_,prod_accum_124__75_,prod_accum_124__74_,prod_accum_124__73_,
  prod_accum_124__72_,prod_accum_124__71_,prod_accum_124__70_,prod_accum_124__69_,
  prod_accum_124__68_,prod_accum_124__67_,prod_accum_124__66_,prod_accum_124__65_,
  prod_accum_124__64_,prod_accum_124__63_,prod_accum_124__62_,prod_accum_124__61_,
  prod_accum_124__60_,prod_accum_124__59_,prod_accum_124__58_,prod_accum_124__57_,
  prod_accum_124__56_,prod_accum_124__55_,prod_accum_124__54_,prod_accum_124__53_,
  prod_accum_124__52_,prod_accum_124__51_,prod_accum_124__50_,prod_accum_124__49_,
  prod_accum_124__48_,prod_accum_124__47_,prod_accum_124__46_,prod_accum_124__45_,
  prod_accum_124__44_,prod_accum_124__43_,prod_accum_124__42_,prod_accum_124__41_,
  prod_accum_124__40_,prod_accum_124__39_,prod_accum_124__38_,prod_accum_124__37_,
  prod_accum_124__36_,prod_accum_124__35_,prod_accum_124__34_,prod_accum_124__33_,
  prod_accum_124__32_,prod_accum_124__31_,prod_accum_124__30_,prod_accum_124__29_,
  prod_accum_124__28_,prod_accum_124__27_,prod_accum_124__26_,prod_accum_124__25_,
  prod_accum_124__24_,prod_accum_124__23_,prod_accum_124__22_,prod_accum_124__21_,
  prod_accum_124__20_,prod_accum_124__19_,prod_accum_124__18_,prod_accum_124__17_,
  prod_accum_124__16_,prod_accum_124__15_,prod_accum_124__14_,prod_accum_124__13_,
  prod_accum_124__12_,prod_accum_124__11_,prod_accum_124__10_,prod_accum_124__9_,
  prod_accum_124__8_,prod_accum_124__7_,prod_accum_124__6_,prod_accum_124__5_,
  prod_accum_124__4_,prod_accum_124__3_,prod_accum_124__2_,prod_accum_124__1_,prod_accum_124__0_,
  prod_accum_123__124_,prod_accum_123__123_,prod_accum_123__122_,
  prod_accum_123__121_,prod_accum_123__120_,prod_accum_123__119_,prod_accum_123__118_,
  prod_accum_123__117_,prod_accum_123__116_,prod_accum_123__115_,prod_accum_123__114_,
  prod_accum_123__113_,prod_accum_123__112_,prod_accum_123__111_,prod_accum_123__110_,
  prod_accum_123__109_,prod_accum_123__108_,prod_accum_123__107_,prod_accum_123__106_,
  prod_accum_123__105_,prod_accum_123__104_,prod_accum_123__103_,prod_accum_123__102_,
  prod_accum_123__101_,prod_accum_123__100_,prod_accum_123__99_,
  prod_accum_123__98_,prod_accum_123__97_,prod_accum_123__96_,prod_accum_123__95_,
  prod_accum_123__94_,prod_accum_123__93_,prod_accum_123__92_,prod_accum_123__91_,
  prod_accum_123__90_,prod_accum_123__89_,prod_accum_123__88_,prod_accum_123__87_,
  prod_accum_123__86_,prod_accum_123__85_,prod_accum_123__84_,prod_accum_123__83_,
  prod_accum_123__82_,prod_accum_123__81_,prod_accum_123__80_,prod_accum_123__79_,
  prod_accum_123__78_,prod_accum_123__77_,prod_accum_123__76_,prod_accum_123__75_,
  prod_accum_123__74_,prod_accum_123__73_,prod_accum_123__72_,prod_accum_123__71_,
  prod_accum_123__70_,prod_accum_123__69_,prod_accum_123__68_,prod_accum_123__67_,
  prod_accum_123__66_,prod_accum_123__65_,prod_accum_123__64_,prod_accum_123__63_,
  prod_accum_123__62_,prod_accum_123__61_,prod_accum_123__60_,prod_accum_123__59_,
  prod_accum_123__58_,prod_accum_123__57_,prod_accum_123__56_,prod_accum_123__55_,
  prod_accum_123__54_,prod_accum_123__53_,prod_accum_123__52_,prod_accum_123__51_,
  prod_accum_123__50_,prod_accum_123__49_,prod_accum_123__48_,prod_accum_123__47_,
  prod_accum_123__46_,prod_accum_123__45_,prod_accum_123__44_,prod_accum_123__43_,
  prod_accum_123__42_,prod_accum_123__41_,prod_accum_123__40_,prod_accum_123__39_,
  prod_accum_123__38_,prod_accum_123__37_,prod_accum_123__36_,prod_accum_123__35_,
  prod_accum_123__34_,prod_accum_123__33_,prod_accum_123__32_,prod_accum_123__31_,
  prod_accum_123__30_,prod_accum_123__29_,prod_accum_123__28_,prod_accum_123__27_,
  prod_accum_123__26_,prod_accum_123__25_,prod_accum_123__24_,prod_accum_123__23_,
  prod_accum_123__22_,prod_accum_123__21_,prod_accum_123__20_,prod_accum_123__19_,
  prod_accum_123__18_,prod_accum_123__17_,prod_accum_123__16_,prod_accum_123__15_,
  prod_accum_123__14_,prod_accum_123__13_,prod_accum_123__12_,prod_accum_123__11_,
  prod_accum_123__10_,prod_accum_123__9_,prod_accum_123__8_,prod_accum_123__7_,prod_accum_123__6_,
  prod_accum_123__5_,prod_accum_123__4_,prod_accum_123__3_,prod_accum_123__2_,
  prod_accum_123__1_,prod_accum_123__0_,SYNOPSYS_UNCONNECTED_1,SYNOPSYS_UNCONNECTED_2,
  SYNOPSYS_UNCONNECTED_3,SYNOPSYS_UNCONNECTED_4,SYNOPSYS_UNCONNECTED_5,
  SYNOPSYS_UNCONNECTED_6,SYNOPSYS_UNCONNECTED_7,SYNOPSYS_UNCONNECTED_8,SYNOPSYS_UNCONNECTED_9,
  SYNOPSYS_UNCONNECTED_10,SYNOPSYS_UNCONNECTED_11,SYNOPSYS_UNCONNECTED_12,
  SYNOPSYS_UNCONNECTED_13,SYNOPSYS_UNCONNECTED_14,SYNOPSYS_UNCONNECTED_15,
  SYNOPSYS_UNCONNECTED_16,SYNOPSYS_UNCONNECTED_17,SYNOPSYS_UNCONNECTED_18,SYNOPSYS_UNCONNECTED_19,
  SYNOPSYS_UNCONNECTED_20,SYNOPSYS_UNCONNECTED_21,SYNOPSYS_UNCONNECTED_22,
  SYNOPSYS_UNCONNECTED_23,SYNOPSYS_UNCONNECTED_24,SYNOPSYS_UNCONNECTED_25,
  SYNOPSYS_UNCONNECTED_26,SYNOPSYS_UNCONNECTED_27,SYNOPSYS_UNCONNECTED_28,SYNOPSYS_UNCONNECTED_29,
  SYNOPSYS_UNCONNECTED_30,SYNOPSYS_UNCONNECTED_31,SYNOPSYS_UNCONNECTED_32,
  SYNOPSYS_UNCONNECTED_33,SYNOPSYS_UNCONNECTED_34,SYNOPSYS_UNCONNECTED_35,
  SYNOPSYS_UNCONNECTED_36,SYNOPSYS_UNCONNECTED_37,SYNOPSYS_UNCONNECTED_38,SYNOPSYS_UNCONNECTED_39,
  SYNOPSYS_UNCONNECTED_40,SYNOPSYS_UNCONNECTED_41,SYNOPSYS_UNCONNECTED_42,
  SYNOPSYS_UNCONNECTED_43,SYNOPSYS_UNCONNECTED_44,SYNOPSYS_UNCONNECTED_45,
  SYNOPSYS_UNCONNECTED_46,SYNOPSYS_UNCONNECTED_47,SYNOPSYS_UNCONNECTED_48,SYNOPSYS_UNCONNECTED_49,
  SYNOPSYS_UNCONNECTED_50,SYNOPSYS_UNCONNECTED_51,SYNOPSYS_UNCONNECTED_52,
  SYNOPSYS_UNCONNECTED_53,SYNOPSYS_UNCONNECTED_54,SYNOPSYS_UNCONNECTED_55,
  SYNOPSYS_UNCONNECTED_56,SYNOPSYS_UNCONNECTED_57,SYNOPSYS_UNCONNECTED_58,SYNOPSYS_UNCONNECTED_59,
  SYNOPSYS_UNCONNECTED_60,SYNOPSYS_UNCONNECTED_61,SYNOPSYS_UNCONNECTED_62,
  SYNOPSYS_UNCONNECTED_63,SYNOPSYS_UNCONNECTED_64,SYNOPSYS_UNCONNECTED_65,
  SYNOPSYS_UNCONNECTED_66,SYNOPSYS_UNCONNECTED_67,SYNOPSYS_UNCONNECTED_68,SYNOPSYS_UNCONNECTED_69,
  SYNOPSYS_UNCONNECTED_70,SYNOPSYS_UNCONNECTED_71,SYNOPSYS_UNCONNECTED_72,
  SYNOPSYS_UNCONNECTED_73,SYNOPSYS_UNCONNECTED_74,SYNOPSYS_UNCONNECTED_75,
  SYNOPSYS_UNCONNECTED_76,SYNOPSYS_UNCONNECTED_77,SYNOPSYS_UNCONNECTED_78,SYNOPSYS_UNCONNECTED_79,
  SYNOPSYS_UNCONNECTED_80,SYNOPSYS_UNCONNECTED_81,SYNOPSYS_UNCONNECTED_82,
  SYNOPSYS_UNCONNECTED_83,SYNOPSYS_UNCONNECTED_84,SYNOPSYS_UNCONNECTED_85,
  SYNOPSYS_UNCONNECTED_86,SYNOPSYS_UNCONNECTED_87,SYNOPSYS_UNCONNECTED_88,SYNOPSYS_UNCONNECTED_89,
  SYNOPSYS_UNCONNECTED_90,SYNOPSYS_UNCONNECTED_91,SYNOPSYS_UNCONNECTED_92,
  SYNOPSYS_UNCONNECTED_93,SYNOPSYS_UNCONNECTED_94,SYNOPSYS_UNCONNECTED_95,
  SYNOPSYS_UNCONNECTED_96,SYNOPSYS_UNCONNECTED_97,SYNOPSYS_UNCONNECTED_98,SYNOPSYS_UNCONNECTED_99,
  SYNOPSYS_UNCONNECTED_100,SYNOPSYS_UNCONNECTED_101,SYNOPSYS_UNCONNECTED_102,
  SYNOPSYS_UNCONNECTED_103,SYNOPSYS_UNCONNECTED_104,SYNOPSYS_UNCONNECTED_105,
  SYNOPSYS_UNCONNECTED_106,SYNOPSYS_UNCONNECTED_107,SYNOPSYS_UNCONNECTED_108,
  SYNOPSYS_UNCONNECTED_109,SYNOPSYS_UNCONNECTED_110,SYNOPSYS_UNCONNECTED_111,
  SYNOPSYS_UNCONNECTED_112,SYNOPSYS_UNCONNECTED_113,SYNOPSYS_UNCONNECTED_114,SYNOPSYS_UNCONNECTED_115,
  SYNOPSYS_UNCONNECTED_116,SYNOPSYS_UNCONNECTED_117,SYNOPSYS_UNCONNECTED_118,
  SYNOPSYS_UNCONNECTED_119,SYNOPSYS_UNCONNECTED_120,SYNOPSYS_UNCONNECTED_121,
  SYNOPSYS_UNCONNECTED_122,SYNOPSYS_UNCONNECTED_123,SYNOPSYS_UNCONNECTED_124,
  SYNOPSYS_UNCONNECTED_125,SYNOPSYS_UNCONNECTED_126,SYNOPSYS_UNCONNECTED_127,
  SYNOPSYS_UNCONNECTED_128,SYNOPSYS_UNCONNECTED_129,SYNOPSYS_UNCONNECTED_130,SYNOPSYS_UNCONNECTED_131,
  SYNOPSYS_UNCONNECTED_132,SYNOPSYS_UNCONNECTED_133,SYNOPSYS_UNCONNECTED_134,
  SYNOPSYS_UNCONNECTED_135,SYNOPSYS_UNCONNECTED_136,SYNOPSYS_UNCONNECTED_137,
  SYNOPSYS_UNCONNECTED_138,SYNOPSYS_UNCONNECTED_139,SYNOPSYS_UNCONNECTED_140,
  SYNOPSYS_UNCONNECTED_141,SYNOPSYS_UNCONNECTED_142,SYNOPSYS_UNCONNECTED_143,
  SYNOPSYS_UNCONNECTED_144,SYNOPSYS_UNCONNECTED_145,SYNOPSYS_UNCONNECTED_146,SYNOPSYS_UNCONNECTED_147,
  SYNOPSYS_UNCONNECTED_148,SYNOPSYS_UNCONNECTED_149,SYNOPSYS_UNCONNECTED_150,
  SYNOPSYS_UNCONNECTED_151,SYNOPSYS_UNCONNECTED_152,SYNOPSYS_UNCONNECTED_153,
  SYNOPSYS_UNCONNECTED_154,SYNOPSYS_UNCONNECTED_155,SYNOPSYS_UNCONNECTED_156,
  SYNOPSYS_UNCONNECTED_157,SYNOPSYS_UNCONNECTED_158,SYNOPSYS_UNCONNECTED_159,
  SYNOPSYS_UNCONNECTED_160,SYNOPSYS_UNCONNECTED_161,SYNOPSYS_UNCONNECTED_162,SYNOPSYS_UNCONNECTED_163,
  SYNOPSYS_UNCONNECTED_164,SYNOPSYS_UNCONNECTED_165,SYNOPSYS_UNCONNECTED_166,
  SYNOPSYS_UNCONNECTED_167,SYNOPSYS_UNCONNECTED_168,SYNOPSYS_UNCONNECTED_169,
  SYNOPSYS_UNCONNECTED_170,SYNOPSYS_UNCONNECTED_171,SYNOPSYS_UNCONNECTED_172,
  SYNOPSYS_UNCONNECTED_173,SYNOPSYS_UNCONNECTED_174,SYNOPSYS_UNCONNECTED_175,
  SYNOPSYS_UNCONNECTED_176,SYNOPSYS_UNCONNECTED_177,SYNOPSYS_UNCONNECTED_178,SYNOPSYS_UNCONNECTED_179,
  SYNOPSYS_UNCONNECTED_180,SYNOPSYS_UNCONNECTED_181,SYNOPSYS_UNCONNECTED_182,
  SYNOPSYS_UNCONNECTED_183,SYNOPSYS_UNCONNECTED_184,SYNOPSYS_UNCONNECTED_185,
  SYNOPSYS_UNCONNECTED_186,SYNOPSYS_UNCONNECTED_187,SYNOPSYS_UNCONNECTED_188,
  SYNOPSYS_UNCONNECTED_189,SYNOPSYS_UNCONNECTED_190,SYNOPSYS_UNCONNECTED_191,
  SYNOPSYS_UNCONNECTED_192,SYNOPSYS_UNCONNECTED_193,SYNOPSYS_UNCONNECTED_194,SYNOPSYS_UNCONNECTED_195,
  SYNOPSYS_UNCONNECTED_196,SYNOPSYS_UNCONNECTED_197,SYNOPSYS_UNCONNECTED_198,
  SYNOPSYS_UNCONNECTED_199,SYNOPSYS_UNCONNECTED_200,SYNOPSYS_UNCONNECTED_201,
  SYNOPSYS_UNCONNECTED_202,SYNOPSYS_UNCONNECTED_203,SYNOPSYS_UNCONNECTED_204,
  SYNOPSYS_UNCONNECTED_205,SYNOPSYS_UNCONNECTED_206,SYNOPSYS_UNCONNECTED_207,
  SYNOPSYS_UNCONNECTED_208,SYNOPSYS_UNCONNECTED_209,SYNOPSYS_UNCONNECTED_210,SYNOPSYS_UNCONNECTED_211,
  SYNOPSYS_UNCONNECTED_212,SYNOPSYS_UNCONNECTED_213,SYNOPSYS_UNCONNECTED_214,
  SYNOPSYS_UNCONNECTED_215,SYNOPSYS_UNCONNECTED_216,SYNOPSYS_UNCONNECTED_217,
  SYNOPSYS_UNCONNECTED_218,SYNOPSYS_UNCONNECTED_219,SYNOPSYS_UNCONNECTED_220,
  SYNOPSYS_UNCONNECTED_221,SYNOPSYS_UNCONNECTED_222,SYNOPSYS_UNCONNECTED_223,
  SYNOPSYS_UNCONNECTED_224,SYNOPSYS_UNCONNECTED_225,SYNOPSYS_UNCONNECTED_226,SYNOPSYS_UNCONNECTED_227,
  SYNOPSYS_UNCONNECTED_228,SYNOPSYS_UNCONNECTED_229,SYNOPSYS_UNCONNECTED_230,
  SYNOPSYS_UNCONNECTED_231,SYNOPSYS_UNCONNECTED_232,SYNOPSYS_UNCONNECTED_233,
  SYNOPSYS_UNCONNECTED_234,SYNOPSYS_UNCONNECTED_235,SYNOPSYS_UNCONNECTED_236,
  SYNOPSYS_UNCONNECTED_237,SYNOPSYS_UNCONNECTED_238,SYNOPSYS_UNCONNECTED_239,
  SYNOPSYS_UNCONNECTED_240,SYNOPSYS_UNCONNECTED_241,SYNOPSYS_UNCONNECTED_242,SYNOPSYS_UNCONNECTED_243,
  SYNOPSYS_UNCONNECTED_244,SYNOPSYS_UNCONNECTED_245,SYNOPSYS_UNCONNECTED_246,
  SYNOPSYS_UNCONNECTED_247,SYNOPSYS_UNCONNECTED_248,SYNOPSYS_UNCONNECTED_249,
  SYNOPSYS_UNCONNECTED_250,SYNOPSYS_UNCONNECTED_251,SYNOPSYS_UNCONNECTED_252,
  SYNOPSYS_UNCONNECTED_253,SYNOPSYS_UNCONNECTED_254,SYNOPSYS_UNCONNECTED_255,
  SYNOPSYS_UNCONNECTED_256;
  wire [127:0] pp0;
  wire [16127:0] a_r,b_r;
  wire [125:0] c_r;

  bsg_and_width_p128
  and0
  (
    .a_i(a_i),
    .b_i({ b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0], b_i[0:0] }),
    .o(pp0)
  );


  bsg_mul_array_row_128_0_0
  genblk1_0__genblk1_first_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_i),
    .b_i(b_i),
    .s_i(pp0),
    .c_i(1'b0),
    .prod_accum_i(pp0[0]),
    .a_o(a_r[127:0]),
    .b_o(b_r[127:0]),
    .s_o({ s_r_0__127_, s_r_0__126_, s_r_0__125_, s_r_0__124_, s_r_0__123_, s_r_0__122_, s_r_0__121_, s_r_0__120_, s_r_0__119_, s_r_0__118_, s_r_0__117_, s_r_0__116_, s_r_0__115_, s_r_0__114_, s_r_0__113_, s_r_0__112_, s_r_0__111_, s_r_0__110_, s_r_0__109_, s_r_0__108_, s_r_0__107_, s_r_0__106_, s_r_0__105_, s_r_0__104_, s_r_0__103_, s_r_0__102_, s_r_0__101_, s_r_0__100_, s_r_0__99_, s_r_0__98_, s_r_0__97_, s_r_0__96_, s_r_0__95_, s_r_0__94_, s_r_0__93_, s_r_0__92_, s_r_0__91_, s_r_0__90_, s_r_0__89_, s_r_0__88_, s_r_0__87_, s_r_0__86_, s_r_0__85_, s_r_0__84_, s_r_0__83_, s_r_0__82_, s_r_0__81_, s_r_0__80_, s_r_0__79_, s_r_0__78_, s_r_0__77_, s_r_0__76_, s_r_0__75_, s_r_0__74_, s_r_0__73_, s_r_0__72_, s_r_0__71_, s_r_0__70_, s_r_0__69_, s_r_0__68_, s_r_0__67_, s_r_0__66_, s_r_0__65_, s_r_0__64_, s_r_0__63_, s_r_0__62_, s_r_0__61_, s_r_0__60_, s_r_0__59_, s_r_0__58_, s_r_0__57_, s_r_0__56_, s_r_0__55_, s_r_0__54_, s_r_0__53_, s_r_0__52_, s_r_0__51_, s_r_0__50_, s_r_0__49_, s_r_0__48_, s_r_0__47_, s_r_0__46_, s_r_0__45_, s_r_0__44_, s_r_0__43_, s_r_0__42_, s_r_0__41_, s_r_0__40_, s_r_0__39_, s_r_0__38_, s_r_0__37_, s_r_0__36_, s_r_0__35_, s_r_0__34_, s_r_0__33_, s_r_0__32_, s_r_0__31_, s_r_0__30_, s_r_0__29_, s_r_0__28_, s_r_0__27_, s_r_0__26_, s_r_0__25_, s_r_0__24_, s_r_0__23_, s_r_0__22_, s_r_0__21_, s_r_0__20_, s_r_0__19_, s_r_0__18_, s_r_0__17_, s_r_0__16_, s_r_0__15_, s_r_0__14_, s_r_0__13_, s_r_0__12_, s_r_0__11_, s_r_0__10_, s_r_0__9_, s_r_0__8_, s_r_0__7_, s_r_0__6_, s_r_0__5_, s_r_0__4_, s_r_0__3_, s_r_0__2_, s_r_0__1_, s_r_0__0_ }),
    .c_o(c_r[0]),
    .prod_accum_o({ prod_accum_0__1_, prod_accum_0__0_ })
  );


  bsg_mul_array_row_128_1_0
  genblk1_1__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[127:0]),
    .b_i(b_r[127:0]),
    .s_i({ s_r_0__127_, s_r_0__126_, s_r_0__125_, s_r_0__124_, s_r_0__123_, s_r_0__122_, s_r_0__121_, s_r_0__120_, s_r_0__119_, s_r_0__118_, s_r_0__117_, s_r_0__116_, s_r_0__115_, s_r_0__114_, s_r_0__113_, s_r_0__112_, s_r_0__111_, s_r_0__110_, s_r_0__109_, s_r_0__108_, s_r_0__107_, s_r_0__106_, s_r_0__105_, s_r_0__104_, s_r_0__103_, s_r_0__102_, s_r_0__101_, s_r_0__100_, s_r_0__99_, s_r_0__98_, s_r_0__97_, s_r_0__96_, s_r_0__95_, s_r_0__94_, s_r_0__93_, s_r_0__92_, s_r_0__91_, s_r_0__90_, s_r_0__89_, s_r_0__88_, s_r_0__87_, s_r_0__86_, s_r_0__85_, s_r_0__84_, s_r_0__83_, s_r_0__82_, s_r_0__81_, s_r_0__80_, s_r_0__79_, s_r_0__78_, s_r_0__77_, s_r_0__76_, s_r_0__75_, s_r_0__74_, s_r_0__73_, s_r_0__72_, s_r_0__71_, s_r_0__70_, s_r_0__69_, s_r_0__68_, s_r_0__67_, s_r_0__66_, s_r_0__65_, s_r_0__64_, s_r_0__63_, s_r_0__62_, s_r_0__61_, s_r_0__60_, s_r_0__59_, s_r_0__58_, s_r_0__57_, s_r_0__56_, s_r_0__55_, s_r_0__54_, s_r_0__53_, s_r_0__52_, s_r_0__51_, s_r_0__50_, s_r_0__49_, s_r_0__48_, s_r_0__47_, s_r_0__46_, s_r_0__45_, s_r_0__44_, s_r_0__43_, s_r_0__42_, s_r_0__41_, s_r_0__40_, s_r_0__39_, s_r_0__38_, s_r_0__37_, s_r_0__36_, s_r_0__35_, s_r_0__34_, s_r_0__33_, s_r_0__32_, s_r_0__31_, s_r_0__30_, s_r_0__29_, s_r_0__28_, s_r_0__27_, s_r_0__26_, s_r_0__25_, s_r_0__24_, s_r_0__23_, s_r_0__22_, s_r_0__21_, s_r_0__20_, s_r_0__19_, s_r_0__18_, s_r_0__17_, s_r_0__16_, s_r_0__15_, s_r_0__14_, s_r_0__13_, s_r_0__12_, s_r_0__11_, s_r_0__10_, s_r_0__9_, s_r_0__8_, s_r_0__7_, s_r_0__6_, s_r_0__5_, s_r_0__4_, s_r_0__3_, s_r_0__2_, s_r_0__1_, s_r_0__0_ }),
    .c_i(c_r[0]),
    .prod_accum_i({ prod_accum_0__1_, prod_accum_0__0_ }),
    .a_o(a_r[255:128]),
    .b_o(b_r[255:128]),
    .s_o({ s_r_1__127_, s_r_1__126_, s_r_1__125_, s_r_1__124_, s_r_1__123_, s_r_1__122_, s_r_1__121_, s_r_1__120_, s_r_1__119_, s_r_1__118_, s_r_1__117_, s_r_1__116_, s_r_1__115_, s_r_1__114_, s_r_1__113_, s_r_1__112_, s_r_1__111_, s_r_1__110_, s_r_1__109_, s_r_1__108_, s_r_1__107_, s_r_1__106_, s_r_1__105_, s_r_1__104_, s_r_1__103_, s_r_1__102_, s_r_1__101_, s_r_1__100_, s_r_1__99_, s_r_1__98_, s_r_1__97_, s_r_1__96_, s_r_1__95_, s_r_1__94_, s_r_1__93_, s_r_1__92_, s_r_1__91_, s_r_1__90_, s_r_1__89_, s_r_1__88_, s_r_1__87_, s_r_1__86_, s_r_1__85_, s_r_1__84_, s_r_1__83_, s_r_1__82_, s_r_1__81_, s_r_1__80_, s_r_1__79_, s_r_1__78_, s_r_1__77_, s_r_1__76_, s_r_1__75_, s_r_1__74_, s_r_1__73_, s_r_1__72_, s_r_1__71_, s_r_1__70_, s_r_1__69_, s_r_1__68_, s_r_1__67_, s_r_1__66_, s_r_1__65_, s_r_1__64_, s_r_1__63_, s_r_1__62_, s_r_1__61_, s_r_1__60_, s_r_1__59_, s_r_1__58_, s_r_1__57_, s_r_1__56_, s_r_1__55_, s_r_1__54_, s_r_1__53_, s_r_1__52_, s_r_1__51_, s_r_1__50_, s_r_1__49_, s_r_1__48_, s_r_1__47_, s_r_1__46_, s_r_1__45_, s_r_1__44_, s_r_1__43_, s_r_1__42_, s_r_1__41_, s_r_1__40_, s_r_1__39_, s_r_1__38_, s_r_1__37_, s_r_1__36_, s_r_1__35_, s_r_1__34_, s_r_1__33_, s_r_1__32_, s_r_1__31_, s_r_1__30_, s_r_1__29_, s_r_1__28_, s_r_1__27_, s_r_1__26_, s_r_1__25_, s_r_1__24_, s_r_1__23_, s_r_1__22_, s_r_1__21_, s_r_1__20_, s_r_1__19_, s_r_1__18_, s_r_1__17_, s_r_1__16_, s_r_1__15_, s_r_1__14_, s_r_1__13_, s_r_1__12_, s_r_1__11_, s_r_1__10_, s_r_1__9_, s_r_1__8_, s_r_1__7_, s_r_1__6_, s_r_1__5_, s_r_1__4_, s_r_1__3_, s_r_1__2_, s_r_1__1_, s_r_1__0_ }),
    .c_o(c_r[1]),
    .prod_accum_o({ prod_accum_1__2_, prod_accum_1__1_, prod_accum_1__0_ })
  );


  bsg_mul_array_row_128_2_0
  genblk1_2__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[255:128]),
    .b_i(b_r[255:128]),
    .s_i({ s_r_1__127_, s_r_1__126_, s_r_1__125_, s_r_1__124_, s_r_1__123_, s_r_1__122_, s_r_1__121_, s_r_1__120_, s_r_1__119_, s_r_1__118_, s_r_1__117_, s_r_1__116_, s_r_1__115_, s_r_1__114_, s_r_1__113_, s_r_1__112_, s_r_1__111_, s_r_1__110_, s_r_1__109_, s_r_1__108_, s_r_1__107_, s_r_1__106_, s_r_1__105_, s_r_1__104_, s_r_1__103_, s_r_1__102_, s_r_1__101_, s_r_1__100_, s_r_1__99_, s_r_1__98_, s_r_1__97_, s_r_1__96_, s_r_1__95_, s_r_1__94_, s_r_1__93_, s_r_1__92_, s_r_1__91_, s_r_1__90_, s_r_1__89_, s_r_1__88_, s_r_1__87_, s_r_1__86_, s_r_1__85_, s_r_1__84_, s_r_1__83_, s_r_1__82_, s_r_1__81_, s_r_1__80_, s_r_1__79_, s_r_1__78_, s_r_1__77_, s_r_1__76_, s_r_1__75_, s_r_1__74_, s_r_1__73_, s_r_1__72_, s_r_1__71_, s_r_1__70_, s_r_1__69_, s_r_1__68_, s_r_1__67_, s_r_1__66_, s_r_1__65_, s_r_1__64_, s_r_1__63_, s_r_1__62_, s_r_1__61_, s_r_1__60_, s_r_1__59_, s_r_1__58_, s_r_1__57_, s_r_1__56_, s_r_1__55_, s_r_1__54_, s_r_1__53_, s_r_1__52_, s_r_1__51_, s_r_1__50_, s_r_1__49_, s_r_1__48_, s_r_1__47_, s_r_1__46_, s_r_1__45_, s_r_1__44_, s_r_1__43_, s_r_1__42_, s_r_1__41_, s_r_1__40_, s_r_1__39_, s_r_1__38_, s_r_1__37_, s_r_1__36_, s_r_1__35_, s_r_1__34_, s_r_1__33_, s_r_1__32_, s_r_1__31_, s_r_1__30_, s_r_1__29_, s_r_1__28_, s_r_1__27_, s_r_1__26_, s_r_1__25_, s_r_1__24_, s_r_1__23_, s_r_1__22_, s_r_1__21_, s_r_1__20_, s_r_1__19_, s_r_1__18_, s_r_1__17_, s_r_1__16_, s_r_1__15_, s_r_1__14_, s_r_1__13_, s_r_1__12_, s_r_1__11_, s_r_1__10_, s_r_1__9_, s_r_1__8_, s_r_1__7_, s_r_1__6_, s_r_1__5_, s_r_1__4_, s_r_1__3_, s_r_1__2_, s_r_1__1_, s_r_1__0_ }),
    .c_i(c_r[1]),
    .prod_accum_i({ prod_accum_1__2_, prod_accum_1__1_, prod_accum_1__0_ }),
    .a_o(a_r[383:256]),
    .b_o(b_r[383:256]),
    .s_o({ s_r_2__127_, s_r_2__126_, s_r_2__125_, s_r_2__124_, s_r_2__123_, s_r_2__122_, s_r_2__121_, s_r_2__120_, s_r_2__119_, s_r_2__118_, s_r_2__117_, s_r_2__116_, s_r_2__115_, s_r_2__114_, s_r_2__113_, s_r_2__112_, s_r_2__111_, s_r_2__110_, s_r_2__109_, s_r_2__108_, s_r_2__107_, s_r_2__106_, s_r_2__105_, s_r_2__104_, s_r_2__103_, s_r_2__102_, s_r_2__101_, s_r_2__100_, s_r_2__99_, s_r_2__98_, s_r_2__97_, s_r_2__96_, s_r_2__95_, s_r_2__94_, s_r_2__93_, s_r_2__92_, s_r_2__91_, s_r_2__90_, s_r_2__89_, s_r_2__88_, s_r_2__87_, s_r_2__86_, s_r_2__85_, s_r_2__84_, s_r_2__83_, s_r_2__82_, s_r_2__81_, s_r_2__80_, s_r_2__79_, s_r_2__78_, s_r_2__77_, s_r_2__76_, s_r_2__75_, s_r_2__74_, s_r_2__73_, s_r_2__72_, s_r_2__71_, s_r_2__70_, s_r_2__69_, s_r_2__68_, s_r_2__67_, s_r_2__66_, s_r_2__65_, s_r_2__64_, s_r_2__63_, s_r_2__62_, s_r_2__61_, s_r_2__60_, s_r_2__59_, s_r_2__58_, s_r_2__57_, s_r_2__56_, s_r_2__55_, s_r_2__54_, s_r_2__53_, s_r_2__52_, s_r_2__51_, s_r_2__50_, s_r_2__49_, s_r_2__48_, s_r_2__47_, s_r_2__46_, s_r_2__45_, s_r_2__44_, s_r_2__43_, s_r_2__42_, s_r_2__41_, s_r_2__40_, s_r_2__39_, s_r_2__38_, s_r_2__37_, s_r_2__36_, s_r_2__35_, s_r_2__34_, s_r_2__33_, s_r_2__32_, s_r_2__31_, s_r_2__30_, s_r_2__29_, s_r_2__28_, s_r_2__27_, s_r_2__26_, s_r_2__25_, s_r_2__24_, s_r_2__23_, s_r_2__22_, s_r_2__21_, s_r_2__20_, s_r_2__19_, s_r_2__18_, s_r_2__17_, s_r_2__16_, s_r_2__15_, s_r_2__14_, s_r_2__13_, s_r_2__12_, s_r_2__11_, s_r_2__10_, s_r_2__9_, s_r_2__8_, s_r_2__7_, s_r_2__6_, s_r_2__5_, s_r_2__4_, s_r_2__3_, s_r_2__2_, s_r_2__1_, s_r_2__0_ }),
    .c_o(c_r[2]),
    .prod_accum_o({ prod_accum_2__3_, prod_accum_2__2_, prod_accum_2__1_, prod_accum_2__0_ })
  );


  bsg_mul_array_row_128_3_0
  genblk1_3__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[383:256]),
    .b_i(b_r[383:256]),
    .s_i({ s_r_2__127_, s_r_2__126_, s_r_2__125_, s_r_2__124_, s_r_2__123_, s_r_2__122_, s_r_2__121_, s_r_2__120_, s_r_2__119_, s_r_2__118_, s_r_2__117_, s_r_2__116_, s_r_2__115_, s_r_2__114_, s_r_2__113_, s_r_2__112_, s_r_2__111_, s_r_2__110_, s_r_2__109_, s_r_2__108_, s_r_2__107_, s_r_2__106_, s_r_2__105_, s_r_2__104_, s_r_2__103_, s_r_2__102_, s_r_2__101_, s_r_2__100_, s_r_2__99_, s_r_2__98_, s_r_2__97_, s_r_2__96_, s_r_2__95_, s_r_2__94_, s_r_2__93_, s_r_2__92_, s_r_2__91_, s_r_2__90_, s_r_2__89_, s_r_2__88_, s_r_2__87_, s_r_2__86_, s_r_2__85_, s_r_2__84_, s_r_2__83_, s_r_2__82_, s_r_2__81_, s_r_2__80_, s_r_2__79_, s_r_2__78_, s_r_2__77_, s_r_2__76_, s_r_2__75_, s_r_2__74_, s_r_2__73_, s_r_2__72_, s_r_2__71_, s_r_2__70_, s_r_2__69_, s_r_2__68_, s_r_2__67_, s_r_2__66_, s_r_2__65_, s_r_2__64_, s_r_2__63_, s_r_2__62_, s_r_2__61_, s_r_2__60_, s_r_2__59_, s_r_2__58_, s_r_2__57_, s_r_2__56_, s_r_2__55_, s_r_2__54_, s_r_2__53_, s_r_2__52_, s_r_2__51_, s_r_2__50_, s_r_2__49_, s_r_2__48_, s_r_2__47_, s_r_2__46_, s_r_2__45_, s_r_2__44_, s_r_2__43_, s_r_2__42_, s_r_2__41_, s_r_2__40_, s_r_2__39_, s_r_2__38_, s_r_2__37_, s_r_2__36_, s_r_2__35_, s_r_2__34_, s_r_2__33_, s_r_2__32_, s_r_2__31_, s_r_2__30_, s_r_2__29_, s_r_2__28_, s_r_2__27_, s_r_2__26_, s_r_2__25_, s_r_2__24_, s_r_2__23_, s_r_2__22_, s_r_2__21_, s_r_2__20_, s_r_2__19_, s_r_2__18_, s_r_2__17_, s_r_2__16_, s_r_2__15_, s_r_2__14_, s_r_2__13_, s_r_2__12_, s_r_2__11_, s_r_2__10_, s_r_2__9_, s_r_2__8_, s_r_2__7_, s_r_2__6_, s_r_2__5_, s_r_2__4_, s_r_2__3_, s_r_2__2_, s_r_2__1_, s_r_2__0_ }),
    .c_i(c_r[2]),
    .prod_accum_i({ prod_accum_2__3_, prod_accum_2__2_, prod_accum_2__1_, prod_accum_2__0_ }),
    .a_o(a_r[511:384]),
    .b_o(b_r[511:384]),
    .s_o({ s_r_3__127_, s_r_3__126_, s_r_3__125_, s_r_3__124_, s_r_3__123_, s_r_3__122_, s_r_3__121_, s_r_3__120_, s_r_3__119_, s_r_3__118_, s_r_3__117_, s_r_3__116_, s_r_3__115_, s_r_3__114_, s_r_3__113_, s_r_3__112_, s_r_3__111_, s_r_3__110_, s_r_3__109_, s_r_3__108_, s_r_3__107_, s_r_3__106_, s_r_3__105_, s_r_3__104_, s_r_3__103_, s_r_3__102_, s_r_3__101_, s_r_3__100_, s_r_3__99_, s_r_3__98_, s_r_3__97_, s_r_3__96_, s_r_3__95_, s_r_3__94_, s_r_3__93_, s_r_3__92_, s_r_3__91_, s_r_3__90_, s_r_3__89_, s_r_3__88_, s_r_3__87_, s_r_3__86_, s_r_3__85_, s_r_3__84_, s_r_3__83_, s_r_3__82_, s_r_3__81_, s_r_3__80_, s_r_3__79_, s_r_3__78_, s_r_3__77_, s_r_3__76_, s_r_3__75_, s_r_3__74_, s_r_3__73_, s_r_3__72_, s_r_3__71_, s_r_3__70_, s_r_3__69_, s_r_3__68_, s_r_3__67_, s_r_3__66_, s_r_3__65_, s_r_3__64_, s_r_3__63_, s_r_3__62_, s_r_3__61_, s_r_3__60_, s_r_3__59_, s_r_3__58_, s_r_3__57_, s_r_3__56_, s_r_3__55_, s_r_3__54_, s_r_3__53_, s_r_3__52_, s_r_3__51_, s_r_3__50_, s_r_3__49_, s_r_3__48_, s_r_3__47_, s_r_3__46_, s_r_3__45_, s_r_3__44_, s_r_3__43_, s_r_3__42_, s_r_3__41_, s_r_3__40_, s_r_3__39_, s_r_3__38_, s_r_3__37_, s_r_3__36_, s_r_3__35_, s_r_3__34_, s_r_3__33_, s_r_3__32_, s_r_3__31_, s_r_3__30_, s_r_3__29_, s_r_3__28_, s_r_3__27_, s_r_3__26_, s_r_3__25_, s_r_3__24_, s_r_3__23_, s_r_3__22_, s_r_3__21_, s_r_3__20_, s_r_3__19_, s_r_3__18_, s_r_3__17_, s_r_3__16_, s_r_3__15_, s_r_3__14_, s_r_3__13_, s_r_3__12_, s_r_3__11_, s_r_3__10_, s_r_3__9_, s_r_3__8_, s_r_3__7_, s_r_3__6_, s_r_3__5_, s_r_3__4_, s_r_3__3_, s_r_3__2_, s_r_3__1_, s_r_3__0_ }),
    .c_o(c_r[3]),
    .prod_accum_o({ prod_accum_3__4_, prod_accum_3__3_, prod_accum_3__2_, prod_accum_3__1_, prod_accum_3__0_ })
  );


  bsg_mul_array_row_128_4_0
  genblk1_4__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[511:384]),
    .b_i(b_r[511:384]),
    .s_i({ s_r_3__127_, s_r_3__126_, s_r_3__125_, s_r_3__124_, s_r_3__123_, s_r_3__122_, s_r_3__121_, s_r_3__120_, s_r_3__119_, s_r_3__118_, s_r_3__117_, s_r_3__116_, s_r_3__115_, s_r_3__114_, s_r_3__113_, s_r_3__112_, s_r_3__111_, s_r_3__110_, s_r_3__109_, s_r_3__108_, s_r_3__107_, s_r_3__106_, s_r_3__105_, s_r_3__104_, s_r_3__103_, s_r_3__102_, s_r_3__101_, s_r_3__100_, s_r_3__99_, s_r_3__98_, s_r_3__97_, s_r_3__96_, s_r_3__95_, s_r_3__94_, s_r_3__93_, s_r_3__92_, s_r_3__91_, s_r_3__90_, s_r_3__89_, s_r_3__88_, s_r_3__87_, s_r_3__86_, s_r_3__85_, s_r_3__84_, s_r_3__83_, s_r_3__82_, s_r_3__81_, s_r_3__80_, s_r_3__79_, s_r_3__78_, s_r_3__77_, s_r_3__76_, s_r_3__75_, s_r_3__74_, s_r_3__73_, s_r_3__72_, s_r_3__71_, s_r_3__70_, s_r_3__69_, s_r_3__68_, s_r_3__67_, s_r_3__66_, s_r_3__65_, s_r_3__64_, s_r_3__63_, s_r_3__62_, s_r_3__61_, s_r_3__60_, s_r_3__59_, s_r_3__58_, s_r_3__57_, s_r_3__56_, s_r_3__55_, s_r_3__54_, s_r_3__53_, s_r_3__52_, s_r_3__51_, s_r_3__50_, s_r_3__49_, s_r_3__48_, s_r_3__47_, s_r_3__46_, s_r_3__45_, s_r_3__44_, s_r_3__43_, s_r_3__42_, s_r_3__41_, s_r_3__40_, s_r_3__39_, s_r_3__38_, s_r_3__37_, s_r_3__36_, s_r_3__35_, s_r_3__34_, s_r_3__33_, s_r_3__32_, s_r_3__31_, s_r_3__30_, s_r_3__29_, s_r_3__28_, s_r_3__27_, s_r_3__26_, s_r_3__25_, s_r_3__24_, s_r_3__23_, s_r_3__22_, s_r_3__21_, s_r_3__20_, s_r_3__19_, s_r_3__18_, s_r_3__17_, s_r_3__16_, s_r_3__15_, s_r_3__14_, s_r_3__13_, s_r_3__12_, s_r_3__11_, s_r_3__10_, s_r_3__9_, s_r_3__8_, s_r_3__7_, s_r_3__6_, s_r_3__5_, s_r_3__4_, s_r_3__3_, s_r_3__2_, s_r_3__1_, s_r_3__0_ }),
    .c_i(c_r[3]),
    .prod_accum_i({ prod_accum_3__4_, prod_accum_3__3_, prod_accum_3__2_, prod_accum_3__1_, prod_accum_3__0_ }),
    .a_o(a_r[639:512]),
    .b_o(b_r[639:512]),
    .s_o({ s_r_4__127_, s_r_4__126_, s_r_4__125_, s_r_4__124_, s_r_4__123_, s_r_4__122_, s_r_4__121_, s_r_4__120_, s_r_4__119_, s_r_4__118_, s_r_4__117_, s_r_4__116_, s_r_4__115_, s_r_4__114_, s_r_4__113_, s_r_4__112_, s_r_4__111_, s_r_4__110_, s_r_4__109_, s_r_4__108_, s_r_4__107_, s_r_4__106_, s_r_4__105_, s_r_4__104_, s_r_4__103_, s_r_4__102_, s_r_4__101_, s_r_4__100_, s_r_4__99_, s_r_4__98_, s_r_4__97_, s_r_4__96_, s_r_4__95_, s_r_4__94_, s_r_4__93_, s_r_4__92_, s_r_4__91_, s_r_4__90_, s_r_4__89_, s_r_4__88_, s_r_4__87_, s_r_4__86_, s_r_4__85_, s_r_4__84_, s_r_4__83_, s_r_4__82_, s_r_4__81_, s_r_4__80_, s_r_4__79_, s_r_4__78_, s_r_4__77_, s_r_4__76_, s_r_4__75_, s_r_4__74_, s_r_4__73_, s_r_4__72_, s_r_4__71_, s_r_4__70_, s_r_4__69_, s_r_4__68_, s_r_4__67_, s_r_4__66_, s_r_4__65_, s_r_4__64_, s_r_4__63_, s_r_4__62_, s_r_4__61_, s_r_4__60_, s_r_4__59_, s_r_4__58_, s_r_4__57_, s_r_4__56_, s_r_4__55_, s_r_4__54_, s_r_4__53_, s_r_4__52_, s_r_4__51_, s_r_4__50_, s_r_4__49_, s_r_4__48_, s_r_4__47_, s_r_4__46_, s_r_4__45_, s_r_4__44_, s_r_4__43_, s_r_4__42_, s_r_4__41_, s_r_4__40_, s_r_4__39_, s_r_4__38_, s_r_4__37_, s_r_4__36_, s_r_4__35_, s_r_4__34_, s_r_4__33_, s_r_4__32_, s_r_4__31_, s_r_4__30_, s_r_4__29_, s_r_4__28_, s_r_4__27_, s_r_4__26_, s_r_4__25_, s_r_4__24_, s_r_4__23_, s_r_4__22_, s_r_4__21_, s_r_4__20_, s_r_4__19_, s_r_4__18_, s_r_4__17_, s_r_4__16_, s_r_4__15_, s_r_4__14_, s_r_4__13_, s_r_4__12_, s_r_4__11_, s_r_4__10_, s_r_4__9_, s_r_4__8_, s_r_4__7_, s_r_4__6_, s_r_4__5_, s_r_4__4_, s_r_4__3_, s_r_4__2_, s_r_4__1_, s_r_4__0_ }),
    .c_o(c_r[4]),
    .prod_accum_o({ prod_accum_4__5_, prod_accum_4__4_, prod_accum_4__3_, prod_accum_4__2_, prod_accum_4__1_, prod_accum_4__0_ })
  );


  bsg_mul_array_row_128_5_0
  genblk1_5__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[639:512]),
    .b_i(b_r[639:512]),
    .s_i({ s_r_4__127_, s_r_4__126_, s_r_4__125_, s_r_4__124_, s_r_4__123_, s_r_4__122_, s_r_4__121_, s_r_4__120_, s_r_4__119_, s_r_4__118_, s_r_4__117_, s_r_4__116_, s_r_4__115_, s_r_4__114_, s_r_4__113_, s_r_4__112_, s_r_4__111_, s_r_4__110_, s_r_4__109_, s_r_4__108_, s_r_4__107_, s_r_4__106_, s_r_4__105_, s_r_4__104_, s_r_4__103_, s_r_4__102_, s_r_4__101_, s_r_4__100_, s_r_4__99_, s_r_4__98_, s_r_4__97_, s_r_4__96_, s_r_4__95_, s_r_4__94_, s_r_4__93_, s_r_4__92_, s_r_4__91_, s_r_4__90_, s_r_4__89_, s_r_4__88_, s_r_4__87_, s_r_4__86_, s_r_4__85_, s_r_4__84_, s_r_4__83_, s_r_4__82_, s_r_4__81_, s_r_4__80_, s_r_4__79_, s_r_4__78_, s_r_4__77_, s_r_4__76_, s_r_4__75_, s_r_4__74_, s_r_4__73_, s_r_4__72_, s_r_4__71_, s_r_4__70_, s_r_4__69_, s_r_4__68_, s_r_4__67_, s_r_4__66_, s_r_4__65_, s_r_4__64_, s_r_4__63_, s_r_4__62_, s_r_4__61_, s_r_4__60_, s_r_4__59_, s_r_4__58_, s_r_4__57_, s_r_4__56_, s_r_4__55_, s_r_4__54_, s_r_4__53_, s_r_4__52_, s_r_4__51_, s_r_4__50_, s_r_4__49_, s_r_4__48_, s_r_4__47_, s_r_4__46_, s_r_4__45_, s_r_4__44_, s_r_4__43_, s_r_4__42_, s_r_4__41_, s_r_4__40_, s_r_4__39_, s_r_4__38_, s_r_4__37_, s_r_4__36_, s_r_4__35_, s_r_4__34_, s_r_4__33_, s_r_4__32_, s_r_4__31_, s_r_4__30_, s_r_4__29_, s_r_4__28_, s_r_4__27_, s_r_4__26_, s_r_4__25_, s_r_4__24_, s_r_4__23_, s_r_4__22_, s_r_4__21_, s_r_4__20_, s_r_4__19_, s_r_4__18_, s_r_4__17_, s_r_4__16_, s_r_4__15_, s_r_4__14_, s_r_4__13_, s_r_4__12_, s_r_4__11_, s_r_4__10_, s_r_4__9_, s_r_4__8_, s_r_4__7_, s_r_4__6_, s_r_4__5_, s_r_4__4_, s_r_4__3_, s_r_4__2_, s_r_4__1_, s_r_4__0_ }),
    .c_i(c_r[4]),
    .prod_accum_i({ prod_accum_4__5_, prod_accum_4__4_, prod_accum_4__3_, prod_accum_4__2_, prod_accum_4__1_, prod_accum_4__0_ }),
    .a_o(a_r[767:640]),
    .b_o(b_r[767:640]),
    .s_o({ s_r_5__127_, s_r_5__126_, s_r_5__125_, s_r_5__124_, s_r_5__123_, s_r_5__122_, s_r_5__121_, s_r_5__120_, s_r_5__119_, s_r_5__118_, s_r_5__117_, s_r_5__116_, s_r_5__115_, s_r_5__114_, s_r_5__113_, s_r_5__112_, s_r_5__111_, s_r_5__110_, s_r_5__109_, s_r_5__108_, s_r_5__107_, s_r_5__106_, s_r_5__105_, s_r_5__104_, s_r_5__103_, s_r_5__102_, s_r_5__101_, s_r_5__100_, s_r_5__99_, s_r_5__98_, s_r_5__97_, s_r_5__96_, s_r_5__95_, s_r_5__94_, s_r_5__93_, s_r_5__92_, s_r_5__91_, s_r_5__90_, s_r_5__89_, s_r_5__88_, s_r_5__87_, s_r_5__86_, s_r_5__85_, s_r_5__84_, s_r_5__83_, s_r_5__82_, s_r_5__81_, s_r_5__80_, s_r_5__79_, s_r_5__78_, s_r_5__77_, s_r_5__76_, s_r_5__75_, s_r_5__74_, s_r_5__73_, s_r_5__72_, s_r_5__71_, s_r_5__70_, s_r_5__69_, s_r_5__68_, s_r_5__67_, s_r_5__66_, s_r_5__65_, s_r_5__64_, s_r_5__63_, s_r_5__62_, s_r_5__61_, s_r_5__60_, s_r_5__59_, s_r_5__58_, s_r_5__57_, s_r_5__56_, s_r_5__55_, s_r_5__54_, s_r_5__53_, s_r_5__52_, s_r_5__51_, s_r_5__50_, s_r_5__49_, s_r_5__48_, s_r_5__47_, s_r_5__46_, s_r_5__45_, s_r_5__44_, s_r_5__43_, s_r_5__42_, s_r_5__41_, s_r_5__40_, s_r_5__39_, s_r_5__38_, s_r_5__37_, s_r_5__36_, s_r_5__35_, s_r_5__34_, s_r_5__33_, s_r_5__32_, s_r_5__31_, s_r_5__30_, s_r_5__29_, s_r_5__28_, s_r_5__27_, s_r_5__26_, s_r_5__25_, s_r_5__24_, s_r_5__23_, s_r_5__22_, s_r_5__21_, s_r_5__20_, s_r_5__19_, s_r_5__18_, s_r_5__17_, s_r_5__16_, s_r_5__15_, s_r_5__14_, s_r_5__13_, s_r_5__12_, s_r_5__11_, s_r_5__10_, s_r_5__9_, s_r_5__8_, s_r_5__7_, s_r_5__6_, s_r_5__5_, s_r_5__4_, s_r_5__3_, s_r_5__2_, s_r_5__1_, s_r_5__0_ }),
    .c_o(c_r[5]),
    .prod_accum_o({ prod_accum_5__6_, prod_accum_5__5_, prod_accum_5__4_, prod_accum_5__3_, prod_accum_5__2_, prod_accum_5__1_, prod_accum_5__0_ })
  );


  bsg_mul_array_row_128_6_0
  genblk1_6__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[767:640]),
    .b_i(b_r[767:640]),
    .s_i({ s_r_5__127_, s_r_5__126_, s_r_5__125_, s_r_5__124_, s_r_5__123_, s_r_5__122_, s_r_5__121_, s_r_5__120_, s_r_5__119_, s_r_5__118_, s_r_5__117_, s_r_5__116_, s_r_5__115_, s_r_5__114_, s_r_5__113_, s_r_5__112_, s_r_5__111_, s_r_5__110_, s_r_5__109_, s_r_5__108_, s_r_5__107_, s_r_5__106_, s_r_5__105_, s_r_5__104_, s_r_5__103_, s_r_5__102_, s_r_5__101_, s_r_5__100_, s_r_5__99_, s_r_5__98_, s_r_5__97_, s_r_5__96_, s_r_5__95_, s_r_5__94_, s_r_5__93_, s_r_5__92_, s_r_5__91_, s_r_5__90_, s_r_5__89_, s_r_5__88_, s_r_5__87_, s_r_5__86_, s_r_5__85_, s_r_5__84_, s_r_5__83_, s_r_5__82_, s_r_5__81_, s_r_5__80_, s_r_5__79_, s_r_5__78_, s_r_5__77_, s_r_5__76_, s_r_5__75_, s_r_5__74_, s_r_5__73_, s_r_5__72_, s_r_5__71_, s_r_5__70_, s_r_5__69_, s_r_5__68_, s_r_5__67_, s_r_5__66_, s_r_5__65_, s_r_5__64_, s_r_5__63_, s_r_5__62_, s_r_5__61_, s_r_5__60_, s_r_5__59_, s_r_5__58_, s_r_5__57_, s_r_5__56_, s_r_5__55_, s_r_5__54_, s_r_5__53_, s_r_5__52_, s_r_5__51_, s_r_5__50_, s_r_5__49_, s_r_5__48_, s_r_5__47_, s_r_5__46_, s_r_5__45_, s_r_5__44_, s_r_5__43_, s_r_5__42_, s_r_5__41_, s_r_5__40_, s_r_5__39_, s_r_5__38_, s_r_5__37_, s_r_5__36_, s_r_5__35_, s_r_5__34_, s_r_5__33_, s_r_5__32_, s_r_5__31_, s_r_5__30_, s_r_5__29_, s_r_5__28_, s_r_5__27_, s_r_5__26_, s_r_5__25_, s_r_5__24_, s_r_5__23_, s_r_5__22_, s_r_5__21_, s_r_5__20_, s_r_5__19_, s_r_5__18_, s_r_5__17_, s_r_5__16_, s_r_5__15_, s_r_5__14_, s_r_5__13_, s_r_5__12_, s_r_5__11_, s_r_5__10_, s_r_5__9_, s_r_5__8_, s_r_5__7_, s_r_5__6_, s_r_5__5_, s_r_5__4_, s_r_5__3_, s_r_5__2_, s_r_5__1_, s_r_5__0_ }),
    .c_i(c_r[5]),
    .prod_accum_i({ prod_accum_5__6_, prod_accum_5__5_, prod_accum_5__4_, prod_accum_5__3_, prod_accum_5__2_, prod_accum_5__1_, prod_accum_5__0_ }),
    .a_o(a_r[895:768]),
    .b_o(b_r[895:768]),
    .s_o({ s_r_6__127_, s_r_6__126_, s_r_6__125_, s_r_6__124_, s_r_6__123_, s_r_6__122_, s_r_6__121_, s_r_6__120_, s_r_6__119_, s_r_6__118_, s_r_6__117_, s_r_6__116_, s_r_6__115_, s_r_6__114_, s_r_6__113_, s_r_6__112_, s_r_6__111_, s_r_6__110_, s_r_6__109_, s_r_6__108_, s_r_6__107_, s_r_6__106_, s_r_6__105_, s_r_6__104_, s_r_6__103_, s_r_6__102_, s_r_6__101_, s_r_6__100_, s_r_6__99_, s_r_6__98_, s_r_6__97_, s_r_6__96_, s_r_6__95_, s_r_6__94_, s_r_6__93_, s_r_6__92_, s_r_6__91_, s_r_6__90_, s_r_6__89_, s_r_6__88_, s_r_6__87_, s_r_6__86_, s_r_6__85_, s_r_6__84_, s_r_6__83_, s_r_6__82_, s_r_6__81_, s_r_6__80_, s_r_6__79_, s_r_6__78_, s_r_6__77_, s_r_6__76_, s_r_6__75_, s_r_6__74_, s_r_6__73_, s_r_6__72_, s_r_6__71_, s_r_6__70_, s_r_6__69_, s_r_6__68_, s_r_6__67_, s_r_6__66_, s_r_6__65_, s_r_6__64_, s_r_6__63_, s_r_6__62_, s_r_6__61_, s_r_6__60_, s_r_6__59_, s_r_6__58_, s_r_6__57_, s_r_6__56_, s_r_6__55_, s_r_6__54_, s_r_6__53_, s_r_6__52_, s_r_6__51_, s_r_6__50_, s_r_6__49_, s_r_6__48_, s_r_6__47_, s_r_6__46_, s_r_6__45_, s_r_6__44_, s_r_6__43_, s_r_6__42_, s_r_6__41_, s_r_6__40_, s_r_6__39_, s_r_6__38_, s_r_6__37_, s_r_6__36_, s_r_6__35_, s_r_6__34_, s_r_6__33_, s_r_6__32_, s_r_6__31_, s_r_6__30_, s_r_6__29_, s_r_6__28_, s_r_6__27_, s_r_6__26_, s_r_6__25_, s_r_6__24_, s_r_6__23_, s_r_6__22_, s_r_6__21_, s_r_6__20_, s_r_6__19_, s_r_6__18_, s_r_6__17_, s_r_6__16_, s_r_6__15_, s_r_6__14_, s_r_6__13_, s_r_6__12_, s_r_6__11_, s_r_6__10_, s_r_6__9_, s_r_6__8_, s_r_6__7_, s_r_6__6_, s_r_6__5_, s_r_6__4_, s_r_6__3_, s_r_6__2_, s_r_6__1_, s_r_6__0_ }),
    .c_o(c_r[6]),
    .prod_accum_o({ prod_accum_6__7_, prod_accum_6__6_, prod_accum_6__5_, prod_accum_6__4_, prod_accum_6__3_, prod_accum_6__2_, prod_accum_6__1_, prod_accum_6__0_ })
  );


  bsg_mul_array_row_128_7_0
  genblk1_7__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[895:768]),
    .b_i(b_r[895:768]),
    .s_i({ s_r_6__127_, s_r_6__126_, s_r_6__125_, s_r_6__124_, s_r_6__123_, s_r_6__122_, s_r_6__121_, s_r_6__120_, s_r_6__119_, s_r_6__118_, s_r_6__117_, s_r_6__116_, s_r_6__115_, s_r_6__114_, s_r_6__113_, s_r_6__112_, s_r_6__111_, s_r_6__110_, s_r_6__109_, s_r_6__108_, s_r_6__107_, s_r_6__106_, s_r_6__105_, s_r_6__104_, s_r_6__103_, s_r_6__102_, s_r_6__101_, s_r_6__100_, s_r_6__99_, s_r_6__98_, s_r_6__97_, s_r_6__96_, s_r_6__95_, s_r_6__94_, s_r_6__93_, s_r_6__92_, s_r_6__91_, s_r_6__90_, s_r_6__89_, s_r_6__88_, s_r_6__87_, s_r_6__86_, s_r_6__85_, s_r_6__84_, s_r_6__83_, s_r_6__82_, s_r_6__81_, s_r_6__80_, s_r_6__79_, s_r_6__78_, s_r_6__77_, s_r_6__76_, s_r_6__75_, s_r_6__74_, s_r_6__73_, s_r_6__72_, s_r_6__71_, s_r_6__70_, s_r_6__69_, s_r_6__68_, s_r_6__67_, s_r_6__66_, s_r_6__65_, s_r_6__64_, s_r_6__63_, s_r_6__62_, s_r_6__61_, s_r_6__60_, s_r_6__59_, s_r_6__58_, s_r_6__57_, s_r_6__56_, s_r_6__55_, s_r_6__54_, s_r_6__53_, s_r_6__52_, s_r_6__51_, s_r_6__50_, s_r_6__49_, s_r_6__48_, s_r_6__47_, s_r_6__46_, s_r_6__45_, s_r_6__44_, s_r_6__43_, s_r_6__42_, s_r_6__41_, s_r_6__40_, s_r_6__39_, s_r_6__38_, s_r_6__37_, s_r_6__36_, s_r_6__35_, s_r_6__34_, s_r_6__33_, s_r_6__32_, s_r_6__31_, s_r_6__30_, s_r_6__29_, s_r_6__28_, s_r_6__27_, s_r_6__26_, s_r_6__25_, s_r_6__24_, s_r_6__23_, s_r_6__22_, s_r_6__21_, s_r_6__20_, s_r_6__19_, s_r_6__18_, s_r_6__17_, s_r_6__16_, s_r_6__15_, s_r_6__14_, s_r_6__13_, s_r_6__12_, s_r_6__11_, s_r_6__10_, s_r_6__9_, s_r_6__8_, s_r_6__7_, s_r_6__6_, s_r_6__5_, s_r_6__4_, s_r_6__3_, s_r_6__2_, s_r_6__1_, s_r_6__0_ }),
    .c_i(c_r[6]),
    .prod_accum_i({ prod_accum_6__7_, prod_accum_6__6_, prod_accum_6__5_, prod_accum_6__4_, prod_accum_6__3_, prod_accum_6__2_, prod_accum_6__1_, prod_accum_6__0_ }),
    .a_o(a_r[1023:896]),
    .b_o(b_r[1023:896]),
    .s_o({ s_r_7__127_, s_r_7__126_, s_r_7__125_, s_r_7__124_, s_r_7__123_, s_r_7__122_, s_r_7__121_, s_r_7__120_, s_r_7__119_, s_r_7__118_, s_r_7__117_, s_r_7__116_, s_r_7__115_, s_r_7__114_, s_r_7__113_, s_r_7__112_, s_r_7__111_, s_r_7__110_, s_r_7__109_, s_r_7__108_, s_r_7__107_, s_r_7__106_, s_r_7__105_, s_r_7__104_, s_r_7__103_, s_r_7__102_, s_r_7__101_, s_r_7__100_, s_r_7__99_, s_r_7__98_, s_r_7__97_, s_r_7__96_, s_r_7__95_, s_r_7__94_, s_r_7__93_, s_r_7__92_, s_r_7__91_, s_r_7__90_, s_r_7__89_, s_r_7__88_, s_r_7__87_, s_r_7__86_, s_r_7__85_, s_r_7__84_, s_r_7__83_, s_r_7__82_, s_r_7__81_, s_r_7__80_, s_r_7__79_, s_r_7__78_, s_r_7__77_, s_r_7__76_, s_r_7__75_, s_r_7__74_, s_r_7__73_, s_r_7__72_, s_r_7__71_, s_r_7__70_, s_r_7__69_, s_r_7__68_, s_r_7__67_, s_r_7__66_, s_r_7__65_, s_r_7__64_, s_r_7__63_, s_r_7__62_, s_r_7__61_, s_r_7__60_, s_r_7__59_, s_r_7__58_, s_r_7__57_, s_r_7__56_, s_r_7__55_, s_r_7__54_, s_r_7__53_, s_r_7__52_, s_r_7__51_, s_r_7__50_, s_r_7__49_, s_r_7__48_, s_r_7__47_, s_r_7__46_, s_r_7__45_, s_r_7__44_, s_r_7__43_, s_r_7__42_, s_r_7__41_, s_r_7__40_, s_r_7__39_, s_r_7__38_, s_r_7__37_, s_r_7__36_, s_r_7__35_, s_r_7__34_, s_r_7__33_, s_r_7__32_, s_r_7__31_, s_r_7__30_, s_r_7__29_, s_r_7__28_, s_r_7__27_, s_r_7__26_, s_r_7__25_, s_r_7__24_, s_r_7__23_, s_r_7__22_, s_r_7__21_, s_r_7__20_, s_r_7__19_, s_r_7__18_, s_r_7__17_, s_r_7__16_, s_r_7__15_, s_r_7__14_, s_r_7__13_, s_r_7__12_, s_r_7__11_, s_r_7__10_, s_r_7__9_, s_r_7__8_, s_r_7__7_, s_r_7__6_, s_r_7__5_, s_r_7__4_, s_r_7__3_, s_r_7__2_, s_r_7__1_, s_r_7__0_ }),
    .c_o(c_r[7]),
    .prod_accum_o({ prod_accum_7__8_, prod_accum_7__7_, prod_accum_7__6_, prod_accum_7__5_, prod_accum_7__4_, prod_accum_7__3_, prod_accum_7__2_, prod_accum_7__1_, prod_accum_7__0_ })
  );


  bsg_mul_array_row_128_8_0
  genblk1_8__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[1023:896]),
    .b_i(b_r[1023:896]),
    .s_i({ s_r_7__127_, s_r_7__126_, s_r_7__125_, s_r_7__124_, s_r_7__123_, s_r_7__122_, s_r_7__121_, s_r_7__120_, s_r_7__119_, s_r_7__118_, s_r_7__117_, s_r_7__116_, s_r_7__115_, s_r_7__114_, s_r_7__113_, s_r_7__112_, s_r_7__111_, s_r_7__110_, s_r_7__109_, s_r_7__108_, s_r_7__107_, s_r_7__106_, s_r_7__105_, s_r_7__104_, s_r_7__103_, s_r_7__102_, s_r_7__101_, s_r_7__100_, s_r_7__99_, s_r_7__98_, s_r_7__97_, s_r_7__96_, s_r_7__95_, s_r_7__94_, s_r_7__93_, s_r_7__92_, s_r_7__91_, s_r_7__90_, s_r_7__89_, s_r_7__88_, s_r_7__87_, s_r_7__86_, s_r_7__85_, s_r_7__84_, s_r_7__83_, s_r_7__82_, s_r_7__81_, s_r_7__80_, s_r_7__79_, s_r_7__78_, s_r_7__77_, s_r_7__76_, s_r_7__75_, s_r_7__74_, s_r_7__73_, s_r_7__72_, s_r_7__71_, s_r_7__70_, s_r_7__69_, s_r_7__68_, s_r_7__67_, s_r_7__66_, s_r_7__65_, s_r_7__64_, s_r_7__63_, s_r_7__62_, s_r_7__61_, s_r_7__60_, s_r_7__59_, s_r_7__58_, s_r_7__57_, s_r_7__56_, s_r_7__55_, s_r_7__54_, s_r_7__53_, s_r_7__52_, s_r_7__51_, s_r_7__50_, s_r_7__49_, s_r_7__48_, s_r_7__47_, s_r_7__46_, s_r_7__45_, s_r_7__44_, s_r_7__43_, s_r_7__42_, s_r_7__41_, s_r_7__40_, s_r_7__39_, s_r_7__38_, s_r_7__37_, s_r_7__36_, s_r_7__35_, s_r_7__34_, s_r_7__33_, s_r_7__32_, s_r_7__31_, s_r_7__30_, s_r_7__29_, s_r_7__28_, s_r_7__27_, s_r_7__26_, s_r_7__25_, s_r_7__24_, s_r_7__23_, s_r_7__22_, s_r_7__21_, s_r_7__20_, s_r_7__19_, s_r_7__18_, s_r_7__17_, s_r_7__16_, s_r_7__15_, s_r_7__14_, s_r_7__13_, s_r_7__12_, s_r_7__11_, s_r_7__10_, s_r_7__9_, s_r_7__8_, s_r_7__7_, s_r_7__6_, s_r_7__5_, s_r_7__4_, s_r_7__3_, s_r_7__2_, s_r_7__1_, s_r_7__0_ }),
    .c_i(c_r[7]),
    .prod_accum_i({ prod_accum_7__8_, prod_accum_7__7_, prod_accum_7__6_, prod_accum_7__5_, prod_accum_7__4_, prod_accum_7__3_, prod_accum_7__2_, prod_accum_7__1_, prod_accum_7__0_ }),
    .a_o(a_r[1151:1024]),
    .b_o(b_r[1151:1024]),
    .s_o({ s_r_8__127_, s_r_8__126_, s_r_8__125_, s_r_8__124_, s_r_8__123_, s_r_8__122_, s_r_8__121_, s_r_8__120_, s_r_8__119_, s_r_8__118_, s_r_8__117_, s_r_8__116_, s_r_8__115_, s_r_8__114_, s_r_8__113_, s_r_8__112_, s_r_8__111_, s_r_8__110_, s_r_8__109_, s_r_8__108_, s_r_8__107_, s_r_8__106_, s_r_8__105_, s_r_8__104_, s_r_8__103_, s_r_8__102_, s_r_8__101_, s_r_8__100_, s_r_8__99_, s_r_8__98_, s_r_8__97_, s_r_8__96_, s_r_8__95_, s_r_8__94_, s_r_8__93_, s_r_8__92_, s_r_8__91_, s_r_8__90_, s_r_8__89_, s_r_8__88_, s_r_8__87_, s_r_8__86_, s_r_8__85_, s_r_8__84_, s_r_8__83_, s_r_8__82_, s_r_8__81_, s_r_8__80_, s_r_8__79_, s_r_8__78_, s_r_8__77_, s_r_8__76_, s_r_8__75_, s_r_8__74_, s_r_8__73_, s_r_8__72_, s_r_8__71_, s_r_8__70_, s_r_8__69_, s_r_8__68_, s_r_8__67_, s_r_8__66_, s_r_8__65_, s_r_8__64_, s_r_8__63_, s_r_8__62_, s_r_8__61_, s_r_8__60_, s_r_8__59_, s_r_8__58_, s_r_8__57_, s_r_8__56_, s_r_8__55_, s_r_8__54_, s_r_8__53_, s_r_8__52_, s_r_8__51_, s_r_8__50_, s_r_8__49_, s_r_8__48_, s_r_8__47_, s_r_8__46_, s_r_8__45_, s_r_8__44_, s_r_8__43_, s_r_8__42_, s_r_8__41_, s_r_8__40_, s_r_8__39_, s_r_8__38_, s_r_8__37_, s_r_8__36_, s_r_8__35_, s_r_8__34_, s_r_8__33_, s_r_8__32_, s_r_8__31_, s_r_8__30_, s_r_8__29_, s_r_8__28_, s_r_8__27_, s_r_8__26_, s_r_8__25_, s_r_8__24_, s_r_8__23_, s_r_8__22_, s_r_8__21_, s_r_8__20_, s_r_8__19_, s_r_8__18_, s_r_8__17_, s_r_8__16_, s_r_8__15_, s_r_8__14_, s_r_8__13_, s_r_8__12_, s_r_8__11_, s_r_8__10_, s_r_8__9_, s_r_8__8_, s_r_8__7_, s_r_8__6_, s_r_8__5_, s_r_8__4_, s_r_8__3_, s_r_8__2_, s_r_8__1_, s_r_8__0_ }),
    .c_o(c_r[8]),
    .prod_accum_o({ prod_accum_8__9_, prod_accum_8__8_, prod_accum_8__7_, prod_accum_8__6_, prod_accum_8__5_, prod_accum_8__4_, prod_accum_8__3_, prod_accum_8__2_, prod_accum_8__1_, prod_accum_8__0_ })
  );


  bsg_mul_array_row_128_9_0
  genblk1_9__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[1151:1024]),
    .b_i(b_r[1151:1024]),
    .s_i({ s_r_8__127_, s_r_8__126_, s_r_8__125_, s_r_8__124_, s_r_8__123_, s_r_8__122_, s_r_8__121_, s_r_8__120_, s_r_8__119_, s_r_8__118_, s_r_8__117_, s_r_8__116_, s_r_8__115_, s_r_8__114_, s_r_8__113_, s_r_8__112_, s_r_8__111_, s_r_8__110_, s_r_8__109_, s_r_8__108_, s_r_8__107_, s_r_8__106_, s_r_8__105_, s_r_8__104_, s_r_8__103_, s_r_8__102_, s_r_8__101_, s_r_8__100_, s_r_8__99_, s_r_8__98_, s_r_8__97_, s_r_8__96_, s_r_8__95_, s_r_8__94_, s_r_8__93_, s_r_8__92_, s_r_8__91_, s_r_8__90_, s_r_8__89_, s_r_8__88_, s_r_8__87_, s_r_8__86_, s_r_8__85_, s_r_8__84_, s_r_8__83_, s_r_8__82_, s_r_8__81_, s_r_8__80_, s_r_8__79_, s_r_8__78_, s_r_8__77_, s_r_8__76_, s_r_8__75_, s_r_8__74_, s_r_8__73_, s_r_8__72_, s_r_8__71_, s_r_8__70_, s_r_8__69_, s_r_8__68_, s_r_8__67_, s_r_8__66_, s_r_8__65_, s_r_8__64_, s_r_8__63_, s_r_8__62_, s_r_8__61_, s_r_8__60_, s_r_8__59_, s_r_8__58_, s_r_8__57_, s_r_8__56_, s_r_8__55_, s_r_8__54_, s_r_8__53_, s_r_8__52_, s_r_8__51_, s_r_8__50_, s_r_8__49_, s_r_8__48_, s_r_8__47_, s_r_8__46_, s_r_8__45_, s_r_8__44_, s_r_8__43_, s_r_8__42_, s_r_8__41_, s_r_8__40_, s_r_8__39_, s_r_8__38_, s_r_8__37_, s_r_8__36_, s_r_8__35_, s_r_8__34_, s_r_8__33_, s_r_8__32_, s_r_8__31_, s_r_8__30_, s_r_8__29_, s_r_8__28_, s_r_8__27_, s_r_8__26_, s_r_8__25_, s_r_8__24_, s_r_8__23_, s_r_8__22_, s_r_8__21_, s_r_8__20_, s_r_8__19_, s_r_8__18_, s_r_8__17_, s_r_8__16_, s_r_8__15_, s_r_8__14_, s_r_8__13_, s_r_8__12_, s_r_8__11_, s_r_8__10_, s_r_8__9_, s_r_8__8_, s_r_8__7_, s_r_8__6_, s_r_8__5_, s_r_8__4_, s_r_8__3_, s_r_8__2_, s_r_8__1_, s_r_8__0_ }),
    .c_i(c_r[8]),
    .prod_accum_i({ prod_accum_8__9_, prod_accum_8__8_, prod_accum_8__7_, prod_accum_8__6_, prod_accum_8__5_, prod_accum_8__4_, prod_accum_8__3_, prod_accum_8__2_, prod_accum_8__1_, prod_accum_8__0_ }),
    .a_o(a_r[1279:1152]),
    .b_o(b_r[1279:1152]),
    .s_o({ s_r_9__127_, s_r_9__126_, s_r_9__125_, s_r_9__124_, s_r_9__123_, s_r_9__122_, s_r_9__121_, s_r_9__120_, s_r_9__119_, s_r_9__118_, s_r_9__117_, s_r_9__116_, s_r_9__115_, s_r_9__114_, s_r_9__113_, s_r_9__112_, s_r_9__111_, s_r_9__110_, s_r_9__109_, s_r_9__108_, s_r_9__107_, s_r_9__106_, s_r_9__105_, s_r_9__104_, s_r_9__103_, s_r_9__102_, s_r_9__101_, s_r_9__100_, s_r_9__99_, s_r_9__98_, s_r_9__97_, s_r_9__96_, s_r_9__95_, s_r_9__94_, s_r_9__93_, s_r_9__92_, s_r_9__91_, s_r_9__90_, s_r_9__89_, s_r_9__88_, s_r_9__87_, s_r_9__86_, s_r_9__85_, s_r_9__84_, s_r_9__83_, s_r_9__82_, s_r_9__81_, s_r_9__80_, s_r_9__79_, s_r_9__78_, s_r_9__77_, s_r_9__76_, s_r_9__75_, s_r_9__74_, s_r_9__73_, s_r_9__72_, s_r_9__71_, s_r_9__70_, s_r_9__69_, s_r_9__68_, s_r_9__67_, s_r_9__66_, s_r_9__65_, s_r_9__64_, s_r_9__63_, s_r_9__62_, s_r_9__61_, s_r_9__60_, s_r_9__59_, s_r_9__58_, s_r_9__57_, s_r_9__56_, s_r_9__55_, s_r_9__54_, s_r_9__53_, s_r_9__52_, s_r_9__51_, s_r_9__50_, s_r_9__49_, s_r_9__48_, s_r_9__47_, s_r_9__46_, s_r_9__45_, s_r_9__44_, s_r_9__43_, s_r_9__42_, s_r_9__41_, s_r_9__40_, s_r_9__39_, s_r_9__38_, s_r_9__37_, s_r_9__36_, s_r_9__35_, s_r_9__34_, s_r_9__33_, s_r_9__32_, s_r_9__31_, s_r_9__30_, s_r_9__29_, s_r_9__28_, s_r_9__27_, s_r_9__26_, s_r_9__25_, s_r_9__24_, s_r_9__23_, s_r_9__22_, s_r_9__21_, s_r_9__20_, s_r_9__19_, s_r_9__18_, s_r_9__17_, s_r_9__16_, s_r_9__15_, s_r_9__14_, s_r_9__13_, s_r_9__12_, s_r_9__11_, s_r_9__10_, s_r_9__9_, s_r_9__8_, s_r_9__7_, s_r_9__6_, s_r_9__5_, s_r_9__4_, s_r_9__3_, s_r_9__2_, s_r_9__1_, s_r_9__0_ }),
    .c_o(c_r[9]),
    .prod_accum_o({ prod_accum_9__10_, prod_accum_9__9_, prod_accum_9__8_, prod_accum_9__7_, prod_accum_9__6_, prod_accum_9__5_, prod_accum_9__4_, prod_accum_9__3_, prod_accum_9__2_, prod_accum_9__1_, prod_accum_9__0_ })
  );


  bsg_mul_array_row_128_10_0
  genblk1_10__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[1279:1152]),
    .b_i(b_r[1279:1152]),
    .s_i({ s_r_9__127_, s_r_9__126_, s_r_9__125_, s_r_9__124_, s_r_9__123_, s_r_9__122_, s_r_9__121_, s_r_9__120_, s_r_9__119_, s_r_9__118_, s_r_9__117_, s_r_9__116_, s_r_9__115_, s_r_9__114_, s_r_9__113_, s_r_9__112_, s_r_9__111_, s_r_9__110_, s_r_9__109_, s_r_9__108_, s_r_9__107_, s_r_9__106_, s_r_9__105_, s_r_9__104_, s_r_9__103_, s_r_9__102_, s_r_9__101_, s_r_9__100_, s_r_9__99_, s_r_9__98_, s_r_9__97_, s_r_9__96_, s_r_9__95_, s_r_9__94_, s_r_9__93_, s_r_9__92_, s_r_9__91_, s_r_9__90_, s_r_9__89_, s_r_9__88_, s_r_9__87_, s_r_9__86_, s_r_9__85_, s_r_9__84_, s_r_9__83_, s_r_9__82_, s_r_9__81_, s_r_9__80_, s_r_9__79_, s_r_9__78_, s_r_9__77_, s_r_9__76_, s_r_9__75_, s_r_9__74_, s_r_9__73_, s_r_9__72_, s_r_9__71_, s_r_9__70_, s_r_9__69_, s_r_9__68_, s_r_9__67_, s_r_9__66_, s_r_9__65_, s_r_9__64_, s_r_9__63_, s_r_9__62_, s_r_9__61_, s_r_9__60_, s_r_9__59_, s_r_9__58_, s_r_9__57_, s_r_9__56_, s_r_9__55_, s_r_9__54_, s_r_9__53_, s_r_9__52_, s_r_9__51_, s_r_9__50_, s_r_9__49_, s_r_9__48_, s_r_9__47_, s_r_9__46_, s_r_9__45_, s_r_9__44_, s_r_9__43_, s_r_9__42_, s_r_9__41_, s_r_9__40_, s_r_9__39_, s_r_9__38_, s_r_9__37_, s_r_9__36_, s_r_9__35_, s_r_9__34_, s_r_9__33_, s_r_9__32_, s_r_9__31_, s_r_9__30_, s_r_9__29_, s_r_9__28_, s_r_9__27_, s_r_9__26_, s_r_9__25_, s_r_9__24_, s_r_9__23_, s_r_9__22_, s_r_9__21_, s_r_9__20_, s_r_9__19_, s_r_9__18_, s_r_9__17_, s_r_9__16_, s_r_9__15_, s_r_9__14_, s_r_9__13_, s_r_9__12_, s_r_9__11_, s_r_9__10_, s_r_9__9_, s_r_9__8_, s_r_9__7_, s_r_9__6_, s_r_9__5_, s_r_9__4_, s_r_9__3_, s_r_9__2_, s_r_9__1_, s_r_9__0_ }),
    .c_i(c_r[9]),
    .prod_accum_i({ prod_accum_9__10_, prod_accum_9__9_, prod_accum_9__8_, prod_accum_9__7_, prod_accum_9__6_, prod_accum_9__5_, prod_accum_9__4_, prod_accum_9__3_, prod_accum_9__2_, prod_accum_9__1_, prod_accum_9__0_ }),
    .a_o(a_r[1407:1280]),
    .b_o(b_r[1407:1280]),
    .s_o({ s_r_10__127_, s_r_10__126_, s_r_10__125_, s_r_10__124_, s_r_10__123_, s_r_10__122_, s_r_10__121_, s_r_10__120_, s_r_10__119_, s_r_10__118_, s_r_10__117_, s_r_10__116_, s_r_10__115_, s_r_10__114_, s_r_10__113_, s_r_10__112_, s_r_10__111_, s_r_10__110_, s_r_10__109_, s_r_10__108_, s_r_10__107_, s_r_10__106_, s_r_10__105_, s_r_10__104_, s_r_10__103_, s_r_10__102_, s_r_10__101_, s_r_10__100_, s_r_10__99_, s_r_10__98_, s_r_10__97_, s_r_10__96_, s_r_10__95_, s_r_10__94_, s_r_10__93_, s_r_10__92_, s_r_10__91_, s_r_10__90_, s_r_10__89_, s_r_10__88_, s_r_10__87_, s_r_10__86_, s_r_10__85_, s_r_10__84_, s_r_10__83_, s_r_10__82_, s_r_10__81_, s_r_10__80_, s_r_10__79_, s_r_10__78_, s_r_10__77_, s_r_10__76_, s_r_10__75_, s_r_10__74_, s_r_10__73_, s_r_10__72_, s_r_10__71_, s_r_10__70_, s_r_10__69_, s_r_10__68_, s_r_10__67_, s_r_10__66_, s_r_10__65_, s_r_10__64_, s_r_10__63_, s_r_10__62_, s_r_10__61_, s_r_10__60_, s_r_10__59_, s_r_10__58_, s_r_10__57_, s_r_10__56_, s_r_10__55_, s_r_10__54_, s_r_10__53_, s_r_10__52_, s_r_10__51_, s_r_10__50_, s_r_10__49_, s_r_10__48_, s_r_10__47_, s_r_10__46_, s_r_10__45_, s_r_10__44_, s_r_10__43_, s_r_10__42_, s_r_10__41_, s_r_10__40_, s_r_10__39_, s_r_10__38_, s_r_10__37_, s_r_10__36_, s_r_10__35_, s_r_10__34_, s_r_10__33_, s_r_10__32_, s_r_10__31_, s_r_10__30_, s_r_10__29_, s_r_10__28_, s_r_10__27_, s_r_10__26_, s_r_10__25_, s_r_10__24_, s_r_10__23_, s_r_10__22_, s_r_10__21_, s_r_10__20_, s_r_10__19_, s_r_10__18_, s_r_10__17_, s_r_10__16_, s_r_10__15_, s_r_10__14_, s_r_10__13_, s_r_10__12_, s_r_10__11_, s_r_10__10_, s_r_10__9_, s_r_10__8_, s_r_10__7_, s_r_10__6_, s_r_10__5_, s_r_10__4_, s_r_10__3_, s_r_10__2_, s_r_10__1_, s_r_10__0_ }),
    .c_o(c_r[10]),
    .prod_accum_o({ prod_accum_10__11_, prod_accum_10__10_, prod_accum_10__9_, prod_accum_10__8_, prod_accum_10__7_, prod_accum_10__6_, prod_accum_10__5_, prod_accum_10__4_, prod_accum_10__3_, prod_accum_10__2_, prod_accum_10__1_, prod_accum_10__0_ })
  );


  bsg_mul_array_row_128_11_0
  genblk1_11__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[1407:1280]),
    .b_i(b_r[1407:1280]),
    .s_i({ s_r_10__127_, s_r_10__126_, s_r_10__125_, s_r_10__124_, s_r_10__123_, s_r_10__122_, s_r_10__121_, s_r_10__120_, s_r_10__119_, s_r_10__118_, s_r_10__117_, s_r_10__116_, s_r_10__115_, s_r_10__114_, s_r_10__113_, s_r_10__112_, s_r_10__111_, s_r_10__110_, s_r_10__109_, s_r_10__108_, s_r_10__107_, s_r_10__106_, s_r_10__105_, s_r_10__104_, s_r_10__103_, s_r_10__102_, s_r_10__101_, s_r_10__100_, s_r_10__99_, s_r_10__98_, s_r_10__97_, s_r_10__96_, s_r_10__95_, s_r_10__94_, s_r_10__93_, s_r_10__92_, s_r_10__91_, s_r_10__90_, s_r_10__89_, s_r_10__88_, s_r_10__87_, s_r_10__86_, s_r_10__85_, s_r_10__84_, s_r_10__83_, s_r_10__82_, s_r_10__81_, s_r_10__80_, s_r_10__79_, s_r_10__78_, s_r_10__77_, s_r_10__76_, s_r_10__75_, s_r_10__74_, s_r_10__73_, s_r_10__72_, s_r_10__71_, s_r_10__70_, s_r_10__69_, s_r_10__68_, s_r_10__67_, s_r_10__66_, s_r_10__65_, s_r_10__64_, s_r_10__63_, s_r_10__62_, s_r_10__61_, s_r_10__60_, s_r_10__59_, s_r_10__58_, s_r_10__57_, s_r_10__56_, s_r_10__55_, s_r_10__54_, s_r_10__53_, s_r_10__52_, s_r_10__51_, s_r_10__50_, s_r_10__49_, s_r_10__48_, s_r_10__47_, s_r_10__46_, s_r_10__45_, s_r_10__44_, s_r_10__43_, s_r_10__42_, s_r_10__41_, s_r_10__40_, s_r_10__39_, s_r_10__38_, s_r_10__37_, s_r_10__36_, s_r_10__35_, s_r_10__34_, s_r_10__33_, s_r_10__32_, s_r_10__31_, s_r_10__30_, s_r_10__29_, s_r_10__28_, s_r_10__27_, s_r_10__26_, s_r_10__25_, s_r_10__24_, s_r_10__23_, s_r_10__22_, s_r_10__21_, s_r_10__20_, s_r_10__19_, s_r_10__18_, s_r_10__17_, s_r_10__16_, s_r_10__15_, s_r_10__14_, s_r_10__13_, s_r_10__12_, s_r_10__11_, s_r_10__10_, s_r_10__9_, s_r_10__8_, s_r_10__7_, s_r_10__6_, s_r_10__5_, s_r_10__4_, s_r_10__3_, s_r_10__2_, s_r_10__1_, s_r_10__0_ }),
    .c_i(c_r[10]),
    .prod_accum_i({ prod_accum_10__11_, prod_accum_10__10_, prod_accum_10__9_, prod_accum_10__8_, prod_accum_10__7_, prod_accum_10__6_, prod_accum_10__5_, prod_accum_10__4_, prod_accum_10__3_, prod_accum_10__2_, prod_accum_10__1_, prod_accum_10__0_ }),
    .a_o(a_r[1535:1408]),
    .b_o(b_r[1535:1408]),
    .s_o({ s_r_11__127_, s_r_11__126_, s_r_11__125_, s_r_11__124_, s_r_11__123_, s_r_11__122_, s_r_11__121_, s_r_11__120_, s_r_11__119_, s_r_11__118_, s_r_11__117_, s_r_11__116_, s_r_11__115_, s_r_11__114_, s_r_11__113_, s_r_11__112_, s_r_11__111_, s_r_11__110_, s_r_11__109_, s_r_11__108_, s_r_11__107_, s_r_11__106_, s_r_11__105_, s_r_11__104_, s_r_11__103_, s_r_11__102_, s_r_11__101_, s_r_11__100_, s_r_11__99_, s_r_11__98_, s_r_11__97_, s_r_11__96_, s_r_11__95_, s_r_11__94_, s_r_11__93_, s_r_11__92_, s_r_11__91_, s_r_11__90_, s_r_11__89_, s_r_11__88_, s_r_11__87_, s_r_11__86_, s_r_11__85_, s_r_11__84_, s_r_11__83_, s_r_11__82_, s_r_11__81_, s_r_11__80_, s_r_11__79_, s_r_11__78_, s_r_11__77_, s_r_11__76_, s_r_11__75_, s_r_11__74_, s_r_11__73_, s_r_11__72_, s_r_11__71_, s_r_11__70_, s_r_11__69_, s_r_11__68_, s_r_11__67_, s_r_11__66_, s_r_11__65_, s_r_11__64_, s_r_11__63_, s_r_11__62_, s_r_11__61_, s_r_11__60_, s_r_11__59_, s_r_11__58_, s_r_11__57_, s_r_11__56_, s_r_11__55_, s_r_11__54_, s_r_11__53_, s_r_11__52_, s_r_11__51_, s_r_11__50_, s_r_11__49_, s_r_11__48_, s_r_11__47_, s_r_11__46_, s_r_11__45_, s_r_11__44_, s_r_11__43_, s_r_11__42_, s_r_11__41_, s_r_11__40_, s_r_11__39_, s_r_11__38_, s_r_11__37_, s_r_11__36_, s_r_11__35_, s_r_11__34_, s_r_11__33_, s_r_11__32_, s_r_11__31_, s_r_11__30_, s_r_11__29_, s_r_11__28_, s_r_11__27_, s_r_11__26_, s_r_11__25_, s_r_11__24_, s_r_11__23_, s_r_11__22_, s_r_11__21_, s_r_11__20_, s_r_11__19_, s_r_11__18_, s_r_11__17_, s_r_11__16_, s_r_11__15_, s_r_11__14_, s_r_11__13_, s_r_11__12_, s_r_11__11_, s_r_11__10_, s_r_11__9_, s_r_11__8_, s_r_11__7_, s_r_11__6_, s_r_11__5_, s_r_11__4_, s_r_11__3_, s_r_11__2_, s_r_11__1_, s_r_11__0_ }),
    .c_o(c_r[11]),
    .prod_accum_o({ prod_accum_11__12_, prod_accum_11__11_, prod_accum_11__10_, prod_accum_11__9_, prod_accum_11__8_, prod_accum_11__7_, prod_accum_11__6_, prod_accum_11__5_, prod_accum_11__4_, prod_accum_11__3_, prod_accum_11__2_, prod_accum_11__1_, prod_accum_11__0_ })
  );


  bsg_mul_array_row_128_12_0
  genblk1_12__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[1535:1408]),
    .b_i(b_r[1535:1408]),
    .s_i({ s_r_11__127_, s_r_11__126_, s_r_11__125_, s_r_11__124_, s_r_11__123_, s_r_11__122_, s_r_11__121_, s_r_11__120_, s_r_11__119_, s_r_11__118_, s_r_11__117_, s_r_11__116_, s_r_11__115_, s_r_11__114_, s_r_11__113_, s_r_11__112_, s_r_11__111_, s_r_11__110_, s_r_11__109_, s_r_11__108_, s_r_11__107_, s_r_11__106_, s_r_11__105_, s_r_11__104_, s_r_11__103_, s_r_11__102_, s_r_11__101_, s_r_11__100_, s_r_11__99_, s_r_11__98_, s_r_11__97_, s_r_11__96_, s_r_11__95_, s_r_11__94_, s_r_11__93_, s_r_11__92_, s_r_11__91_, s_r_11__90_, s_r_11__89_, s_r_11__88_, s_r_11__87_, s_r_11__86_, s_r_11__85_, s_r_11__84_, s_r_11__83_, s_r_11__82_, s_r_11__81_, s_r_11__80_, s_r_11__79_, s_r_11__78_, s_r_11__77_, s_r_11__76_, s_r_11__75_, s_r_11__74_, s_r_11__73_, s_r_11__72_, s_r_11__71_, s_r_11__70_, s_r_11__69_, s_r_11__68_, s_r_11__67_, s_r_11__66_, s_r_11__65_, s_r_11__64_, s_r_11__63_, s_r_11__62_, s_r_11__61_, s_r_11__60_, s_r_11__59_, s_r_11__58_, s_r_11__57_, s_r_11__56_, s_r_11__55_, s_r_11__54_, s_r_11__53_, s_r_11__52_, s_r_11__51_, s_r_11__50_, s_r_11__49_, s_r_11__48_, s_r_11__47_, s_r_11__46_, s_r_11__45_, s_r_11__44_, s_r_11__43_, s_r_11__42_, s_r_11__41_, s_r_11__40_, s_r_11__39_, s_r_11__38_, s_r_11__37_, s_r_11__36_, s_r_11__35_, s_r_11__34_, s_r_11__33_, s_r_11__32_, s_r_11__31_, s_r_11__30_, s_r_11__29_, s_r_11__28_, s_r_11__27_, s_r_11__26_, s_r_11__25_, s_r_11__24_, s_r_11__23_, s_r_11__22_, s_r_11__21_, s_r_11__20_, s_r_11__19_, s_r_11__18_, s_r_11__17_, s_r_11__16_, s_r_11__15_, s_r_11__14_, s_r_11__13_, s_r_11__12_, s_r_11__11_, s_r_11__10_, s_r_11__9_, s_r_11__8_, s_r_11__7_, s_r_11__6_, s_r_11__5_, s_r_11__4_, s_r_11__3_, s_r_11__2_, s_r_11__1_, s_r_11__0_ }),
    .c_i(c_r[11]),
    .prod_accum_i({ prod_accum_11__12_, prod_accum_11__11_, prod_accum_11__10_, prod_accum_11__9_, prod_accum_11__8_, prod_accum_11__7_, prod_accum_11__6_, prod_accum_11__5_, prod_accum_11__4_, prod_accum_11__3_, prod_accum_11__2_, prod_accum_11__1_, prod_accum_11__0_ }),
    .a_o(a_r[1663:1536]),
    .b_o(b_r[1663:1536]),
    .s_o({ s_r_12__127_, s_r_12__126_, s_r_12__125_, s_r_12__124_, s_r_12__123_, s_r_12__122_, s_r_12__121_, s_r_12__120_, s_r_12__119_, s_r_12__118_, s_r_12__117_, s_r_12__116_, s_r_12__115_, s_r_12__114_, s_r_12__113_, s_r_12__112_, s_r_12__111_, s_r_12__110_, s_r_12__109_, s_r_12__108_, s_r_12__107_, s_r_12__106_, s_r_12__105_, s_r_12__104_, s_r_12__103_, s_r_12__102_, s_r_12__101_, s_r_12__100_, s_r_12__99_, s_r_12__98_, s_r_12__97_, s_r_12__96_, s_r_12__95_, s_r_12__94_, s_r_12__93_, s_r_12__92_, s_r_12__91_, s_r_12__90_, s_r_12__89_, s_r_12__88_, s_r_12__87_, s_r_12__86_, s_r_12__85_, s_r_12__84_, s_r_12__83_, s_r_12__82_, s_r_12__81_, s_r_12__80_, s_r_12__79_, s_r_12__78_, s_r_12__77_, s_r_12__76_, s_r_12__75_, s_r_12__74_, s_r_12__73_, s_r_12__72_, s_r_12__71_, s_r_12__70_, s_r_12__69_, s_r_12__68_, s_r_12__67_, s_r_12__66_, s_r_12__65_, s_r_12__64_, s_r_12__63_, s_r_12__62_, s_r_12__61_, s_r_12__60_, s_r_12__59_, s_r_12__58_, s_r_12__57_, s_r_12__56_, s_r_12__55_, s_r_12__54_, s_r_12__53_, s_r_12__52_, s_r_12__51_, s_r_12__50_, s_r_12__49_, s_r_12__48_, s_r_12__47_, s_r_12__46_, s_r_12__45_, s_r_12__44_, s_r_12__43_, s_r_12__42_, s_r_12__41_, s_r_12__40_, s_r_12__39_, s_r_12__38_, s_r_12__37_, s_r_12__36_, s_r_12__35_, s_r_12__34_, s_r_12__33_, s_r_12__32_, s_r_12__31_, s_r_12__30_, s_r_12__29_, s_r_12__28_, s_r_12__27_, s_r_12__26_, s_r_12__25_, s_r_12__24_, s_r_12__23_, s_r_12__22_, s_r_12__21_, s_r_12__20_, s_r_12__19_, s_r_12__18_, s_r_12__17_, s_r_12__16_, s_r_12__15_, s_r_12__14_, s_r_12__13_, s_r_12__12_, s_r_12__11_, s_r_12__10_, s_r_12__9_, s_r_12__8_, s_r_12__7_, s_r_12__6_, s_r_12__5_, s_r_12__4_, s_r_12__3_, s_r_12__2_, s_r_12__1_, s_r_12__0_ }),
    .c_o(c_r[12]),
    .prod_accum_o({ prod_accum_12__13_, prod_accum_12__12_, prod_accum_12__11_, prod_accum_12__10_, prod_accum_12__9_, prod_accum_12__8_, prod_accum_12__7_, prod_accum_12__6_, prod_accum_12__5_, prod_accum_12__4_, prod_accum_12__3_, prod_accum_12__2_, prod_accum_12__1_, prod_accum_12__0_ })
  );


  bsg_mul_array_row_128_13_0
  genblk1_13__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[1663:1536]),
    .b_i(b_r[1663:1536]),
    .s_i({ s_r_12__127_, s_r_12__126_, s_r_12__125_, s_r_12__124_, s_r_12__123_, s_r_12__122_, s_r_12__121_, s_r_12__120_, s_r_12__119_, s_r_12__118_, s_r_12__117_, s_r_12__116_, s_r_12__115_, s_r_12__114_, s_r_12__113_, s_r_12__112_, s_r_12__111_, s_r_12__110_, s_r_12__109_, s_r_12__108_, s_r_12__107_, s_r_12__106_, s_r_12__105_, s_r_12__104_, s_r_12__103_, s_r_12__102_, s_r_12__101_, s_r_12__100_, s_r_12__99_, s_r_12__98_, s_r_12__97_, s_r_12__96_, s_r_12__95_, s_r_12__94_, s_r_12__93_, s_r_12__92_, s_r_12__91_, s_r_12__90_, s_r_12__89_, s_r_12__88_, s_r_12__87_, s_r_12__86_, s_r_12__85_, s_r_12__84_, s_r_12__83_, s_r_12__82_, s_r_12__81_, s_r_12__80_, s_r_12__79_, s_r_12__78_, s_r_12__77_, s_r_12__76_, s_r_12__75_, s_r_12__74_, s_r_12__73_, s_r_12__72_, s_r_12__71_, s_r_12__70_, s_r_12__69_, s_r_12__68_, s_r_12__67_, s_r_12__66_, s_r_12__65_, s_r_12__64_, s_r_12__63_, s_r_12__62_, s_r_12__61_, s_r_12__60_, s_r_12__59_, s_r_12__58_, s_r_12__57_, s_r_12__56_, s_r_12__55_, s_r_12__54_, s_r_12__53_, s_r_12__52_, s_r_12__51_, s_r_12__50_, s_r_12__49_, s_r_12__48_, s_r_12__47_, s_r_12__46_, s_r_12__45_, s_r_12__44_, s_r_12__43_, s_r_12__42_, s_r_12__41_, s_r_12__40_, s_r_12__39_, s_r_12__38_, s_r_12__37_, s_r_12__36_, s_r_12__35_, s_r_12__34_, s_r_12__33_, s_r_12__32_, s_r_12__31_, s_r_12__30_, s_r_12__29_, s_r_12__28_, s_r_12__27_, s_r_12__26_, s_r_12__25_, s_r_12__24_, s_r_12__23_, s_r_12__22_, s_r_12__21_, s_r_12__20_, s_r_12__19_, s_r_12__18_, s_r_12__17_, s_r_12__16_, s_r_12__15_, s_r_12__14_, s_r_12__13_, s_r_12__12_, s_r_12__11_, s_r_12__10_, s_r_12__9_, s_r_12__8_, s_r_12__7_, s_r_12__6_, s_r_12__5_, s_r_12__4_, s_r_12__3_, s_r_12__2_, s_r_12__1_, s_r_12__0_ }),
    .c_i(c_r[12]),
    .prod_accum_i({ prod_accum_12__13_, prod_accum_12__12_, prod_accum_12__11_, prod_accum_12__10_, prod_accum_12__9_, prod_accum_12__8_, prod_accum_12__7_, prod_accum_12__6_, prod_accum_12__5_, prod_accum_12__4_, prod_accum_12__3_, prod_accum_12__2_, prod_accum_12__1_, prod_accum_12__0_ }),
    .a_o(a_r[1791:1664]),
    .b_o(b_r[1791:1664]),
    .s_o({ s_r_13__127_, s_r_13__126_, s_r_13__125_, s_r_13__124_, s_r_13__123_, s_r_13__122_, s_r_13__121_, s_r_13__120_, s_r_13__119_, s_r_13__118_, s_r_13__117_, s_r_13__116_, s_r_13__115_, s_r_13__114_, s_r_13__113_, s_r_13__112_, s_r_13__111_, s_r_13__110_, s_r_13__109_, s_r_13__108_, s_r_13__107_, s_r_13__106_, s_r_13__105_, s_r_13__104_, s_r_13__103_, s_r_13__102_, s_r_13__101_, s_r_13__100_, s_r_13__99_, s_r_13__98_, s_r_13__97_, s_r_13__96_, s_r_13__95_, s_r_13__94_, s_r_13__93_, s_r_13__92_, s_r_13__91_, s_r_13__90_, s_r_13__89_, s_r_13__88_, s_r_13__87_, s_r_13__86_, s_r_13__85_, s_r_13__84_, s_r_13__83_, s_r_13__82_, s_r_13__81_, s_r_13__80_, s_r_13__79_, s_r_13__78_, s_r_13__77_, s_r_13__76_, s_r_13__75_, s_r_13__74_, s_r_13__73_, s_r_13__72_, s_r_13__71_, s_r_13__70_, s_r_13__69_, s_r_13__68_, s_r_13__67_, s_r_13__66_, s_r_13__65_, s_r_13__64_, s_r_13__63_, s_r_13__62_, s_r_13__61_, s_r_13__60_, s_r_13__59_, s_r_13__58_, s_r_13__57_, s_r_13__56_, s_r_13__55_, s_r_13__54_, s_r_13__53_, s_r_13__52_, s_r_13__51_, s_r_13__50_, s_r_13__49_, s_r_13__48_, s_r_13__47_, s_r_13__46_, s_r_13__45_, s_r_13__44_, s_r_13__43_, s_r_13__42_, s_r_13__41_, s_r_13__40_, s_r_13__39_, s_r_13__38_, s_r_13__37_, s_r_13__36_, s_r_13__35_, s_r_13__34_, s_r_13__33_, s_r_13__32_, s_r_13__31_, s_r_13__30_, s_r_13__29_, s_r_13__28_, s_r_13__27_, s_r_13__26_, s_r_13__25_, s_r_13__24_, s_r_13__23_, s_r_13__22_, s_r_13__21_, s_r_13__20_, s_r_13__19_, s_r_13__18_, s_r_13__17_, s_r_13__16_, s_r_13__15_, s_r_13__14_, s_r_13__13_, s_r_13__12_, s_r_13__11_, s_r_13__10_, s_r_13__9_, s_r_13__8_, s_r_13__7_, s_r_13__6_, s_r_13__5_, s_r_13__4_, s_r_13__3_, s_r_13__2_, s_r_13__1_, s_r_13__0_ }),
    .c_o(c_r[13]),
    .prod_accum_o({ prod_accum_13__14_, prod_accum_13__13_, prod_accum_13__12_, prod_accum_13__11_, prod_accum_13__10_, prod_accum_13__9_, prod_accum_13__8_, prod_accum_13__7_, prod_accum_13__6_, prod_accum_13__5_, prod_accum_13__4_, prod_accum_13__3_, prod_accum_13__2_, prod_accum_13__1_, prod_accum_13__0_ })
  );


  bsg_mul_array_row_128_14_0
  genblk1_14__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[1791:1664]),
    .b_i(b_r[1791:1664]),
    .s_i({ s_r_13__127_, s_r_13__126_, s_r_13__125_, s_r_13__124_, s_r_13__123_, s_r_13__122_, s_r_13__121_, s_r_13__120_, s_r_13__119_, s_r_13__118_, s_r_13__117_, s_r_13__116_, s_r_13__115_, s_r_13__114_, s_r_13__113_, s_r_13__112_, s_r_13__111_, s_r_13__110_, s_r_13__109_, s_r_13__108_, s_r_13__107_, s_r_13__106_, s_r_13__105_, s_r_13__104_, s_r_13__103_, s_r_13__102_, s_r_13__101_, s_r_13__100_, s_r_13__99_, s_r_13__98_, s_r_13__97_, s_r_13__96_, s_r_13__95_, s_r_13__94_, s_r_13__93_, s_r_13__92_, s_r_13__91_, s_r_13__90_, s_r_13__89_, s_r_13__88_, s_r_13__87_, s_r_13__86_, s_r_13__85_, s_r_13__84_, s_r_13__83_, s_r_13__82_, s_r_13__81_, s_r_13__80_, s_r_13__79_, s_r_13__78_, s_r_13__77_, s_r_13__76_, s_r_13__75_, s_r_13__74_, s_r_13__73_, s_r_13__72_, s_r_13__71_, s_r_13__70_, s_r_13__69_, s_r_13__68_, s_r_13__67_, s_r_13__66_, s_r_13__65_, s_r_13__64_, s_r_13__63_, s_r_13__62_, s_r_13__61_, s_r_13__60_, s_r_13__59_, s_r_13__58_, s_r_13__57_, s_r_13__56_, s_r_13__55_, s_r_13__54_, s_r_13__53_, s_r_13__52_, s_r_13__51_, s_r_13__50_, s_r_13__49_, s_r_13__48_, s_r_13__47_, s_r_13__46_, s_r_13__45_, s_r_13__44_, s_r_13__43_, s_r_13__42_, s_r_13__41_, s_r_13__40_, s_r_13__39_, s_r_13__38_, s_r_13__37_, s_r_13__36_, s_r_13__35_, s_r_13__34_, s_r_13__33_, s_r_13__32_, s_r_13__31_, s_r_13__30_, s_r_13__29_, s_r_13__28_, s_r_13__27_, s_r_13__26_, s_r_13__25_, s_r_13__24_, s_r_13__23_, s_r_13__22_, s_r_13__21_, s_r_13__20_, s_r_13__19_, s_r_13__18_, s_r_13__17_, s_r_13__16_, s_r_13__15_, s_r_13__14_, s_r_13__13_, s_r_13__12_, s_r_13__11_, s_r_13__10_, s_r_13__9_, s_r_13__8_, s_r_13__7_, s_r_13__6_, s_r_13__5_, s_r_13__4_, s_r_13__3_, s_r_13__2_, s_r_13__1_, s_r_13__0_ }),
    .c_i(c_r[13]),
    .prod_accum_i({ prod_accum_13__14_, prod_accum_13__13_, prod_accum_13__12_, prod_accum_13__11_, prod_accum_13__10_, prod_accum_13__9_, prod_accum_13__8_, prod_accum_13__7_, prod_accum_13__6_, prod_accum_13__5_, prod_accum_13__4_, prod_accum_13__3_, prod_accum_13__2_, prod_accum_13__1_, prod_accum_13__0_ }),
    .a_o(a_r[1919:1792]),
    .b_o(b_r[1919:1792]),
    .s_o({ s_r_14__127_, s_r_14__126_, s_r_14__125_, s_r_14__124_, s_r_14__123_, s_r_14__122_, s_r_14__121_, s_r_14__120_, s_r_14__119_, s_r_14__118_, s_r_14__117_, s_r_14__116_, s_r_14__115_, s_r_14__114_, s_r_14__113_, s_r_14__112_, s_r_14__111_, s_r_14__110_, s_r_14__109_, s_r_14__108_, s_r_14__107_, s_r_14__106_, s_r_14__105_, s_r_14__104_, s_r_14__103_, s_r_14__102_, s_r_14__101_, s_r_14__100_, s_r_14__99_, s_r_14__98_, s_r_14__97_, s_r_14__96_, s_r_14__95_, s_r_14__94_, s_r_14__93_, s_r_14__92_, s_r_14__91_, s_r_14__90_, s_r_14__89_, s_r_14__88_, s_r_14__87_, s_r_14__86_, s_r_14__85_, s_r_14__84_, s_r_14__83_, s_r_14__82_, s_r_14__81_, s_r_14__80_, s_r_14__79_, s_r_14__78_, s_r_14__77_, s_r_14__76_, s_r_14__75_, s_r_14__74_, s_r_14__73_, s_r_14__72_, s_r_14__71_, s_r_14__70_, s_r_14__69_, s_r_14__68_, s_r_14__67_, s_r_14__66_, s_r_14__65_, s_r_14__64_, s_r_14__63_, s_r_14__62_, s_r_14__61_, s_r_14__60_, s_r_14__59_, s_r_14__58_, s_r_14__57_, s_r_14__56_, s_r_14__55_, s_r_14__54_, s_r_14__53_, s_r_14__52_, s_r_14__51_, s_r_14__50_, s_r_14__49_, s_r_14__48_, s_r_14__47_, s_r_14__46_, s_r_14__45_, s_r_14__44_, s_r_14__43_, s_r_14__42_, s_r_14__41_, s_r_14__40_, s_r_14__39_, s_r_14__38_, s_r_14__37_, s_r_14__36_, s_r_14__35_, s_r_14__34_, s_r_14__33_, s_r_14__32_, s_r_14__31_, s_r_14__30_, s_r_14__29_, s_r_14__28_, s_r_14__27_, s_r_14__26_, s_r_14__25_, s_r_14__24_, s_r_14__23_, s_r_14__22_, s_r_14__21_, s_r_14__20_, s_r_14__19_, s_r_14__18_, s_r_14__17_, s_r_14__16_, s_r_14__15_, s_r_14__14_, s_r_14__13_, s_r_14__12_, s_r_14__11_, s_r_14__10_, s_r_14__9_, s_r_14__8_, s_r_14__7_, s_r_14__6_, s_r_14__5_, s_r_14__4_, s_r_14__3_, s_r_14__2_, s_r_14__1_, s_r_14__0_ }),
    .c_o(c_r[14]),
    .prod_accum_o({ prod_accum_14__15_, prod_accum_14__14_, prod_accum_14__13_, prod_accum_14__12_, prod_accum_14__11_, prod_accum_14__10_, prod_accum_14__9_, prod_accum_14__8_, prod_accum_14__7_, prod_accum_14__6_, prod_accum_14__5_, prod_accum_14__4_, prod_accum_14__3_, prod_accum_14__2_, prod_accum_14__1_, prod_accum_14__0_ })
  );


  bsg_mul_array_row_128_15_1
  genblk1_15__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[1919:1792]),
    .b_i(b_r[1919:1792]),
    .s_i({ s_r_14__127_, s_r_14__126_, s_r_14__125_, s_r_14__124_, s_r_14__123_, s_r_14__122_, s_r_14__121_, s_r_14__120_, s_r_14__119_, s_r_14__118_, s_r_14__117_, s_r_14__116_, s_r_14__115_, s_r_14__114_, s_r_14__113_, s_r_14__112_, s_r_14__111_, s_r_14__110_, s_r_14__109_, s_r_14__108_, s_r_14__107_, s_r_14__106_, s_r_14__105_, s_r_14__104_, s_r_14__103_, s_r_14__102_, s_r_14__101_, s_r_14__100_, s_r_14__99_, s_r_14__98_, s_r_14__97_, s_r_14__96_, s_r_14__95_, s_r_14__94_, s_r_14__93_, s_r_14__92_, s_r_14__91_, s_r_14__90_, s_r_14__89_, s_r_14__88_, s_r_14__87_, s_r_14__86_, s_r_14__85_, s_r_14__84_, s_r_14__83_, s_r_14__82_, s_r_14__81_, s_r_14__80_, s_r_14__79_, s_r_14__78_, s_r_14__77_, s_r_14__76_, s_r_14__75_, s_r_14__74_, s_r_14__73_, s_r_14__72_, s_r_14__71_, s_r_14__70_, s_r_14__69_, s_r_14__68_, s_r_14__67_, s_r_14__66_, s_r_14__65_, s_r_14__64_, s_r_14__63_, s_r_14__62_, s_r_14__61_, s_r_14__60_, s_r_14__59_, s_r_14__58_, s_r_14__57_, s_r_14__56_, s_r_14__55_, s_r_14__54_, s_r_14__53_, s_r_14__52_, s_r_14__51_, s_r_14__50_, s_r_14__49_, s_r_14__48_, s_r_14__47_, s_r_14__46_, s_r_14__45_, s_r_14__44_, s_r_14__43_, s_r_14__42_, s_r_14__41_, s_r_14__40_, s_r_14__39_, s_r_14__38_, s_r_14__37_, s_r_14__36_, s_r_14__35_, s_r_14__34_, s_r_14__33_, s_r_14__32_, s_r_14__31_, s_r_14__30_, s_r_14__29_, s_r_14__28_, s_r_14__27_, s_r_14__26_, s_r_14__25_, s_r_14__24_, s_r_14__23_, s_r_14__22_, s_r_14__21_, s_r_14__20_, s_r_14__19_, s_r_14__18_, s_r_14__17_, s_r_14__16_, s_r_14__15_, s_r_14__14_, s_r_14__13_, s_r_14__12_, s_r_14__11_, s_r_14__10_, s_r_14__9_, s_r_14__8_, s_r_14__7_, s_r_14__6_, s_r_14__5_, s_r_14__4_, s_r_14__3_, s_r_14__2_, s_r_14__1_, s_r_14__0_ }),
    .c_i(c_r[14]),
    .prod_accum_i({ prod_accum_14__15_, prod_accum_14__14_, prod_accum_14__13_, prod_accum_14__12_, prod_accum_14__11_, prod_accum_14__10_, prod_accum_14__9_, prod_accum_14__8_, prod_accum_14__7_, prod_accum_14__6_, prod_accum_14__5_, prod_accum_14__4_, prod_accum_14__3_, prod_accum_14__2_, prod_accum_14__1_, prod_accum_14__0_ }),
    .a_o(a_r[2047:1920]),
    .b_o(b_r[2047:1920]),
    .s_o({ s_r_15__127_, s_r_15__126_, s_r_15__125_, s_r_15__124_, s_r_15__123_, s_r_15__122_, s_r_15__121_, s_r_15__120_, s_r_15__119_, s_r_15__118_, s_r_15__117_, s_r_15__116_, s_r_15__115_, s_r_15__114_, s_r_15__113_, s_r_15__112_, s_r_15__111_, s_r_15__110_, s_r_15__109_, s_r_15__108_, s_r_15__107_, s_r_15__106_, s_r_15__105_, s_r_15__104_, s_r_15__103_, s_r_15__102_, s_r_15__101_, s_r_15__100_, s_r_15__99_, s_r_15__98_, s_r_15__97_, s_r_15__96_, s_r_15__95_, s_r_15__94_, s_r_15__93_, s_r_15__92_, s_r_15__91_, s_r_15__90_, s_r_15__89_, s_r_15__88_, s_r_15__87_, s_r_15__86_, s_r_15__85_, s_r_15__84_, s_r_15__83_, s_r_15__82_, s_r_15__81_, s_r_15__80_, s_r_15__79_, s_r_15__78_, s_r_15__77_, s_r_15__76_, s_r_15__75_, s_r_15__74_, s_r_15__73_, s_r_15__72_, s_r_15__71_, s_r_15__70_, s_r_15__69_, s_r_15__68_, s_r_15__67_, s_r_15__66_, s_r_15__65_, s_r_15__64_, s_r_15__63_, s_r_15__62_, s_r_15__61_, s_r_15__60_, s_r_15__59_, s_r_15__58_, s_r_15__57_, s_r_15__56_, s_r_15__55_, s_r_15__54_, s_r_15__53_, s_r_15__52_, s_r_15__51_, s_r_15__50_, s_r_15__49_, s_r_15__48_, s_r_15__47_, s_r_15__46_, s_r_15__45_, s_r_15__44_, s_r_15__43_, s_r_15__42_, s_r_15__41_, s_r_15__40_, s_r_15__39_, s_r_15__38_, s_r_15__37_, s_r_15__36_, s_r_15__35_, s_r_15__34_, s_r_15__33_, s_r_15__32_, s_r_15__31_, s_r_15__30_, s_r_15__29_, s_r_15__28_, s_r_15__27_, s_r_15__26_, s_r_15__25_, s_r_15__24_, s_r_15__23_, s_r_15__22_, s_r_15__21_, s_r_15__20_, s_r_15__19_, s_r_15__18_, s_r_15__17_, s_r_15__16_, s_r_15__15_, s_r_15__14_, s_r_15__13_, s_r_15__12_, s_r_15__11_, s_r_15__10_, s_r_15__9_, s_r_15__8_, s_r_15__7_, s_r_15__6_, s_r_15__5_, s_r_15__4_, s_r_15__3_, s_r_15__2_, s_r_15__1_, s_r_15__0_ }),
    .c_o(c_r[15]),
    .prod_accum_o({ prod_accum_15__16_, prod_accum_15__15_, prod_accum_15__14_, prod_accum_15__13_, prod_accum_15__12_, prod_accum_15__11_, prod_accum_15__10_, prod_accum_15__9_, prod_accum_15__8_, prod_accum_15__7_, prod_accum_15__6_, prod_accum_15__5_, prod_accum_15__4_, prod_accum_15__3_, prod_accum_15__2_, prod_accum_15__1_, prod_accum_15__0_ })
  );


  bsg_mul_array_row_128_16_0
  genblk1_16__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[2047:1920]),
    .b_i(b_r[2047:1920]),
    .s_i({ s_r_15__127_, s_r_15__126_, s_r_15__125_, s_r_15__124_, s_r_15__123_, s_r_15__122_, s_r_15__121_, s_r_15__120_, s_r_15__119_, s_r_15__118_, s_r_15__117_, s_r_15__116_, s_r_15__115_, s_r_15__114_, s_r_15__113_, s_r_15__112_, s_r_15__111_, s_r_15__110_, s_r_15__109_, s_r_15__108_, s_r_15__107_, s_r_15__106_, s_r_15__105_, s_r_15__104_, s_r_15__103_, s_r_15__102_, s_r_15__101_, s_r_15__100_, s_r_15__99_, s_r_15__98_, s_r_15__97_, s_r_15__96_, s_r_15__95_, s_r_15__94_, s_r_15__93_, s_r_15__92_, s_r_15__91_, s_r_15__90_, s_r_15__89_, s_r_15__88_, s_r_15__87_, s_r_15__86_, s_r_15__85_, s_r_15__84_, s_r_15__83_, s_r_15__82_, s_r_15__81_, s_r_15__80_, s_r_15__79_, s_r_15__78_, s_r_15__77_, s_r_15__76_, s_r_15__75_, s_r_15__74_, s_r_15__73_, s_r_15__72_, s_r_15__71_, s_r_15__70_, s_r_15__69_, s_r_15__68_, s_r_15__67_, s_r_15__66_, s_r_15__65_, s_r_15__64_, s_r_15__63_, s_r_15__62_, s_r_15__61_, s_r_15__60_, s_r_15__59_, s_r_15__58_, s_r_15__57_, s_r_15__56_, s_r_15__55_, s_r_15__54_, s_r_15__53_, s_r_15__52_, s_r_15__51_, s_r_15__50_, s_r_15__49_, s_r_15__48_, s_r_15__47_, s_r_15__46_, s_r_15__45_, s_r_15__44_, s_r_15__43_, s_r_15__42_, s_r_15__41_, s_r_15__40_, s_r_15__39_, s_r_15__38_, s_r_15__37_, s_r_15__36_, s_r_15__35_, s_r_15__34_, s_r_15__33_, s_r_15__32_, s_r_15__31_, s_r_15__30_, s_r_15__29_, s_r_15__28_, s_r_15__27_, s_r_15__26_, s_r_15__25_, s_r_15__24_, s_r_15__23_, s_r_15__22_, s_r_15__21_, s_r_15__20_, s_r_15__19_, s_r_15__18_, s_r_15__17_, s_r_15__16_, s_r_15__15_, s_r_15__14_, s_r_15__13_, s_r_15__12_, s_r_15__11_, s_r_15__10_, s_r_15__9_, s_r_15__8_, s_r_15__7_, s_r_15__6_, s_r_15__5_, s_r_15__4_, s_r_15__3_, s_r_15__2_, s_r_15__1_, s_r_15__0_ }),
    .c_i(c_r[15]),
    .prod_accum_i({ prod_accum_15__16_, prod_accum_15__15_, prod_accum_15__14_, prod_accum_15__13_, prod_accum_15__12_, prod_accum_15__11_, prod_accum_15__10_, prod_accum_15__9_, prod_accum_15__8_, prod_accum_15__7_, prod_accum_15__6_, prod_accum_15__5_, prod_accum_15__4_, prod_accum_15__3_, prod_accum_15__2_, prod_accum_15__1_, prod_accum_15__0_ }),
    .a_o(a_r[2175:2048]),
    .b_o(b_r[2175:2048]),
    .s_o({ s_r_16__127_, s_r_16__126_, s_r_16__125_, s_r_16__124_, s_r_16__123_, s_r_16__122_, s_r_16__121_, s_r_16__120_, s_r_16__119_, s_r_16__118_, s_r_16__117_, s_r_16__116_, s_r_16__115_, s_r_16__114_, s_r_16__113_, s_r_16__112_, s_r_16__111_, s_r_16__110_, s_r_16__109_, s_r_16__108_, s_r_16__107_, s_r_16__106_, s_r_16__105_, s_r_16__104_, s_r_16__103_, s_r_16__102_, s_r_16__101_, s_r_16__100_, s_r_16__99_, s_r_16__98_, s_r_16__97_, s_r_16__96_, s_r_16__95_, s_r_16__94_, s_r_16__93_, s_r_16__92_, s_r_16__91_, s_r_16__90_, s_r_16__89_, s_r_16__88_, s_r_16__87_, s_r_16__86_, s_r_16__85_, s_r_16__84_, s_r_16__83_, s_r_16__82_, s_r_16__81_, s_r_16__80_, s_r_16__79_, s_r_16__78_, s_r_16__77_, s_r_16__76_, s_r_16__75_, s_r_16__74_, s_r_16__73_, s_r_16__72_, s_r_16__71_, s_r_16__70_, s_r_16__69_, s_r_16__68_, s_r_16__67_, s_r_16__66_, s_r_16__65_, s_r_16__64_, s_r_16__63_, s_r_16__62_, s_r_16__61_, s_r_16__60_, s_r_16__59_, s_r_16__58_, s_r_16__57_, s_r_16__56_, s_r_16__55_, s_r_16__54_, s_r_16__53_, s_r_16__52_, s_r_16__51_, s_r_16__50_, s_r_16__49_, s_r_16__48_, s_r_16__47_, s_r_16__46_, s_r_16__45_, s_r_16__44_, s_r_16__43_, s_r_16__42_, s_r_16__41_, s_r_16__40_, s_r_16__39_, s_r_16__38_, s_r_16__37_, s_r_16__36_, s_r_16__35_, s_r_16__34_, s_r_16__33_, s_r_16__32_, s_r_16__31_, s_r_16__30_, s_r_16__29_, s_r_16__28_, s_r_16__27_, s_r_16__26_, s_r_16__25_, s_r_16__24_, s_r_16__23_, s_r_16__22_, s_r_16__21_, s_r_16__20_, s_r_16__19_, s_r_16__18_, s_r_16__17_, s_r_16__16_, s_r_16__15_, s_r_16__14_, s_r_16__13_, s_r_16__12_, s_r_16__11_, s_r_16__10_, s_r_16__9_, s_r_16__8_, s_r_16__7_, s_r_16__6_, s_r_16__5_, s_r_16__4_, s_r_16__3_, s_r_16__2_, s_r_16__1_, s_r_16__0_ }),
    .c_o(c_r[16]),
    .prod_accum_o({ prod_accum_16__17_, prod_accum_16__16_, prod_accum_16__15_, prod_accum_16__14_, prod_accum_16__13_, prod_accum_16__12_, prod_accum_16__11_, prod_accum_16__10_, prod_accum_16__9_, prod_accum_16__8_, prod_accum_16__7_, prod_accum_16__6_, prod_accum_16__5_, prod_accum_16__4_, prod_accum_16__3_, prod_accum_16__2_, prod_accum_16__1_, prod_accum_16__0_ })
  );


  bsg_mul_array_row_128_17_0
  genblk1_17__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[2175:2048]),
    .b_i(b_r[2175:2048]),
    .s_i({ s_r_16__127_, s_r_16__126_, s_r_16__125_, s_r_16__124_, s_r_16__123_, s_r_16__122_, s_r_16__121_, s_r_16__120_, s_r_16__119_, s_r_16__118_, s_r_16__117_, s_r_16__116_, s_r_16__115_, s_r_16__114_, s_r_16__113_, s_r_16__112_, s_r_16__111_, s_r_16__110_, s_r_16__109_, s_r_16__108_, s_r_16__107_, s_r_16__106_, s_r_16__105_, s_r_16__104_, s_r_16__103_, s_r_16__102_, s_r_16__101_, s_r_16__100_, s_r_16__99_, s_r_16__98_, s_r_16__97_, s_r_16__96_, s_r_16__95_, s_r_16__94_, s_r_16__93_, s_r_16__92_, s_r_16__91_, s_r_16__90_, s_r_16__89_, s_r_16__88_, s_r_16__87_, s_r_16__86_, s_r_16__85_, s_r_16__84_, s_r_16__83_, s_r_16__82_, s_r_16__81_, s_r_16__80_, s_r_16__79_, s_r_16__78_, s_r_16__77_, s_r_16__76_, s_r_16__75_, s_r_16__74_, s_r_16__73_, s_r_16__72_, s_r_16__71_, s_r_16__70_, s_r_16__69_, s_r_16__68_, s_r_16__67_, s_r_16__66_, s_r_16__65_, s_r_16__64_, s_r_16__63_, s_r_16__62_, s_r_16__61_, s_r_16__60_, s_r_16__59_, s_r_16__58_, s_r_16__57_, s_r_16__56_, s_r_16__55_, s_r_16__54_, s_r_16__53_, s_r_16__52_, s_r_16__51_, s_r_16__50_, s_r_16__49_, s_r_16__48_, s_r_16__47_, s_r_16__46_, s_r_16__45_, s_r_16__44_, s_r_16__43_, s_r_16__42_, s_r_16__41_, s_r_16__40_, s_r_16__39_, s_r_16__38_, s_r_16__37_, s_r_16__36_, s_r_16__35_, s_r_16__34_, s_r_16__33_, s_r_16__32_, s_r_16__31_, s_r_16__30_, s_r_16__29_, s_r_16__28_, s_r_16__27_, s_r_16__26_, s_r_16__25_, s_r_16__24_, s_r_16__23_, s_r_16__22_, s_r_16__21_, s_r_16__20_, s_r_16__19_, s_r_16__18_, s_r_16__17_, s_r_16__16_, s_r_16__15_, s_r_16__14_, s_r_16__13_, s_r_16__12_, s_r_16__11_, s_r_16__10_, s_r_16__9_, s_r_16__8_, s_r_16__7_, s_r_16__6_, s_r_16__5_, s_r_16__4_, s_r_16__3_, s_r_16__2_, s_r_16__1_, s_r_16__0_ }),
    .c_i(c_r[16]),
    .prod_accum_i({ prod_accum_16__17_, prod_accum_16__16_, prod_accum_16__15_, prod_accum_16__14_, prod_accum_16__13_, prod_accum_16__12_, prod_accum_16__11_, prod_accum_16__10_, prod_accum_16__9_, prod_accum_16__8_, prod_accum_16__7_, prod_accum_16__6_, prod_accum_16__5_, prod_accum_16__4_, prod_accum_16__3_, prod_accum_16__2_, prod_accum_16__1_, prod_accum_16__0_ }),
    .a_o(a_r[2303:2176]),
    .b_o(b_r[2303:2176]),
    .s_o({ s_r_17__127_, s_r_17__126_, s_r_17__125_, s_r_17__124_, s_r_17__123_, s_r_17__122_, s_r_17__121_, s_r_17__120_, s_r_17__119_, s_r_17__118_, s_r_17__117_, s_r_17__116_, s_r_17__115_, s_r_17__114_, s_r_17__113_, s_r_17__112_, s_r_17__111_, s_r_17__110_, s_r_17__109_, s_r_17__108_, s_r_17__107_, s_r_17__106_, s_r_17__105_, s_r_17__104_, s_r_17__103_, s_r_17__102_, s_r_17__101_, s_r_17__100_, s_r_17__99_, s_r_17__98_, s_r_17__97_, s_r_17__96_, s_r_17__95_, s_r_17__94_, s_r_17__93_, s_r_17__92_, s_r_17__91_, s_r_17__90_, s_r_17__89_, s_r_17__88_, s_r_17__87_, s_r_17__86_, s_r_17__85_, s_r_17__84_, s_r_17__83_, s_r_17__82_, s_r_17__81_, s_r_17__80_, s_r_17__79_, s_r_17__78_, s_r_17__77_, s_r_17__76_, s_r_17__75_, s_r_17__74_, s_r_17__73_, s_r_17__72_, s_r_17__71_, s_r_17__70_, s_r_17__69_, s_r_17__68_, s_r_17__67_, s_r_17__66_, s_r_17__65_, s_r_17__64_, s_r_17__63_, s_r_17__62_, s_r_17__61_, s_r_17__60_, s_r_17__59_, s_r_17__58_, s_r_17__57_, s_r_17__56_, s_r_17__55_, s_r_17__54_, s_r_17__53_, s_r_17__52_, s_r_17__51_, s_r_17__50_, s_r_17__49_, s_r_17__48_, s_r_17__47_, s_r_17__46_, s_r_17__45_, s_r_17__44_, s_r_17__43_, s_r_17__42_, s_r_17__41_, s_r_17__40_, s_r_17__39_, s_r_17__38_, s_r_17__37_, s_r_17__36_, s_r_17__35_, s_r_17__34_, s_r_17__33_, s_r_17__32_, s_r_17__31_, s_r_17__30_, s_r_17__29_, s_r_17__28_, s_r_17__27_, s_r_17__26_, s_r_17__25_, s_r_17__24_, s_r_17__23_, s_r_17__22_, s_r_17__21_, s_r_17__20_, s_r_17__19_, s_r_17__18_, s_r_17__17_, s_r_17__16_, s_r_17__15_, s_r_17__14_, s_r_17__13_, s_r_17__12_, s_r_17__11_, s_r_17__10_, s_r_17__9_, s_r_17__8_, s_r_17__7_, s_r_17__6_, s_r_17__5_, s_r_17__4_, s_r_17__3_, s_r_17__2_, s_r_17__1_, s_r_17__0_ }),
    .c_o(c_r[17]),
    .prod_accum_o({ prod_accum_17__18_, prod_accum_17__17_, prod_accum_17__16_, prod_accum_17__15_, prod_accum_17__14_, prod_accum_17__13_, prod_accum_17__12_, prod_accum_17__11_, prod_accum_17__10_, prod_accum_17__9_, prod_accum_17__8_, prod_accum_17__7_, prod_accum_17__6_, prod_accum_17__5_, prod_accum_17__4_, prod_accum_17__3_, prod_accum_17__2_, prod_accum_17__1_, prod_accum_17__0_ })
  );


  bsg_mul_array_row_128_18_0
  genblk1_18__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[2303:2176]),
    .b_i(b_r[2303:2176]),
    .s_i({ s_r_17__127_, s_r_17__126_, s_r_17__125_, s_r_17__124_, s_r_17__123_, s_r_17__122_, s_r_17__121_, s_r_17__120_, s_r_17__119_, s_r_17__118_, s_r_17__117_, s_r_17__116_, s_r_17__115_, s_r_17__114_, s_r_17__113_, s_r_17__112_, s_r_17__111_, s_r_17__110_, s_r_17__109_, s_r_17__108_, s_r_17__107_, s_r_17__106_, s_r_17__105_, s_r_17__104_, s_r_17__103_, s_r_17__102_, s_r_17__101_, s_r_17__100_, s_r_17__99_, s_r_17__98_, s_r_17__97_, s_r_17__96_, s_r_17__95_, s_r_17__94_, s_r_17__93_, s_r_17__92_, s_r_17__91_, s_r_17__90_, s_r_17__89_, s_r_17__88_, s_r_17__87_, s_r_17__86_, s_r_17__85_, s_r_17__84_, s_r_17__83_, s_r_17__82_, s_r_17__81_, s_r_17__80_, s_r_17__79_, s_r_17__78_, s_r_17__77_, s_r_17__76_, s_r_17__75_, s_r_17__74_, s_r_17__73_, s_r_17__72_, s_r_17__71_, s_r_17__70_, s_r_17__69_, s_r_17__68_, s_r_17__67_, s_r_17__66_, s_r_17__65_, s_r_17__64_, s_r_17__63_, s_r_17__62_, s_r_17__61_, s_r_17__60_, s_r_17__59_, s_r_17__58_, s_r_17__57_, s_r_17__56_, s_r_17__55_, s_r_17__54_, s_r_17__53_, s_r_17__52_, s_r_17__51_, s_r_17__50_, s_r_17__49_, s_r_17__48_, s_r_17__47_, s_r_17__46_, s_r_17__45_, s_r_17__44_, s_r_17__43_, s_r_17__42_, s_r_17__41_, s_r_17__40_, s_r_17__39_, s_r_17__38_, s_r_17__37_, s_r_17__36_, s_r_17__35_, s_r_17__34_, s_r_17__33_, s_r_17__32_, s_r_17__31_, s_r_17__30_, s_r_17__29_, s_r_17__28_, s_r_17__27_, s_r_17__26_, s_r_17__25_, s_r_17__24_, s_r_17__23_, s_r_17__22_, s_r_17__21_, s_r_17__20_, s_r_17__19_, s_r_17__18_, s_r_17__17_, s_r_17__16_, s_r_17__15_, s_r_17__14_, s_r_17__13_, s_r_17__12_, s_r_17__11_, s_r_17__10_, s_r_17__9_, s_r_17__8_, s_r_17__7_, s_r_17__6_, s_r_17__5_, s_r_17__4_, s_r_17__3_, s_r_17__2_, s_r_17__1_, s_r_17__0_ }),
    .c_i(c_r[17]),
    .prod_accum_i({ prod_accum_17__18_, prod_accum_17__17_, prod_accum_17__16_, prod_accum_17__15_, prod_accum_17__14_, prod_accum_17__13_, prod_accum_17__12_, prod_accum_17__11_, prod_accum_17__10_, prod_accum_17__9_, prod_accum_17__8_, prod_accum_17__7_, prod_accum_17__6_, prod_accum_17__5_, prod_accum_17__4_, prod_accum_17__3_, prod_accum_17__2_, prod_accum_17__1_, prod_accum_17__0_ }),
    .a_o(a_r[2431:2304]),
    .b_o(b_r[2431:2304]),
    .s_o({ s_r_18__127_, s_r_18__126_, s_r_18__125_, s_r_18__124_, s_r_18__123_, s_r_18__122_, s_r_18__121_, s_r_18__120_, s_r_18__119_, s_r_18__118_, s_r_18__117_, s_r_18__116_, s_r_18__115_, s_r_18__114_, s_r_18__113_, s_r_18__112_, s_r_18__111_, s_r_18__110_, s_r_18__109_, s_r_18__108_, s_r_18__107_, s_r_18__106_, s_r_18__105_, s_r_18__104_, s_r_18__103_, s_r_18__102_, s_r_18__101_, s_r_18__100_, s_r_18__99_, s_r_18__98_, s_r_18__97_, s_r_18__96_, s_r_18__95_, s_r_18__94_, s_r_18__93_, s_r_18__92_, s_r_18__91_, s_r_18__90_, s_r_18__89_, s_r_18__88_, s_r_18__87_, s_r_18__86_, s_r_18__85_, s_r_18__84_, s_r_18__83_, s_r_18__82_, s_r_18__81_, s_r_18__80_, s_r_18__79_, s_r_18__78_, s_r_18__77_, s_r_18__76_, s_r_18__75_, s_r_18__74_, s_r_18__73_, s_r_18__72_, s_r_18__71_, s_r_18__70_, s_r_18__69_, s_r_18__68_, s_r_18__67_, s_r_18__66_, s_r_18__65_, s_r_18__64_, s_r_18__63_, s_r_18__62_, s_r_18__61_, s_r_18__60_, s_r_18__59_, s_r_18__58_, s_r_18__57_, s_r_18__56_, s_r_18__55_, s_r_18__54_, s_r_18__53_, s_r_18__52_, s_r_18__51_, s_r_18__50_, s_r_18__49_, s_r_18__48_, s_r_18__47_, s_r_18__46_, s_r_18__45_, s_r_18__44_, s_r_18__43_, s_r_18__42_, s_r_18__41_, s_r_18__40_, s_r_18__39_, s_r_18__38_, s_r_18__37_, s_r_18__36_, s_r_18__35_, s_r_18__34_, s_r_18__33_, s_r_18__32_, s_r_18__31_, s_r_18__30_, s_r_18__29_, s_r_18__28_, s_r_18__27_, s_r_18__26_, s_r_18__25_, s_r_18__24_, s_r_18__23_, s_r_18__22_, s_r_18__21_, s_r_18__20_, s_r_18__19_, s_r_18__18_, s_r_18__17_, s_r_18__16_, s_r_18__15_, s_r_18__14_, s_r_18__13_, s_r_18__12_, s_r_18__11_, s_r_18__10_, s_r_18__9_, s_r_18__8_, s_r_18__7_, s_r_18__6_, s_r_18__5_, s_r_18__4_, s_r_18__3_, s_r_18__2_, s_r_18__1_, s_r_18__0_ }),
    .c_o(c_r[18]),
    .prod_accum_o({ prod_accum_18__19_, prod_accum_18__18_, prod_accum_18__17_, prod_accum_18__16_, prod_accum_18__15_, prod_accum_18__14_, prod_accum_18__13_, prod_accum_18__12_, prod_accum_18__11_, prod_accum_18__10_, prod_accum_18__9_, prod_accum_18__8_, prod_accum_18__7_, prod_accum_18__6_, prod_accum_18__5_, prod_accum_18__4_, prod_accum_18__3_, prod_accum_18__2_, prod_accum_18__1_, prod_accum_18__0_ })
  );


  bsg_mul_array_row_128_19_0
  genblk1_19__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[2431:2304]),
    .b_i(b_r[2431:2304]),
    .s_i({ s_r_18__127_, s_r_18__126_, s_r_18__125_, s_r_18__124_, s_r_18__123_, s_r_18__122_, s_r_18__121_, s_r_18__120_, s_r_18__119_, s_r_18__118_, s_r_18__117_, s_r_18__116_, s_r_18__115_, s_r_18__114_, s_r_18__113_, s_r_18__112_, s_r_18__111_, s_r_18__110_, s_r_18__109_, s_r_18__108_, s_r_18__107_, s_r_18__106_, s_r_18__105_, s_r_18__104_, s_r_18__103_, s_r_18__102_, s_r_18__101_, s_r_18__100_, s_r_18__99_, s_r_18__98_, s_r_18__97_, s_r_18__96_, s_r_18__95_, s_r_18__94_, s_r_18__93_, s_r_18__92_, s_r_18__91_, s_r_18__90_, s_r_18__89_, s_r_18__88_, s_r_18__87_, s_r_18__86_, s_r_18__85_, s_r_18__84_, s_r_18__83_, s_r_18__82_, s_r_18__81_, s_r_18__80_, s_r_18__79_, s_r_18__78_, s_r_18__77_, s_r_18__76_, s_r_18__75_, s_r_18__74_, s_r_18__73_, s_r_18__72_, s_r_18__71_, s_r_18__70_, s_r_18__69_, s_r_18__68_, s_r_18__67_, s_r_18__66_, s_r_18__65_, s_r_18__64_, s_r_18__63_, s_r_18__62_, s_r_18__61_, s_r_18__60_, s_r_18__59_, s_r_18__58_, s_r_18__57_, s_r_18__56_, s_r_18__55_, s_r_18__54_, s_r_18__53_, s_r_18__52_, s_r_18__51_, s_r_18__50_, s_r_18__49_, s_r_18__48_, s_r_18__47_, s_r_18__46_, s_r_18__45_, s_r_18__44_, s_r_18__43_, s_r_18__42_, s_r_18__41_, s_r_18__40_, s_r_18__39_, s_r_18__38_, s_r_18__37_, s_r_18__36_, s_r_18__35_, s_r_18__34_, s_r_18__33_, s_r_18__32_, s_r_18__31_, s_r_18__30_, s_r_18__29_, s_r_18__28_, s_r_18__27_, s_r_18__26_, s_r_18__25_, s_r_18__24_, s_r_18__23_, s_r_18__22_, s_r_18__21_, s_r_18__20_, s_r_18__19_, s_r_18__18_, s_r_18__17_, s_r_18__16_, s_r_18__15_, s_r_18__14_, s_r_18__13_, s_r_18__12_, s_r_18__11_, s_r_18__10_, s_r_18__9_, s_r_18__8_, s_r_18__7_, s_r_18__6_, s_r_18__5_, s_r_18__4_, s_r_18__3_, s_r_18__2_, s_r_18__1_, s_r_18__0_ }),
    .c_i(c_r[18]),
    .prod_accum_i({ prod_accum_18__19_, prod_accum_18__18_, prod_accum_18__17_, prod_accum_18__16_, prod_accum_18__15_, prod_accum_18__14_, prod_accum_18__13_, prod_accum_18__12_, prod_accum_18__11_, prod_accum_18__10_, prod_accum_18__9_, prod_accum_18__8_, prod_accum_18__7_, prod_accum_18__6_, prod_accum_18__5_, prod_accum_18__4_, prod_accum_18__3_, prod_accum_18__2_, prod_accum_18__1_, prod_accum_18__0_ }),
    .a_o(a_r[2559:2432]),
    .b_o(b_r[2559:2432]),
    .s_o({ s_r_19__127_, s_r_19__126_, s_r_19__125_, s_r_19__124_, s_r_19__123_, s_r_19__122_, s_r_19__121_, s_r_19__120_, s_r_19__119_, s_r_19__118_, s_r_19__117_, s_r_19__116_, s_r_19__115_, s_r_19__114_, s_r_19__113_, s_r_19__112_, s_r_19__111_, s_r_19__110_, s_r_19__109_, s_r_19__108_, s_r_19__107_, s_r_19__106_, s_r_19__105_, s_r_19__104_, s_r_19__103_, s_r_19__102_, s_r_19__101_, s_r_19__100_, s_r_19__99_, s_r_19__98_, s_r_19__97_, s_r_19__96_, s_r_19__95_, s_r_19__94_, s_r_19__93_, s_r_19__92_, s_r_19__91_, s_r_19__90_, s_r_19__89_, s_r_19__88_, s_r_19__87_, s_r_19__86_, s_r_19__85_, s_r_19__84_, s_r_19__83_, s_r_19__82_, s_r_19__81_, s_r_19__80_, s_r_19__79_, s_r_19__78_, s_r_19__77_, s_r_19__76_, s_r_19__75_, s_r_19__74_, s_r_19__73_, s_r_19__72_, s_r_19__71_, s_r_19__70_, s_r_19__69_, s_r_19__68_, s_r_19__67_, s_r_19__66_, s_r_19__65_, s_r_19__64_, s_r_19__63_, s_r_19__62_, s_r_19__61_, s_r_19__60_, s_r_19__59_, s_r_19__58_, s_r_19__57_, s_r_19__56_, s_r_19__55_, s_r_19__54_, s_r_19__53_, s_r_19__52_, s_r_19__51_, s_r_19__50_, s_r_19__49_, s_r_19__48_, s_r_19__47_, s_r_19__46_, s_r_19__45_, s_r_19__44_, s_r_19__43_, s_r_19__42_, s_r_19__41_, s_r_19__40_, s_r_19__39_, s_r_19__38_, s_r_19__37_, s_r_19__36_, s_r_19__35_, s_r_19__34_, s_r_19__33_, s_r_19__32_, s_r_19__31_, s_r_19__30_, s_r_19__29_, s_r_19__28_, s_r_19__27_, s_r_19__26_, s_r_19__25_, s_r_19__24_, s_r_19__23_, s_r_19__22_, s_r_19__21_, s_r_19__20_, s_r_19__19_, s_r_19__18_, s_r_19__17_, s_r_19__16_, s_r_19__15_, s_r_19__14_, s_r_19__13_, s_r_19__12_, s_r_19__11_, s_r_19__10_, s_r_19__9_, s_r_19__8_, s_r_19__7_, s_r_19__6_, s_r_19__5_, s_r_19__4_, s_r_19__3_, s_r_19__2_, s_r_19__1_, s_r_19__0_ }),
    .c_o(c_r[19]),
    .prod_accum_o({ prod_accum_19__20_, prod_accum_19__19_, prod_accum_19__18_, prod_accum_19__17_, prod_accum_19__16_, prod_accum_19__15_, prod_accum_19__14_, prod_accum_19__13_, prod_accum_19__12_, prod_accum_19__11_, prod_accum_19__10_, prod_accum_19__9_, prod_accum_19__8_, prod_accum_19__7_, prod_accum_19__6_, prod_accum_19__5_, prod_accum_19__4_, prod_accum_19__3_, prod_accum_19__2_, prod_accum_19__1_, prod_accum_19__0_ })
  );


  bsg_mul_array_row_128_20_0
  genblk1_20__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[2559:2432]),
    .b_i(b_r[2559:2432]),
    .s_i({ s_r_19__127_, s_r_19__126_, s_r_19__125_, s_r_19__124_, s_r_19__123_, s_r_19__122_, s_r_19__121_, s_r_19__120_, s_r_19__119_, s_r_19__118_, s_r_19__117_, s_r_19__116_, s_r_19__115_, s_r_19__114_, s_r_19__113_, s_r_19__112_, s_r_19__111_, s_r_19__110_, s_r_19__109_, s_r_19__108_, s_r_19__107_, s_r_19__106_, s_r_19__105_, s_r_19__104_, s_r_19__103_, s_r_19__102_, s_r_19__101_, s_r_19__100_, s_r_19__99_, s_r_19__98_, s_r_19__97_, s_r_19__96_, s_r_19__95_, s_r_19__94_, s_r_19__93_, s_r_19__92_, s_r_19__91_, s_r_19__90_, s_r_19__89_, s_r_19__88_, s_r_19__87_, s_r_19__86_, s_r_19__85_, s_r_19__84_, s_r_19__83_, s_r_19__82_, s_r_19__81_, s_r_19__80_, s_r_19__79_, s_r_19__78_, s_r_19__77_, s_r_19__76_, s_r_19__75_, s_r_19__74_, s_r_19__73_, s_r_19__72_, s_r_19__71_, s_r_19__70_, s_r_19__69_, s_r_19__68_, s_r_19__67_, s_r_19__66_, s_r_19__65_, s_r_19__64_, s_r_19__63_, s_r_19__62_, s_r_19__61_, s_r_19__60_, s_r_19__59_, s_r_19__58_, s_r_19__57_, s_r_19__56_, s_r_19__55_, s_r_19__54_, s_r_19__53_, s_r_19__52_, s_r_19__51_, s_r_19__50_, s_r_19__49_, s_r_19__48_, s_r_19__47_, s_r_19__46_, s_r_19__45_, s_r_19__44_, s_r_19__43_, s_r_19__42_, s_r_19__41_, s_r_19__40_, s_r_19__39_, s_r_19__38_, s_r_19__37_, s_r_19__36_, s_r_19__35_, s_r_19__34_, s_r_19__33_, s_r_19__32_, s_r_19__31_, s_r_19__30_, s_r_19__29_, s_r_19__28_, s_r_19__27_, s_r_19__26_, s_r_19__25_, s_r_19__24_, s_r_19__23_, s_r_19__22_, s_r_19__21_, s_r_19__20_, s_r_19__19_, s_r_19__18_, s_r_19__17_, s_r_19__16_, s_r_19__15_, s_r_19__14_, s_r_19__13_, s_r_19__12_, s_r_19__11_, s_r_19__10_, s_r_19__9_, s_r_19__8_, s_r_19__7_, s_r_19__6_, s_r_19__5_, s_r_19__4_, s_r_19__3_, s_r_19__2_, s_r_19__1_, s_r_19__0_ }),
    .c_i(c_r[19]),
    .prod_accum_i({ prod_accum_19__20_, prod_accum_19__19_, prod_accum_19__18_, prod_accum_19__17_, prod_accum_19__16_, prod_accum_19__15_, prod_accum_19__14_, prod_accum_19__13_, prod_accum_19__12_, prod_accum_19__11_, prod_accum_19__10_, prod_accum_19__9_, prod_accum_19__8_, prod_accum_19__7_, prod_accum_19__6_, prod_accum_19__5_, prod_accum_19__4_, prod_accum_19__3_, prod_accum_19__2_, prod_accum_19__1_, prod_accum_19__0_ }),
    .a_o(a_r[2687:2560]),
    .b_o(b_r[2687:2560]),
    .s_o({ s_r_20__127_, s_r_20__126_, s_r_20__125_, s_r_20__124_, s_r_20__123_, s_r_20__122_, s_r_20__121_, s_r_20__120_, s_r_20__119_, s_r_20__118_, s_r_20__117_, s_r_20__116_, s_r_20__115_, s_r_20__114_, s_r_20__113_, s_r_20__112_, s_r_20__111_, s_r_20__110_, s_r_20__109_, s_r_20__108_, s_r_20__107_, s_r_20__106_, s_r_20__105_, s_r_20__104_, s_r_20__103_, s_r_20__102_, s_r_20__101_, s_r_20__100_, s_r_20__99_, s_r_20__98_, s_r_20__97_, s_r_20__96_, s_r_20__95_, s_r_20__94_, s_r_20__93_, s_r_20__92_, s_r_20__91_, s_r_20__90_, s_r_20__89_, s_r_20__88_, s_r_20__87_, s_r_20__86_, s_r_20__85_, s_r_20__84_, s_r_20__83_, s_r_20__82_, s_r_20__81_, s_r_20__80_, s_r_20__79_, s_r_20__78_, s_r_20__77_, s_r_20__76_, s_r_20__75_, s_r_20__74_, s_r_20__73_, s_r_20__72_, s_r_20__71_, s_r_20__70_, s_r_20__69_, s_r_20__68_, s_r_20__67_, s_r_20__66_, s_r_20__65_, s_r_20__64_, s_r_20__63_, s_r_20__62_, s_r_20__61_, s_r_20__60_, s_r_20__59_, s_r_20__58_, s_r_20__57_, s_r_20__56_, s_r_20__55_, s_r_20__54_, s_r_20__53_, s_r_20__52_, s_r_20__51_, s_r_20__50_, s_r_20__49_, s_r_20__48_, s_r_20__47_, s_r_20__46_, s_r_20__45_, s_r_20__44_, s_r_20__43_, s_r_20__42_, s_r_20__41_, s_r_20__40_, s_r_20__39_, s_r_20__38_, s_r_20__37_, s_r_20__36_, s_r_20__35_, s_r_20__34_, s_r_20__33_, s_r_20__32_, s_r_20__31_, s_r_20__30_, s_r_20__29_, s_r_20__28_, s_r_20__27_, s_r_20__26_, s_r_20__25_, s_r_20__24_, s_r_20__23_, s_r_20__22_, s_r_20__21_, s_r_20__20_, s_r_20__19_, s_r_20__18_, s_r_20__17_, s_r_20__16_, s_r_20__15_, s_r_20__14_, s_r_20__13_, s_r_20__12_, s_r_20__11_, s_r_20__10_, s_r_20__9_, s_r_20__8_, s_r_20__7_, s_r_20__6_, s_r_20__5_, s_r_20__4_, s_r_20__3_, s_r_20__2_, s_r_20__1_, s_r_20__0_ }),
    .c_o(c_r[20]),
    .prod_accum_o({ prod_accum_20__21_, prod_accum_20__20_, prod_accum_20__19_, prod_accum_20__18_, prod_accum_20__17_, prod_accum_20__16_, prod_accum_20__15_, prod_accum_20__14_, prod_accum_20__13_, prod_accum_20__12_, prod_accum_20__11_, prod_accum_20__10_, prod_accum_20__9_, prod_accum_20__8_, prod_accum_20__7_, prod_accum_20__6_, prod_accum_20__5_, prod_accum_20__4_, prod_accum_20__3_, prod_accum_20__2_, prod_accum_20__1_, prod_accum_20__0_ })
  );


  bsg_mul_array_row_128_21_0
  genblk1_21__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[2687:2560]),
    .b_i(b_r[2687:2560]),
    .s_i({ s_r_20__127_, s_r_20__126_, s_r_20__125_, s_r_20__124_, s_r_20__123_, s_r_20__122_, s_r_20__121_, s_r_20__120_, s_r_20__119_, s_r_20__118_, s_r_20__117_, s_r_20__116_, s_r_20__115_, s_r_20__114_, s_r_20__113_, s_r_20__112_, s_r_20__111_, s_r_20__110_, s_r_20__109_, s_r_20__108_, s_r_20__107_, s_r_20__106_, s_r_20__105_, s_r_20__104_, s_r_20__103_, s_r_20__102_, s_r_20__101_, s_r_20__100_, s_r_20__99_, s_r_20__98_, s_r_20__97_, s_r_20__96_, s_r_20__95_, s_r_20__94_, s_r_20__93_, s_r_20__92_, s_r_20__91_, s_r_20__90_, s_r_20__89_, s_r_20__88_, s_r_20__87_, s_r_20__86_, s_r_20__85_, s_r_20__84_, s_r_20__83_, s_r_20__82_, s_r_20__81_, s_r_20__80_, s_r_20__79_, s_r_20__78_, s_r_20__77_, s_r_20__76_, s_r_20__75_, s_r_20__74_, s_r_20__73_, s_r_20__72_, s_r_20__71_, s_r_20__70_, s_r_20__69_, s_r_20__68_, s_r_20__67_, s_r_20__66_, s_r_20__65_, s_r_20__64_, s_r_20__63_, s_r_20__62_, s_r_20__61_, s_r_20__60_, s_r_20__59_, s_r_20__58_, s_r_20__57_, s_r_20__56_, s_r_20__55_, s_r_20__54_, s_r_20__53_, s_r_20__52_, s_r_20__51_, s_r_20__50_, s_r_20__49_, s_r_20__48_, s_r_20__47_, s_r_20__46_, s_r_20__45_, s_r_20__44_, s_r_20__43_, s_r_20__42_, s_r_20__41_, s_r_20__40_, s_r_20__39_, s_r_20__38_, s_r_20__37_, s_r_20__36_, s_r_20__35_, s_r_20__34_, s_r_20__33_, s_r_20__32_, s_r_20__31_, s_r_20__30_, s_r_20__29_, s_r_20__28_, s_r_20__27_, s_r_20__26_, s_r_20__25_, s_r_20__24_, s_r_20__23_, s_r_20__22_, s_r_20__21_, s_r_20__20_, s_r_20__19_, s_r_20__18_, s_r_20__17_, s_r_20__16_, s_r_20__15_, s_r_20__14_, s_r_20__13_, s_r_20__12_, s_r_20__11_, s_r_20__10_, s_r_20__9_, s_r_20__8_, s_r_20__7_, s_r_20__6_, s_r_20__5_, s_r_20__4_, s_r_20__3_, s_r_20__2_, s_r_20__1_, s_r_20__0_ }),
    .c_i(c_r[20]),
    .prod_accum_i({ prod_accum_20__21_, prod_accum_20__20_, prod_accum_20__19_, prod_accum_20__18_, prod_accum_20__17_, prod_accum_20__16_, prod_accum_20__15_, prod_accum_20__14_, prod_accum_20__13_, prod_accum_20__12_, prod_accum_20__11_, prod_accum_20__10_, prod_accum_20__9_, prod_accum_20__8_, prod_accum_20__7_, prod_accum_20__6_, prod_accum_20__5_, prod_accum_20__4_, prod_accum_20__3_, prod_accum_20__2_, prod_accum_20__1_, prod_accum_20__0_ }),
    .a_o(a_r[2815:2688]),
    .b_o(b_r[2815:2688]),
    .s_o({ s_r_21__127_, s_r_21__126_, s_r_21__125_, s_r_21__124_, s_r_21__123_, s_r_21__122_, s_r_21__121_, s_r_21__120_, s_r_21__119_, s_r_21__118_, s_r_21__117_, s_r_21__116_, s_r_21__115_, s_r_21__114_, s_r_21__113_, s_r_21__112_, s_r_21__111_, s_r_21__110_, s_r_21__109_, s_r_21__108_, s_r_21__107_, s_r_21__106_, s_r_21__105_, s_r_21__104_, s_r_21__103_, s_r_21__102_, s_r_21__101_, s_r_21__100_, s_r_21__99_, s_r_21__98_, s_r_21__97_, s_r_21__96_, s_r_21__95_, s_r_21__94_, s_r_21__93_, s_r_21__92_, s_r_21__91_, s_r_21__90_, s_r_21__89_, s_r_21__88_, s_r_21__87_, s_r_21__86_, s_r_21__85_, s_r_21__84_, s_r_21__83_, s_r_21__82_, s_r_21__81_, s_r_21__80_, s_r_21__79_, s_r_21__78_, s_r_21__77_, s_r_21__76_, s_r_21__75_, s_r_21__74_, s_r_21__73_, s_r_21__72_, s_r_21__71_, s_r_21__70_, s_r_21__69_, s_r_21__68_, s_r_21__67_, s_r_21__66_, s_r_21__65_, s_r_21__64_, s_r_21__63_, s_r_21__62_, s_r_21__61_, s_r_21__60_, s_r_21__59_, s_r_21__58_, s_r_21__57_, s_r_21__56_, s_r_21__55_, s_r_21__54_, s_r_21__53_, s_r_21__52_, s_r_21__51_, s_r_21__50_, s_r_21__49_, s_r_21__48_, s_r_21__47_, s_r_21__46_, s_r_21__45_, s_r_21__44_, s_r_21__43_, s_r_21__42_, s_r_21__41_, s_r_21__40_, s_r_21__39_, s_r_21__38_, s_r_21__37_, s_r_21__36_, s_r_21__35_, s_r_21__34_, s_r_21__33_, s_r_21__32_, s_r_21__31_, s_r_21__30_, s_r_21__29_, s_r_21__28_, s_r_21__27_, s_r_21__26_, s_r_21__25_, s_r_21__24_, s_r_21__23_, s_r_21__22_, s_r_21__21_, s_r_21__20_, s_r_21__19_, s_r_21__18_, s_r_21__17_, s_r_21__16_, s_r_21__15_, s_r_21__14_, s_r_21__13_, s_r_21__12_, s_r_21__11_, s_r_21__10_, s_r_21__9_, s_r_21__8_, s_r_21__7_, s_r_21__6_, s_r_21__5_, s_r_21__4_, s_r_21__3_, s_r_21__2_, s_r_21__1_, s_r_21__0_ }),
    .c_o(c_r[21]),
    .prod_accum_o({ prod_accum_21__22_, prod_accum_21__21_, prod_accum_21__20_, prod_accum_21__19_, prod_accum_21__18_, prod_accum_21__17_, prod_accum_21__16_, prod_accum_21__15_, prod_accum_21__14_, prod_accum_21__13_, prod_accum_21__12_, prod_accum_21__11_, prod_accum_21__10_, prod_accum_21__9_, prod_accum_21__8_, prod_accum_21__7_, prod_accum_21__6_, prod_accum_21__5_, prod_accum_21__4_, prod_accum_21__3_, prod_accum_21__2_, prod_accum_21__1_, prod_accum_21__0_ })
  );


  bsg_mul_array_row_128_22_0
  genblk1_22__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[2815:2688]),
    .b_i(b_r[2815:2688]),
    .s_i({ s_r_21__127_, s_r_21__126_, s_r_21__125_, s_r_21__124_, s_r_21__123_, s_r_21__122_, s_r_21__121_, s_r_21__120_, s_r_21__119_, s_r_21__118_, s_r_21__117_, s_r_21__116_, s_r_21__115_, s_r_21__114_, s_r_21__113_, s_r_21__112_, s_r_21__111_, s_r_21__110_, s_r_21__109_, s_r_21__108_, s_r_21__107_, s_r_21__106_, s_r_21__105_, s_r_21__104_, s_r_21__103_, s_r_21__102_, s_r_21__101_, s_r_21__100_, s_r_21__99_, s_r_21__98_, s_r_21__97_, s_r_21__96_, s_r_21__95_, s_r_21__94_, s_r_21__93_, s_r_21__92_, s_r_21__91_, s_r_21__90_, s_r_21__89_, s_r_21__88_, s_r_21__87_, s_r_21__86_, s_r_21__85_, s_r_21__84_, s_r_21__83_, s_r_21__82_, s_r_21__81_, s_r_21__80_, s_r_21__79_, s_r_21__78_, s_r_21__77_, s_r_21__76_, s_r_21__75_, s_r_21__74_, s_r_21__73_, s_r_21__72_, s_r_21__71_, s_r_21__70_, s_r_21__69_, s_r_21__68_, s_r_21__67_, s_r_21__66_, s_r_21__65_, s_r_21__64_, s_r_21__63_, s_r_21__62_, s_r_21__61_, s_r_21__60_, s_r_21__59_, s_r_21__58_, s_r_21__57_, s_r_21__56_, s_r_21__55_, s_r_21__54_, s_r_21__53_, s_r_21__52_, s_r_21__51_, s_r_21__50_, s_r_21__49_, s_r_21__48_, s_r_21__47_, s_r_21__46_, s_r_21__45_, s_r_21__44_, s_r_21__43_, s_r_21__42_, s_r_21__41_, s_r_21__40_, s_r_21__39_, s_r_21__38_, s_r_21__37_, s_r_21__36_, s_r_21__35_, s_r_21__34_, s_r_21__33_, s_r_21__32_, s_r_21__31_, s_r_21__30_, s_r_21__29_, s_r_21__28_, s_r_21__27_, s_r_21__26_, s_r_21__25_, s_r_21__24_, s_r_21__23_, s_r_21__22_, s_r_21__21_, s_r_21__20_, s_r_21__19_, s_r_21__18_, s_r_21__17_, s_r_21__16_, s_r_21__15_, s_r_21__14_, s_r_21__13_, s_r_21__12_, s_r_21__11_, s_r_21__10_, s_r_21__9_, s_r_21__8_, s_r_21__7_, s_r_21__6_, s_r_21__5_, s_r_21__4_, s_r_21__3_, s_r_21__2_, s_r_21__1_, s_r_21__0_ }),
    .c_i(c_r[21]),
    .prod_accum_i({ prod_accum_21__22_, prod_accum_21__21_, prod_accum_21__20_, prod_accum_21__19_, prod_accum_21__18_, prod_accum_21__17_, prod_accum_21__16_, prod_accum_21__15_, prod_accum_21__14_, prod_accum_21__13_, prod_accum_21__12_, prod_accum_21__11_, prod_accum_21__10_, prod_accum_21__9_, prod_accum_21__8_, prod_accum_21__7_, prod_accum_21__6_, prod_accum_21__5_, prod_accum_21__4_, prod_accum_21__3_, prod_accum_21__2_, prod_accum_21__1_, prod_accum_21__0_ }),
    .a_o(a_r[2943:2816]),
    .b_o(b_r[2943:2816]),
    .s_o({ s_r_22__127_, s_r_22__126_, s_r_22__125_, s_r_22__124_, s_r_22__123_, s_r_22__122_, s_r_22__121_, s_r_22__120_, s_r_22__119_, s_r_22__118_, s_r_22__117_, s_r_22__116_, s_r_22__115_, s_r_22__114_, s_r_22__113_, s_r_22__112_, s_r_22__111_, s_r_22__110_, s_r_22__109_, s_r_22__108_, s_r_22__107_, s_r_22__106_, s_r_22__105_, s_r_22__104_, s_r_22__103_, s_r_22__102_, s_r_22__101_, s_r_22__100_, s_r_22__99_, s_r_22__98_, s_r_22__97_, s_r_22__96_, s_r_22__95_, s_r_22__94_, s_r_22__93_, s_r_22__92_, s_r_22__91_, s_r_22__90_, s_r_22__89_, s_r_22__88_, s_r_22__87_, s_r_22__86_, s_r_22__85_, s_r_22__84_, s_r_22__83_, s_r_22__82_, s_r_22__81_, s_r_22__80_, s_r_22__79_, s_r_22__78_, s_r_22__77_, s_r_22__76_, s_r_22__75_, s_r_22__74_, s_r_22__73_, s_r_22__72_, s_r_22__71_, s_r_22__70_, s_r_22__69_, s_r_22__68_, s_r_22__67_, s_r_22__66_, s_r_22__65_, s_r_22__64_, s_r_22__63_, s_r_22__62_, s_r_22__61_, s_r_22__60_, s_r_22__59_, s_r_22__58_, s_r_22__57_, s_r_22__56_, s_r_22__55_, s_r_22__54_, s_r_22__53_, s_r_22__52_, s_r_22__51_, s_r_22__50_, s_r_22__49_, s_r_22__48_, s_r_22__47_, s_r_22__46_, s_r_22__45_, s_r_22__44_, s_r_22__43_, s_r_22__42_, s_r_22__41_, s_r_22__40_, s_r_22__39_, s_r_22__38_, s_r_22__37_, s_r_22__36_, s_r_22__35_, s_r_22__34_, s_r_22__33_, s_r_22__32_, s_r_22__31_, s_r_22__30_, s_r_22__29_, s_r_22__28_, s_r_22__27_, s_r_22__26_, s_r_22__25_, s_r_22__24_, s_r_22__23_, s_r_22__22_, s_r_22__21_, s_r_22__20_, s_r_22__19_, s_r_22__18_, s_r_22__17_, s_r_22__16_, s_r_22__15_, s_r_22__14_, s_r_22__13_, s_r_22__12_, s_r_22__11_, s_r_22__10_, s_r_22__9_, s_r_22__8_, s_r_22__7_, s_r_22__6_, s_r_22__5_, s_r_22__4_, s_r_22__3_, s_r_22__2_, s_r_22__1_, s_r_22__0_ }),
    .c_o(c_r[22]),
    .prod_accum_o({ prod_accum_22__23_, prod_accum_22__22_, prod_accum_22__21_, prod_accum_22__20_, prod_accum_22__19_, prod_accum_22__18_, prod_accum_22__17_, prod_accum_22__16_, prod_accum_22__15_, prod_accum_22__14_, prod_accum_22__13_, prod_accum_22__12_, prod_accum_22__11_, prod_accum_22__10_, prod_accum_22__9_, prod_accum_22__8_, prod_accum_22__7_, prod_accum_22__6_, prod_accum_22__5_, prod_accum_22__4_, prod_accum_22__3_, prod_accum_22__2_, prod_accum_22__1_, prod_accum_22__0_ })
  );


  bsg_mul_array_row_128_23_0
  genblk1_23__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[2943:2816]),
    .b_i(b_r[2943:2816]),
    .s_i({ s_r_22__127_, s_r_22__126_, s_r_22__125_, s_r_22__124_, s_r_22__123_, s_r_22__122_, s_r_22__121_, s_r_22__120_, s_r_22__119_, s_r_22__118_, s_r_22__117_, s_r_22__116_, s_r_22__115_, s_r_22__114_, s_r_22__113_, s_r_22__112_, s_r_22__111_, s_r_22__110_, s_r_22__109_, s_r_22__108_, s_r_22__107_, s_r_22__106_, s_r_22__105_, s_r_22__104_, s_r_22__103_, s_r_22__102_, s_r_22__101_, s_r_22__100_, s_r_22__99_, s_r_22__98_, s_r_22__97_, s_r_22__96_, s_r_22__95_, s_r_22__94_, s_r_22__93_, s_r_22__92_, s_r_22__91_, s_r_22__90_, s_r_22__89_, s_r_22__88_, s_r_22__87_, s_r_22__86_, s_r_22__85_, s_r_22__84_, s_r_22__83_, s_r_22__82_, s_r_22__81_, s_r_22__80_, s_r_22__79_, s_r_22__78_, s_r_22__77_, s_r_22__76_, s_r_22__75_, s_r_22__74_, s_r_22__73_, s_r_22__72_, s_r_22__71_, s_r_22__70_, s_r_22__69_, s_r_22__68_, s_r_22__67_, s_r_22__66_, s_r_22__65_, s_r_22__64_, s_r_22__63_, s_r_22__62_, s_r_22__61_, s_r_22__60_, s_r_22__59_, s_r_22__58_, s_r_22__57_, s_r_22__56_, s_r_22__55_, s_r_22__54_, s_r_22__53_, s_r_22__52_, s_r_22__51_, s_r_22__50_, s_r_22__49_, s_r_22__48_, s_r_22__47_, s_r_22__46_, s_r_22__45_, s_r_22__44_, s_r_22__43_, s_r_22__42_, s_r_22__41_, s_r_22__40_, s_r_22__39_, s_r_22__38_, s_r_22__37_, s_r_22__36_, s_r_22__35_, s_r_22__34_, s_r_22__33_, s_r_22__32_, s_r_22__31_, s_r_22__30_, s_r_22__29_, s_r_22__28_, s_r_22__27_, s_r_22__26_, s_r_22__25_, s_r_22__24_, s_r_22__23_, s_r_22__22_, s_r_22__21_, s_r_22__20_, s_r_22__19_, s_r_22__18_, s_r_22__17_, s_r_22__16_, s_r_22__15_, s_r_22__14_, s_r_22__13_, s_r_22__12_, s_r_22__11_, s_r_22__10_, s_r_22__9_, s_r_22__8_, s_r_22__7_, s_r_22__6_, s_r_22__5_, s_r_22__4_, s_r_22__3_, s_r_22__2_, s_r_22__1_, s_r_22__0_ }),
    .c_i(c_r[22]),
    .prod_accum_i({ prod_accum_22__23_, prod_accum_22__22_, prod_accum_22__21_, prod_accum_22__20_, prod_accum_22__19_, prod_accum_22__18_, prod_accum_22__17_, prod_accum_22__16_, prod_accum_22__15_, prod_accum_22__14_, prod_accum_22__13_, prod_accum_22__12_, prod_accum_22__11_, prod_accum_22__10_, prod_accum_22__9_, prod_accum_22__8_, prod_accum_22__7_, prod_accum_22__6_, prod_accum_22__5_, prod_accum_22__4_, prod_accum_22__3_, prod_accum_22__2_, prod_accum_22__1_, prod_accum_22__0_ }),
    .a_o(a_r[3071:2944]),
    .b_o(b_r[3071:2944]),
    .s_o({ s_r_23__127_, s_r_23__126_, s_r_23__125_, s_r_23__124_, s_r_23__123_, s_r_23__122_, s_r_23__121_, s_r_23__120_, s_r_23__119_, s_r_23__118_, s_r_23__117_, s_r_23__116_, s_r_23__115_, s_r_23__114_, s_r_23__113_, s_r_23__112_, s_r_23__111_, s_r_23__110_, s_r_23__109_, s_r_23__108_, s_r_23__107_, s_r_23__106_, s_r_23__105_, s_r_23__104_, s_r_23__103_, s_r_23__102_, s_r_23__101_, s_r_23__100_, s_r_23__99_, s_r_23__98_, s_r_23__97_, s_r_23__96_, s_r_23__95_, s_r_23__94_, s_r_23__93_, s_r_23__92_, s_r_23__91_, s_r_23__90_, s_r_23__89_, s_r_23__88_, s_r_23__87_, s_r_23__86_, s_r_23__85_, s_r_23__84_, s_r_23__83_, s_r_23__82_, s_r_23__81_, s_r_23__80_, s_r_23__79_, s_r_23__78_, s_r_23__77_, s_r_23__76_, s_r_23__75_, s_r_23__74_, s_r_23__73_, s_r_23__72_, s_r_23__71_, s_r_23__70_, s_r_23__69_, s_r_23__68_, s_r_23__67_, s_r_23__66_, s_r_23__65_, s_r_23__64_, s_r_23__63_, s_r_23__62_, s_r_23__61_, s_r_23__60_, s_r_23__59_, s_r_23__58_, s_r_23__57_, s_r_23__56_, s_r_23__55_, s_r_23__54_, s_r_23__53_, s_r_23__52_, s_r_23__51_, s_r_23__50_, s_r_23__49_, s_r_23__48_, s_r_23__47_, s_r_23__46_, s_r_23__45_, s_r_23__44_, s_r_23__43_, s_r_23__42_, s_r_23__41_, s_r_23__40_, s_r_23__39_, s_r_23__38_, s_r_23__37_, s_r_23__36_, s_r_23__35_, s_r_23__34_, s_r_23__33_, s_r_23__32_, s_r_23__31_, s_r_23__30_, s_r_23__29_, s_r_23__28_, s_r_23__27_, s_r_23__26_, s_r_23__25_, s_r_23__24_, s_r_23__23_, s_r_23__22_, s_r_23__21_, s_r_23__20_, s_r_23__19_, s_r_23__18_, s_r_23__17_, s_r_23__16_, s_r_23__15_, s_r_23__14_, s_r_23__13_, s_r_23__12_, s_r_23__11_, s_r_23__10_, s_r_23__9_, s_r_23__8_, s_r_23__7_, s_r_23__6_, s_r_23__5_, s_r_23__4_, s_r_23__3_, s_r_23__2_, s_r_23__1_, s_r_23__0_ }),
    .c_o(c_r[23]),
    .prod_accum_o({ prod_accum_23__24_, prod_accum_23__23_, prod_accum_23__22_, prod_accum_23__21_, prod_accum_23__20_, prod_accum_23__19_, prod_accum_23__18_, prod_accum_23__17_, prod_accum_23__16_, prod_accum_23__15_, prod_accum_23__14_, prod_accum_23__13_, prod_accum_23__12_, prod_accum_23__11_, prod_accum_23__10_, prod_accum_23__9_, prod_accum_23__8_, prod_accum_23__7_, prod_accum_23__6_, prod_accum_23__5_, prod_accum_23__4_, prod_accum_23__3_, prod_accum_23__2_, prod_accum_23__1_, prod_accum_23__0_ })
  );


  bsg_mul_array_row_128_24_0
  genblk1_24__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[3071:2944]),
    .b_i(b_r[3071:2944]),
    .s_i({ s_r_23__127_, s_r_23__126_, s_r_23__125_, s_r_23__124_, s_r_23__123_, s_r_23__122_, s_r_23__121_, s_r_23__120_, s_r_23__119_, s_r_23__118_, s_r_23__117_, s_r_23__116_, s_r_23__115_, s_r_23__114_, s_r_23__113_, s_r_23__112_, s_r_23__111_, s_r_23__110_, s_r_23__109_, s_r_23__108_, s_r_23__107_, s_r_23__106_, s_r_23__105_, s_r_23__104_, s_r_23__103_, s_r_23__102_, s_r_23__101_, s_r_23__100_, s_r_23__99_, s_r_23__98_, s_r_23__97_, s_r_23__96_, s_r_23__95_, s_r_23__94_, s_r_23__93_, s_r_23__92_, s_r_23__91_, s_r_23__90_, s_r_23__89_, s_r_23__88_, s_r_23__87_, s_r_23__86_, s_r_23__85_, s_r_23__84_, s_r_23__83_, s_r_23__82_, s_r_23__81_, s_r_23__80_, s_r_23__79_, s_r_23__78_, s_r_23__77_, s_r_23__76_, s_r_23__75_, s_r_23__74_, s_r_23__73_, s_r_23__72_, s_r_23__71_, s_r_23__70_, s_r_23__69_, s_r_23__68_, s_r_23__67_, s_r_23__66_, s_r_23__65_, s_r_23__64_, s_r_23__63_, s_r_23__62_, s_r_23__61_, s_r_23__60_, s_r_23__59_, s_r_23__58_, s_r_23__57_, s_r_23__56_, s_r_23__55_, s_r_23__54_, s_r_23__53_, s_r_23__52_, s_r_23__51_, s_r_23__50_, s_r_23__49_, s_r_23__48_, s_r_23__47_, s_r_23__46_, s_r_23__45_, s_r_23__44_, s_r_23__43_, s_r_23__42_, s_r_23__41_, s_r_23__40_, s_r_23__39_, s_r_23__38_, s_r_23__37_, s_r_23__36_, s_r_23__35_, s_r_23__34_, s_r_23__33_, s_r_23__32_, s_r_23__31_, s_r_23__30_, s_r_23__29_, s_r_23__28_, s_r_23__27_, s_r_23__26_, s_r_23__25_, s_r_23__24_, s_r_23__23_, s_r_23__22_, s_r_23__21_, s_r_23__20_, s_r_23__19_, s_r_23__18_, s_r_23__17_, s_r_23__16_, s_r_23__15_, s_r_23__14_, s_r_23__13_, s_r_23__12_, s_r_23__11_, s_r_23__10_, s_r_23__9_, s_r_23__8_, s_r_23__7_, s_r_23__6_, s_r_23__5_, s_r_23__4_, s_r_23__3_, s_r_23__2_, s_r_23__1_, s_r_23__0_ }),
    .c_i(c_r[23]),
    .prod_accum_i({ prod_accum_23__24_, prod_accum_23__23_, prod_accum_23__22_, prod_accum_23__21_, prod_accum_23__20_, prod_accum_23__19_, prod_accum_23__18_, prod_accum_23__17_, prod_accum_23__16_, prod_accum_23__15_, prod_accum_23__14_, prod_accum_23__13_, prod_accum_23__12_, prod_accum_23__11_, prod_accum_23__10_, prod_accum_23__9_, prod_accum_23__8_, prod_accum_23__7_, prod_accum_23__6_, prod_accum_23__5_, prod_accum_23__4_, prod_accum_23__3_, prod_accum_23__2_, prod_accum_23__1_, prod_accum_23__0_ }),
    .a_o(a_r[3199:3072]),
    .b_o(b_r[3199:3072]),
    .s_o({ s_r_24__127_, s_r_24__126_, s_r_24__125_, s_r_24__124_, s_r_24__123_, s_r_24__122_, s_r_24__121_, s_r_24__120_, s_r_24__119_, s_r_24__118_, s_r_24__117_, s_r_24__116_, s_r_24__115_, s_r_24__114_, s_r_24__113_, s_r_24__112_, s_r_24__111_, s_r_24__110_, s_r_24__109_, s_r_24__108_, s_r_24__107_, s_r_24__106_, s_r_24__105_, s_r_24__104_, s_r_24__103_, s_r_24__102_, s_r_24__101_, s_r_24__100_, s_r_24__99_, s_r_24__98_, s_r_24__97_, s_r_24__96_, s_r_24__95_, s_r_24__94_, s_r_24__93_, s_r_24__92_, s_r_24__91_, s_r_24__90_, s_r_24__89_, s_r_24__88_, s_r_24__87_, s_r_24__86_, s_r_24__85_, s_r_24__84_, s_r_24__83_, s_r_24__82_, s_r_24__81_, s_r_24__80_, s_r_24__79_, s_r_24__78_, s_r_24__77_, s_r_24__76_, s_r_24__75_, s_r_24__74_, s_r_24__73_, s_r_24__72_, s_r_24__71_, s_r_24__70_, s_r_24__69_, s_r_24__68_, s_r_24__67_, s_r_24__66_, s_r_24__65_, s_r_24__64_, s_r_24__63_, s_r_24__62_, s_r_24__61_, s_r_24__60_, s_r_24__59_, s_r_24__58_, s_r_24__57_, s_r_24__56_, s_r_24__55_, s_r_24__54_, s_r_24__53_, s_r_24__52_, s_r_24__51_, s_r_24__50_, s_r_24__49_, s_r_24__48_, s_r_24__47_, s_r_24__46_, s_r_24__45_, s_r_24__44_, s_r_24__43_, s_r_24__42_, s_r_24__41_, s_r_24__40_, s_r_24__39_, s_r_24__38_, s_r_24__37_, s_r_24__36_, s_r_24__35_, s_r_24__34_, s_r_24__33_, s_r_24__32_, s_r_24__31_, s_r_24__30_, s_r_24__29_, s_r_24__28_, s_r_24__27_, s_r_24__26_, s_r_24__25_, s_r_24__24_, s_r_24__23_, s_r_24__22_, s_r_24__21_, s_r_24__20_, s_r_24__19_, s_r_24__18_, s_r_24__17_, s_r_24__16_, s_r_24__15_, s_r_24__14_, s_r_24__13_, s_r_24__12_, s_r_24__11_, s_r_24__10_, s_r_24__9_, s_r_24__8_, s_r_24__7_, s_r_24__6_, s_r_24__5_, s_r_24__4_, s_r_24__3_, s_r_24__2_, s_r_24__1_, s_r_24__0_ }),
    .c_o(c_r[24]),
    .prod_accum_o({ prod_accum_24__25_, prod_accum_24__24_, prod_accum_24__23_, prod_accum_24__22_, prod_accum_24__21_, prod_accum_24__20_, prod_accum_24__19_, prod_accum_24__18_, prod_accum_24__17_, prod_accum_24__16_, prod_accum_24__15_, prod_accum_24__14_, prod_accum_24__13_, prod_accum_24__12_, prod_accum_24__11_, prod_accum_24__10_, prod_accum_24__9_, prod_accum_24__8_, prod_accum_24__7_, prod_accum_24__6_, prod_accum_24__5_, prod_accum_24__4_, prod_accum_24__3_, prod_accum_24__2_, prod_accum_24__1_, prod_accum_24__0_ })
  );


  bsg_mul_array_row_128_25_0
  genblk1_25__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[3199:3072]),
    .b_i(b_r[3199:3072]),
    .s_i({ s_r_24__127_, s_r_24__126_, s_r_24__125_, s_r_24__124_, s_r_24__123_, s_r_24__122_, s_r_24__121_, s_r_24__120_, s_r_24__119_, s_r_24__118_, s_r_24__117_, s_r_24__116_, s_r_24__115_, s_r_24__114_, s_r_24__113_, s_r_24__112_, s_r_24__111_, s_r_24__110_, s_r_24__109_, s_r_24__108_, s_r_24__107_, s_r_24__106_, s_r_24__105_, s_r_24__104_, s_r_24__103_, s_r_24__102_, s_r_24__101_, s_r_24__100_, s_r_24__99_, s_r_24__98_, s_r_24__97_, s_r_24__96_, s_r_24__95_, s_r_24__94_, s_r_24__93_, s_r_24__92_, s_r_24__91_, s_r_24__90_, s_r_24__89_, s_r_24__88_, s_r_24__87_, s_r_24__86_, s_r_24__85_, s_r_24__84_, s_r_24__83_, s_r_24__82_, s_r_24__81_, s_r_24__80_, s_r_24__79_, s_r_24__78_, s_r_24__77_, s_r_24__76_, s_r_24__75_, s_r_24__74_, s_r_24__73_, s_r_24__72_, s_r_24__71_, s_r_24__70_, s_r_24__69_, s_r_24__68_, s_r_24__67_, s_r_24__66_, s_r_24__65_, s_r_24__64_, s_r_24__63_, s_r_24__62_, s_r_24__61_, s_r_24__60_, s_r_24__59_, s_r_24__58_, s_r_24__57_, s_r_24__56_, s_r_24__55_, s_r_24__54_, s_r_24__53_, s_r_24__52_, s_r_24__51_, s_r_24__50_, s_r_24__49_, s_r_24__48_, s_r_24__47_, s_r_24__46_, s_r_24__45_, s_r_24__44_, s_r_24__43_, s_r_24__42_, s_r_24__41_, s_r_24__40_, s_r_24__39_, s_r_24__38_, s_r_24__37_, s_r_24__36_, s_r_24__35_, s_r_24__34_, s_r_24__33_, s_r_24__32_, s_r_24__31_, s_r_24__30_, s_r_24__29_, s_r_24__28_, s_r_24__27_, s_r_24__26_, s_r_24__25_, s_r_24__24_, s_r_24__23_, s_r_24__22_, s_r_24__21_, s_r_24__20_, s_r_24__19_, s_r_24__18_, s_r_24__17_, s_r_24__16_, s_r_24__15_, s_r_24__14_, s_r_24__13_, s_r_24__12_, s_r_24__11_, s_r_24__10_, s_r_24__9_, s_r_24__8_, s_r_24__7_, s_r_24__6_, s_r_24__5_, s_r_24__4_, s_r_24__3_, s_r_24__2_, s_r_24__1_, s_r_24__0_ }),
    .c_i(c_r[24]),
    .prod_accum_i({ prod_accum_24__25_, prod_accum_24__24_, prod_accum_24__23_, prod_accum_24__22_, prod_accum_24__21_, prod_accum_24__20_, prod_accum_24__19_, prod_accum_24__18_, prod_accum_24__17_, prod_accum_24__16_, prod_accum_24__15_, prod_accum_24__14_, prod_accum_24__13_, prod_accum_24__12_, prod_accum_24__11_, prod_accum_24__10_, prod_accum_24__9_, prod_accum_24__8_, prod_accum_24__7_, prod_accum_24__6_, prod_accum_24__5_, prod_accum_24__4_, prod_accum_24__3_, prod_accum_24__2_, prod_accum_24__1_, prod_accum_24__0_ }),
    .a_o(a_r[3327:3200]),
    .b_o(b_r[3327:3200]),
    .s_o({ s_r_25__127_, s_r_25__126_, s_r_25__125_, s_r_25__124_, s_r_25__123_, s_r_25__122_, s_r_25__121_, s_r_25__120_, s_r_25__119_, s_r_25__118_, s_r_25__117_, s_r_25__116_, s_r_25__115_, s_r_25__114_, s_r_25__113_, s_r_25__112_, s_r_25__111_, s_r_25__110_, s_r_25__109_, s_r_25__108_, s_r_25__107_, s_r_25__106_, s_r_25__105_, s_r_25__104_, s_r_25__103_, s_r_25__102_, s_r_25__101_, s_r_25__100_, s_r_25__99_, s_r_25__98_, s_r_25__97_, s_r_25__96_, s_r_25__95_, s_r_25__94_, s_r_25__93_, s_r_25__92_, s_r_25__91_, s_r_25__90_, s_r_25__89_, s_r_25__88_, s_r_25__87_, s_r_25__86_, s_r_25__85_, s_r_25__84_, s_r_25__83_, s_r_25__82_, s_r_25__81_, s_r_25__80_, s_r_25__79_, s_r_25__78_, s_r_25__77_, s_r_25__76_, s_r_25__75_, s_r_25__74_, s_r_25__73_, s_r_25__72_, s_r_25__71_, s_r_25__70_, s_r_25__69_, s_r_25__68_, s_r_25__67_, s_r_25__66_, s_r_25__65_, s_r_25__64_, s_r_25__63_, s_r_25__62_, s_r_25__61_, s_r_25__60_, s_r_25__59_, s_r_25__58_, s_r_25__57_, s_r_25__56_, s_r_25__55_, s_r_25__54_, s_r_25__53_, s_r_25__52_, s_r_25__51_, s_r_25__50_, s_r_25__49_, s_r_25__48_, s_r_25__47_, s_r_25__46_, s_r_25__45_, s_r_25__44_, s_r_25__43_, s_r_25__42_, s_r_25__41_, s_r_25__40_, s_r_25__39_, s_r_25__38_, s_r_25__37_, s_r_25__36_, s_r_25__35_, s_r_25__34_, s_r_25__33_, s_r_25__32_, s_r_25__31_, s_r_25__30_, s_r_25__29_, s_r_25__28_, s_r_25__27_, s_r_25__26_, s_r_25__25_, s_r_25__24_, s_r_25__23_, s_r_25__22_, s_r_25__21_, s_r_25__20_, s_r_25__19_, s_r_25__18_, s_r_25__17_, s_r_25__16_, s_r_25__15_, s_r_25__14_, s_r_25__13_, s_r_25__12_, s_r_25__11_, s_r_25__10_, s_r_25__9_, s_r_25__8_, s_r_25__7_, s_r_25__6_, s_r_25__5_, s_r_25__4_, s_r_25__3_, s_r_25__2_, s_r_25__1_, s_r_25__0_ }),
    .c_o(c_r[25]),
    .prod_accum_o({ prod_accum_25__26_, prod_accum_25__25_, prod_accum_25__24_, prod_accum_25__23_, prod_accum_25__22_, prod_accum_25__21_, prod_accum_25__20_, prod_accum_25__19_, prod_accum_25__18_, prod_accum_25__17_, prod_accum_25__16_, prod_accum_25__15_, prod_accum_25__14_, prod_accum_25__13_, prod_accum_25__12_, prod_accum_25__11_, prod_accum_25__10_, prod_accum_25__9_, prod_accum_25__8_, prod_accum_25__7_, prod_accum_25__6_, prod_accum_25__5_, prod_accum_25__4_, prod_accum_25__3_, prod_accum_25__2_, prod_accum_25__1_, prod_accum_25__0_ })
  );


  bsg_mul_array_row_128_26_0
  genblk1_26__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[3327:3200]),
    .b_i(b_r[3327:3200]),
    .s_i({ s_r_25__127_, s_r_25__126_, s_r_25__125_, s_r_25__124_, s_r_25__123_, s_r_25__122_, s_r_25__121_, s_r_25__120_, s_r_25__119_, s_r_25__118_, s_r_25__117_, s_r_25__116_, s_r_25__115_, s_r_25__114_, s_r_25__113_, s_r_25__112_, s_r_25__111_, s_r_25__110_, s_r_25__109_, s_r_25__108_, s_r_25__107_, s_r_25__106_, s_r_25__105_, s_r_25__104_, s_r_25__103_, s_r_25__102_, s_r_25__101_, s_r_25__100_, s_r_25__99_, s_r_25__98_, s_r_25__97_, s_r_25__96_, s_r_25__95_, s_r_25__94_, s_r_25__93_, s_r_25__92_, s_r_25__91_, s_r_25__90_, s_r_25__89_, s_r_25__88_, s_r_25__87_, s_r_25__86_, s_r_25__85_, s_r_25__84_, s_r_25__83_, s_r_25__82_, s_r_25__81_, s_r_25__80_, s_r_25__79_, s_r_25__78_, s_r_25__77_, s_r_25__76_, s_r_25__75_, s_r_25__74_, s_r_25__73_, s_r_25__72_, s_r_25__71_, s_r_25__70_, s_r_25__69_, s_r_25__68_, s_r_25__67_, s_r_25__66_, s_r_25__65_, s_r_25__64_, s_r_25__63_, s_r_25__62_, s_r_25__61_, s_r_25__60_, s_r_25__59_, s_r_25__58_, s_r_25__57_, s_r_25__56_, s_r_25__55_, s_r_25__54_, s_r_25__53_, s_r_25__52_, s_r_25__51_, s_r_25__50_, s_r_25__49_, s_r_25__48_, s_r_25__47_, s_r_25__46_, s_r_25__45_, s_r_25__44_, s_r_25__43_, s_r_25__42_, s_r_25__41_, s_r_25__40_, s_r_25__39_, s_r_25__38_, s_r_25__37_, s_r_25__36_, s_r_25__35_, s_r_25__34_, s_r_25__33_, s_r_25__32_, s_r_25__31_, s_r_25__30_, s_r_25__29_, s_r_25__28_, s_r_25__27_, s_r_25__26_, s_r_25__25_, s_r_25__24_, s_r_25__23_, s_r_25__22_, s_r_25__21_, s_r_25__20_, s_r_25__19_, s_r_25__18_, s_r_25__17_, s_r_25__16_, s_r_25__15_, s_r_25__14_, s_r_25__13_, s_r_25__12_, s_r_25__11_, s_r_25__10_, s_r_25__9_, s_r_25__8_, s_r_25__7_, s_r_25__6_, s_r_25__5_, s_r_25__4_, s_r_25__3_, s_r_25__2_, s_r_25__1_, s_r_25__0_ }),
    .c_i(c_r[25]),
    .prod_accum_i({ prod_accum_25__26_, prod_accum_25__25_, prod_accum_25__24_, prod_accum_25__23_, prod_accum_25__22_, prod_accum_25__21_, prod_accum_25__20_, prod_accum_25__19_, prod_accum_25__18_, prod_accum_25__17_, prod_accum_25__16_, prod_accum_25__15_, prod_accum_25__14_, prod_accum_25__13_, prod_accum_25__12_, prod_accum_25__11_, prod_accum_25__10_, prod_accum_25__9_, prod_accum_25__8_, prod_accum_25__7_, prod_accum_25__6_, prod_accum_25__5_, prod_accum_25__4_, prod_accum_25__3_, prod_accum_25__2_, prod_accum_25__1_, prod_accum_25__0_ }),
    .a_o(a_r[3455:3328]),
    .b_o(b_r[3455:3328]),
    .s_o({ s_r_26__127_, s_r_26__126_, s_r_26__125_, s_r_26__124_, s_r_26__123_, s_r_26__122_, s_r_26__121_, s_r_26__120_, s_r_26__119_, s_r_26__118_, s_r_26__117_, s_r_26__116_, s_r_26__115_, s_r_26__114_, s_r_26__113_, s_r_26__112_, s_r_26__111_, s_r_26__110_, s_r_26__109_, s_r_26__108_, s_r_26__107_, s_r_26__106_, s_r_26__105_, s_r_26__104_, s_r_26__103_, s_r_26__102_, s_r_26__101_, s_r_26__100_, s_r_26__99_, s_r_26__98_, s_r_26__97_, s_r_26__96_, s_r_26__95_, s_r_26__94_, s_r_26__93_, s_r_26__92_, s_r_26__91_, s_r_26__90_, s_r_26__89_, s_r_26__88_, s_r_26__87_, s_r_26__86_, s_r_26__85_, s_r_26__84_, s_r_26__83_, s_r_26__82_, s_r_26__81_, s_r_26__80_, s_r_26__79_, s_r_26__78_, s_r_26__77_, s_r_26__76_, s_r_26__75_, s_r_26__74_, s_r_26__73_, s_r_26__72_, s_r_26__71_, s_r_26__70_, s_r_26__69_, s_r_26__68_, s_r_26__67_, s_r_26__66_, s_r_26__65_, s_r_26__64_, s_r_26__63_, s_r_26__62_, s_r_26__61_, s_r_26__60_, s_r_26__59_, s_r_26__58_, s_r_26__57_, s_r_26__56_, s_r_26__55_, s_r_26__54_, s_r_26__53_, s_r_26__52_, s_r_26__51_, s_r_26__50_, s_r_26__49_, s_r_26__48_, s_r_26__47_, s_r_26__46_, s_r_26__45_, s_r_26__44_, s_r_26__43_, s_r_26__42_, s_r_26__41_, s_r_26__40_, s_r_26__39_, s_r_26__38_, s_r_26__37_, s_r_26__36_, s_r_26__35_, s_r_26__34_, s_r_26__33_, s_r_26__32_, s_r_26__31_, s_r_26__30_, s_r_26__29_, s_r_26__28_, s_r_26__27_, s_r_26__26_, s_r_26__25_, s_r_26__24_, s_r_26__23_, s_r_26__22_, s_r_26__21_, s_r_26__20_, s_r_26__19_, s_r_26__18_, s_r_26__17_, s_r_26__16_, s_r_26__15_, s_r_26__14_, s_r_26__13_, s_r_26__12_, s_r_26__11_, s_r_26__10_, s_r_26__9_, s_r_26__8_, s_r_26__7_, s_r_26__6_, s_r_26__5_, s_r_26__4_, s_r_26__3_, s_r_26__2_, s_r_26__1_, s_r_26__0_ }),
    .c_o(c_r[26]),
    .prod_accum_o({ prod_accum_26__27_, prod_accum_26__26_, prod_accum_26__25_, prod_accum_26__24_, prod_accum_26__23_, prod_accum_26__22_, prod_accum_26__21_, prod_accum_26__20_, prod_accum_26__19_, prod_accum_26__18_, prod_accum_26__17_, prod_accum_26__16_, prod_accum_26__15_, prod_accum_26__14_, prod_accum_26__13_, prod_accum_26__12_, prod_accum_26__11_, prod_accum_26__10_, prod_accum_26__9_, prod_accum_26__8_, prod_accum_26__7_, prod_accum_26__6_, prod_accum_26__5_, prod_accum_26__4_, prod_accum_26__3_, prod_accum_26__2_, prod_accum_26__1_, prod_accum_26__0_ })
  );


  bsg_mul_array_row_128_27_0
  genblk1_27__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[3455:3328]),
    .b_i(b_r[3455:3328]),
    .s_i({ s_r_26__127_, s_r_26__126_, s_r_26__125_, s_r_26__124_, s_r_26__123_, s_r_26__122_, s_r_26__121_, s_r_26__120_, s_r_26__119_, s_r_26__118_, s_r_26__117_, s_r_26__116_, s_r_26__115_, s_r_26__114_, s_r_26__113_, s_r_26__112_, s_r_26__111_, s_r_26__110_, s_r_26__109_, s_r_26__108_, s_r_26__107_, s_r_26__106_, s_r_26__105_, s_r_26__104_, s_r_26__103_, s_r_26__102_, s_r_26__101_, s_r_26__100_, s_r_26__99_, s_r_26__98_, s_r_26__97_, s_r_26__96_, s_r_26__95_, s_r_26__94_, s_r_26__93_, s_r_26__92_, s_r_26__91_, s_r_26__90_, s_r_26__89_, s_r_26__88_, s_r_26__87_, s_r_26__86_, s_r_26__85_, s_r_26__84_, s_r_26__83_, s_r_26__82_, s_r_26__81_, s_r_26__80_, s_r_26__79_, s_r_26__78_, s_r_26__77_, s_r_26__76_, s_r_26__75_, s_r_26__74_, s_r_26__73_, s_r_26__72_, s_r_26__71_, s_r_26__70_, s_r_26__69_, s_r_26__68_, s_r_26__67_, s_r_26__66_, s_r_26__65_, s_r_26__64_, s_r_26__63_, s_r_26__62_, s_r_26__61_, s_r_26__60_, s_r_26__59_, s_r_26__58_, s_r_26__57_, s_r_26__56_, s_r_26__55_, s_r_26__54_, s_r_26__53_, s_r_26__52_, s_r_26__51_, s_r_26__50_, s_r_26__49_, s_r_26__48_, s_r_26__47_, s_r_26__46_, s_r_26__45_, s_r_26__44_, s_r_26__43_, s_r_26__42_, s_r_26__41_, s_r_26__40_, s_r_26__39_, s_r_26__38_, s_r_26__37_, s_r_26__36_, s_r_26__35_, s_r_26__34_, s_r_26__33_, s_r_26__32_, s_r_26__31_, s_r_26__30_, s_r_26__29_, s_r_26__28_, s_r_26__27_, s_r_26__26_, s_r_26__25_, s_r_26__24_, s_r_26__23_, s_r_26__22_, s_r_26__21_, s_r_26__20_, s_r_26__19_, s_r_26__18_, s_r_26__17_, s_r_26__16_, s_r_26__15_, s_r_26__14_, s_r_26__13_, s_r_26__12_, s_r_26__11_, s_r_26__10_, s_r_26__9_, s_r_26__8_, s_r_26__7_, s_r_26__6_, s_r_26__5_, s_r_26__4_, s_r_26__3_, s_r_26__2_, s_r_26__1_, s_r_26__0_ }),
    .c_i(c_r[26]),
    .prod_accum_i({ prod_accum_26__27_, prod_accum_26__26_, prod_accum_26__25_, prod_accum_26__24_, prod_accum_26__23_, prod_accum_26__22_, prod_accum_26__21_, prod_accum_26__20_, prod_accum_26__19_, prod_accum_26__18_, prod_accum_26__17_, prod_accum_26__16_, prod_accum_26__15_, prod_accum_26__14_, prod_accum_26__13_, prod_accum_26__12_, prod_accum_26__11_, prod_accum_26__10_, prod_accum_26__9_, prod_accum_26__8_, prod_accum_26__7_, prod_accum_26__6_, prod_accum_26__5_, prod_accum_26__4_, prod_accum_26__3_, prod_accum_26__2_, prod_accum_26__1_, prod_accum_26__0_ }),
    .a_o(a_r[3583:3456]),
    .b_o(b_r[3583:3456]),
    .s_o({ s_r_27__127_, s_r_27__126_, s_r_27__125_, s_r_27__124_, s_r_27__123_, s_r_27__122_, s_r_27__121_, s_r_27__120_, s_r_27__119_, s_r_27__118_, s_r_27__117_, s_r_27__116_, s_r_27__115_, s_r_27__114_, s_r_27__113_, s_r_27__112_, s_r_27__111_, s_r_27__110_, s_r_27__109_, s_r_27__108_, s_r_27__107_, s_r_27__106_, s_r_27__105_, s_r_27__104_, s_r_27__103_, s_r_27__102_, s_r_27__101_, s_r_27__100_, s_r_27__99_, s_r_27__98_, s_r_27__97_, s_r_27__96_, s_r_27__95_, s_r_27__94_, s_r_27__93_, s_r_27__92_, s_r_27__91_, s_r_27__90_, s_r_27__89_, s_r_27__88_, s_r_27__87_, s_r_27__86_, s_r_27__85_, s_r_27__84_, s_r_27__83_, s_r_27__82_, s_r_27__81_, s_r_27__80_, s_r_27__79_, s_r_27__78_, s_r_27__77_, s_r_27__76_, s_r_27__75_, s_r_27__74_, s_r_27__73_, s_r_27__72_, s_r_27__71_, s_r_27__70_, s_r_27__69_, s_r_27__68_, s_r_27__67_, s_r_27__66_, s_r_27__65_, s_r_27__64_, s_r_27__63_, s_r_27__62_, s_r_27__61_, s_r_27__60_, s_r_27__59_, s_r_27__58_, s_r_27__57_, s_r_27__56_, s_r_27__55_, s_r_27__54_, s_r_27__53_, s_r_27__52_, s_r_27__51_, s_r_27__50_, s_r_27__49_, s_r_27__48_, s_r_27__47_, s_r_27__46_, s_r_27__45_, s_r_27__44_, s_r_27__43_, s_r_27__42_, s_r_27__41_, s_r_27__40_, s_r_27__39_, s_r_27__38_, s_r_27__37_, s_r_27__36_, s_r_27__35_, s_r_27__34_, s_r_27__33_, s_r_27__32_, s_r_27__31_, s_r_27__30_, s_r_27__29_, s_r_27__28_, s_r_27__27_, s_r_27__26_, s_r_27__25_, s_r_27__24_, s_r_27__23_, s_r_27__22_, s_r_27__21_, s_r_27__20_, s_r_27__19_, s_r_27__18_, s_r_27__17_, s_r_27__16_, s_r_27__15_, s_r_27__14_, s_r_27__13_, s_r_27__12_, s_r_27__11_, s_r_27__10_, s_r_27__9_, s_r_27__8_, s_r_27__7_, s_r_27__6_, s_r_27__5_, s_r_27__4_, s_r_27__3_, s_r_27__2_, s_r_27__1_, s_r_27__0_ }),
    .c_o(c_r[27]),
    .prod_accum_o({ prod_accum_27__28_, prod_accum_27__27_, prod_accum_27__26_, prod_accum_27__25_, prod_accum_27__24_, prod_accum_27__23_, prod_accum_27__22_, prod_accum_27__21_, prod_accum_27__20_, prod_accum_27__19_, prod_accum_27__18_, prod_accum_27__17_, prod_accum_27__16_, prod_accum_27__15_, prod_accum_27__14_, prod_accum_27__13_, prod_accum_27__12_, prod_accum_27__11_, prod_accum_27__10_, prod_accum_27__9_, prod_accum_27__8_, prod_accum_27__7_, prod_accum_27__6_, prod_accum_27__5_, prod_accum_27__4_, prod_accum_27__3_, prod_accum_27__2_, prod_accum_27__1_, prod_accum_27__0_ })
  );


  bsg_mul_array_row_128_28_0
  genblk1_28__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[3583:3456]),
    .b_i(b_r[3583:3456]),
    .s_i({ s_r_27__127_, s_r_27__126_, s_r_27__125_, s_r_27__124_, s_r_27__123_, s_r_27__122_, s_r_27__121_, s_r_27__120_, s_r_27__119_, s_r_27__118_, s_r_27__117_, s_r_27__116_, s_r_27__115_, s_r_27__114_, s_r_27__113_, s_r_27__112_, s_r_27__111_, s_r_27__110_, s_r_27__109_, s_r_27__108_, s_r_27__107_, s_r_27__106_, s_r_27__105_, s_r_27__104_, s_r_27__103_, s_r_27__102_, s_r_27__101_, s_r_27__100_, s_r_27__99_, s_r_27__98_, s_r_27__97_, s_r_27__96_, s_r_27__95_, s_r_27__94_, s_r_27__93_, s_r_27__92_, s_r_27__91_, s_r_27__90_, s_r_27__89_, s_r_27__88_, s_r_27__87_, s_r_27__86_, s_r_27__85_, s_r_27__84_, s_r_27__83_, s_r_27__82_, s_r_27__81_, s_r_27__80_, s_r_27__79_, s_r_27__78_, s_r_27__77_, s_r_27__76_, s_r_27__75_, s_r_27__74_, s_r_27__73_, s_r_27__72_, s_r_27__71_, s_r_27__70_, s_r_27__69_, s_r_27__68_, s_r_27__67_, s_r_27__66_, s_r_27__65_, s_r_27__64_, s_r_27__63_, s_r_27__62_, s_r_27__61_, s_r_27__60_, s_r_27__59_, s_r_27__58_, s_r_27__57_, s_r_27__56_, s_r_27__55_, s_r_27__54_, s_r_27__53_, s_r_27__52_, s_r_27__51_, s_r_27__50_, s_r_27__49_, s_r_27__48_, s_r_27__47_, s_r_27__46_, s_r_27__45_, s_r_27__44_, s_r_27__43_, s_r_27__42_, s_r_27__41_, s_r_27__40_, s_r_27__39_, s_r_27__38_, s_r_27__37_, s_r_27__36_, s_r_27__35_, s_r_27__34_, s_r_27__33_, s_r_27__32_, s_r_27__31_, s_r_27__30_, s_r_27__29_, s_r_27__28_, s_r_27__27_, s_r_27__26_, s_r_27__25_, s_r_27__24_, s_r_27__23_, s_r_27__22_, s_r_27__21_, s_r_27__20_, s_r_27__19_, s_r_27__18_, s_r_27__17_, s_r_27__16_, s_r_27__15_, s_r_27__14_, s_r_27__13_, s_r_27__12_, s_r_27__11_, s_r_27__10_, s_r_27__9_, s_r_27__8_, s_r_27__7_, s_r_27__6_, s_r_27__5_, s_r_27__4_, s_r_27__3_, s_r_27__2_, s_r_27__1_, s_r_27__0_ }),
    .c_i(c_r[27]),
    .prod_accum_i({ prod_accum_27__28_, prod_accum_27__27_, prod_accum_27__26_, prod_accum_27__25_, prod_accum_27__24_, prod_accum_27__23_, prod_accum_27__22_, prod_accum_27__21_, prod_accum_27__20_, prod_accum_27__19_, prod_accum_27__18_, prod_accum_27__17_, prod_accum_27__16_, prod_accum_27__15_, prod_accum_27__14_, prod_accum_27__13_, prod_accum_27__12_, prod_accum_27__11_, prod_accum_27__10_, prod_accum_27__9_, prod_accum_27__8_, prod_accum_27__7_, prod_accum_27__6_, prod_accum_27__5_, prod_accum_27__4_, prod_accum_27__3_, prod_accum_27__2_, prod_accum_27__1_, prod_accum_27__0_ }),
    .a_o(a_r[3711:3584]),
    .b_o(b_r[3711:3584]),
    .s_o({ s_r_28__127_, s_r_28__126_, s_r_28__125_, s_r_28__124_, s_r_28__123_, s_r_28__122_, s_r_28__121_, s_r_28__120_, s_r_28__119_, s_r_28__118_, s_r_28__117_, s_r_28__116_, s_r_28__115_, s_r_28__114_, s_r_28__113_, s_r_28__112_, s_r_28__111_, s_r_28__110_, s_r_28__109_, s_r_28__108_, s_r_28__107_, s_r_28__106_, s_r_28__105_, s_r_28__104_, s_r_28__103_, s_r_28__102_, s_r_28__101_, s_r_28__100_, s_r_28__99_, s_r_28__98_, s_r_28__97_, s_r_28__96_, s_r_28__95_, s_r_28__94_, s_r_28__93_, s_r_28__92_, s_r_28__91_, s_r_28__90_, s_r_28__89_, s_r_28__88_, s_r_28__87_, s_r_28__86_, s_r_28__85_, s_r_28__84_, s_r_28__83_, s_r_28__82_, s_r_28__81_, s_r_28__80_, s_r_28__79_, s_r_28__78_, s_r_28__77_, s_r_28__76_, s_r_28__75_, s_r_28__74_, s_r_28__73_, s_r_28__72_, s_r_28__71_, s_r_28__70_, s_r_28__69_, s_r_28__68_, s_r_28__67_, s_r_28__66_, s_r_28__65_, s_r_28__64_, s_r_28__63_, s_r_28__62_, s_r_28__61_, s_r_28__60_, s_r_28__59_, s_r_28__58_, s_r_28__57_, s_r_28__56_, s_r_28__55_, s_r_28__54_, s_r_28__53_, s_r_28__52_, s_r_28__51_, s_r_28__50_, s_r_28__49_, s_r_28__48_, s_r_28__47_, s_r_28__46_, s_r_28__45_, s_r_28__44_, s_r_28__43_, s_r_28__42_, s_r_28__41_, s_r_28__40_, s_r_28__39_, s_r_28__38_, s_r_28__37_, s_r_28__36_, s_r_28__35_, s_r_28__34_, s_r_28__33_, s_r_28__32_, s_r_28__31_, s_r_28__30_, s_r_28__29_, s_r_28__28_, s_r_28__27_, s_r_28__26_, s_r_28__25_, s_r_28__24_, s_r_28__23_, s_r_28__22_, s_r_28__21_, s_r_28__20_, s_r_28__19_, s_r_28__18_, s_r_28__17_, s_r_28__16_, s_r_28__15_, s_r_28__14_, s_r_28__13_, s_r_28__12_, s_r_28__11_, s_r_28__10_, s_r_28__9_, s_r_28__8_, s_r_28__7_, s_r_28__6_, s_r_28__5_, s_r_28__4_, s_r_28__3_, s_r_28__2_, s_r_28__1_, s_r_28__0_ }),
    .c_o(c_r[28]),
    .prod_accum_o({ prod_accum_28__29_, prod_accum_28__28_, prod_accum_28__27_, prod_accum_28__26_, prod_accum_28__25_, prod_accum_28__24_, prod_accum_28__23_, prod_accum_28__22_, prod_accum_28__21_, prod_accum_28__20_, prod_accum_28__19_, prod_accum_28__18_, prod_accum_28__17_, prod_accum_28__16_, prod_accum_28__15_, prod_accum_28__14_, prod_accum_28__13_, prod_accum_28__12_, prod_accum_28__11_, prod_accum_28__10_, prod_accum_28__9_, prod_accum_28__8_, prod_accum_28__7_, prod_accum_28__6_, prod_accum_28__5_, prod_accum_28__4_, prod_accum_28__3_, prod_accum_28__2_, prod_accum_28__1_, prod_accum_28__0_ })
  );


  bsg_mul_array_row_128_29_0
  genblk1_29__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[3711:3584]),
    .b_i(b_r[3711:3584]),
    .s_i({ s_r_28__127_, s_r_28__126_, s_r_28__125_, s_r_28__124_, s_r_28__123_, s_r_28__122_, s_r_28__121_, s_r_28__120_, s_r_28__119_, s_r_28__118_, s_r_28__117_, s_r_28__116_, s_r_28__115_, s_r_28__114_, s_r_28__113_, s_r_28__112_, s_r_28__111_, s_r_28__110_, s_r_28__109_, s_r_28__108_, s_r_28__107_, s_r_28__106_, s_r_28__105_, s_r_28__104_, s_r_28__103_, s_r_28__102_, s_r_28__101_, s_r_28__100_, s_r_28__99_, s_r_28__98_, s_r_28__97_, s_r_28__96_, s_r_28__95_, s_r_28__94_, s_r_28__93_, s_r_28__92_, s_r_28__91_, s_r_28__90_, s_r_28__89_, s_r_28__88_, s_r_28__87_, s_r_28__86_, s_r_28__85_, s_r_28__84_, s_r_28__83_, s_r_28__82_, s_r_28__81_, s_r_28__80_, s_r_28__79_, s_r_28__78_, s_r_28__77_, s_r_28__76_, s_r_28__75_, s_r_28__74_, s_r_28__73_, s_r_28__72_, s_r_28__71_, s_r_28__70_, s_r_28__69_, s_r_28__68_, s_r_28__67_, s_r_28__66_, s_r_28__65_, s_r_28__64_, s_r_28__63_, s_r_28__62_, s_r_28__61_, s_r_28__60_, s_r_28__59_, s_r_28__58_, s_r_28__57_, s_r_28__56_, s_r_28__55_, s_r_28__54_, s_r_28__53_, s_r_28__52_, s_r_28__51_, s_r_28__50_, s_r_28__49_, s_r_28__48_, s_r_28__47_, s_r_28__46_, s_r_28__45_, s_r_28__44_, s_r_28__43_, s_r_28__42_, s_r_28__41_, s_r_28__40_, s_r_28__39_, s_r_28__38_, s_r_28__37_, s_r_28__36_, s_r_28__35_, s_r_28__34_, s_r_28__33_, s_r_28__32_, s_r_28__31_, s_r_28__30_, s_r_28__29_, s_r_28__28_, s_r_28__27_, s_r_28__26_, s_r_28__25_, s_r_28__24_, s_r_28__23_, s_r_28__22_, s_r_28__21_, s_r_28__20_, s_r_28__19_, s_r_28__18_, s_r_28__17_, s_r_28__16_, s_r_28__15_, s_r_28__14_, s_r_28__13_, s_r_28__12_, s_r_28__11_, s_r_28__10_, s_r_28__9_, s_r_28__8_, s_r_28__7_, s_r_28__6_, s_r_28__5_, s_r_28__4_, s_r_28__3_, s_r_28__2_, s_r_28__1_, s_r_28__0_ }),
    .c_i(c_r[28]),
    .prod_accum_i({ prod_accum_28__29_, prod_accum_28__28_, prod_accum_28__27_, prod_accum_28__26_, prod_accum_28__25_, prod_accum_28__24_, prod_accum_28__23_, prod_accum_28__22_, prod_accum_28__21_, prod_accum_28__20_, prod_accum_28__19_, prod_accum_28__18_, prod_accum_28__17_, prod_accum_28__16_, prod_accum_28__15_, prod_accum_28__14_, prod_accum_28__13_, prod_accum_28__12_, prod_accum_28__11_, prod_accum_28__10_, prod_accum_28__9_, prod_accum_28__8_, prod_accum_28__7_, prod_accum_28__6_, prod_accum_28__5_, prod_accum_28__4_, prod_accum_28__3_, prod_accum_28__2_, prod_accum_28__1_, prod_accum_28__0_ }),
    .a_o(a_r[3839:3712]),
    .b_o(b_r[3839:3712]),
    .s_o({ s_r_29__127_, s_r_29__126_, s_r_29__125_, s_r_29__124_, s_r_29__123_, s_r_29__122_, s_r_29__121_, s_r_29__120_, s_r_29__119_, s_r_29__118_, s_r_29__117_, s_r_29__116_, s_r_29__115_, s_r_29__114_, s_r_29__113_, s_r_29__112_, s_r_29__111_, s_r_29__110_, s_r_29__109_, s_r_29__108_, s_r_29__107_, s_r_29__106_, s_r_29__105_, s_r_29__104_, s_r_29__103_, s_r_29__102_, s_r_29__101_, s_r_29__100_, s_r_29__99_, s_r_29__98_, s_r_29__97_, s_r_29__96_, s_r_29__95_, s_r_29__94_, s_r_29__93_, s_r_29__92_, s_r_29__91_, s_r_29__90_, s_r_29__89_, s_r_29__88_, s_r_29__87_, s_r_29__86_, s_r_29__85_, s_r_29__84_, s_r_29__83_, s_r_29__82_, s_r_29__81_, s_r_29__80_, s_r_29__79_, s_r_29__78_, s_r_29__77_, s_r_29__76_, s_r_29__75_, s_r_29__74_, s_r_29__73_, s_r_29__72_, s_r_29__71_, s_r_29__70_, s_r_29__69_, s_r_29__68_, s_r_29__67_, s_r_29__66_, s_r_29__65_, s_r_29__64_, s_r_29__63_, s_r_29__62_, s_r_29__61_, s_r_29__60_, s_r_29__59_, s_r_29__58_, s_r_29__57_, s_r_29__56_, s_r_29__55_, s_r_29__54_, s_r_29__53_, s_r_29__52_, s_r_29__51_, s_r_29__50_, s_r_29__49_, s_r_29__48_, s_r_29__47_, s_r_29__46_, s_r_29__45_, s_r_29__44_, s_r_29__43_, s_r_29__42_, s_r_29__41_, s_r_29__40_, s_r_29__39_, s_r_29__38_, s_r_29__37_, s_r_29__36_, s_r_29__35_, s_r_29__34_, s_r_29__33_, s_r_29__32_, s_r_29__31_, s_r_29__30_, s_r_29__29_, s_r_29__28_, s_r_29__27_, s_r_29__26_, s_r_29__25_, s_r_29__24_, s_r_29__23_, s_r_29__22_, s_r_29__21_, s_r_29__20_, s_r_29__19_, s_r_29__18_, s_r_29__17_, s_r_29__16_, s_r_29__15_, s_r_29__14_, s_r_29__13_, s_r_29__12_, s_r_29__11_, s_r_29__10_, s_r_29__9_, s_r_29__8_, s_r_29__7_, s_r_29__6_, s_r_29__5_, s_r_29__4_, s_r_29__3_, s_r_29__2_, s_r_29__1_, s_r_29__0_ }),
    .c_o(c_r[29]),
    .prod_accum_o({ prod_accum_29__30_, prod_accum_29__29_, prod_accum_29__28_, prod_accum_29__27_, prod_accum_29__26_, prod_accum_29__25_, prod_accum_29__24_, prod_accum_29__23_, prod_accum_29__22_, prod_accum_29__21_, prod_accum_29__20_, prod_accum_29__19_, prod_accum_29__18_, prod_accum_29__17_, prod_accum_29__16_, prod_accum_29__15_, prod_accum_29__14_, prod_accum_29__13_, prod_accum_29__12_, prod_accum_29__11_, prod_accum_29__10_, prod_accum_29__9_, prod_accum_29__8_, prod_accum_29__7_, prod_accum_29__6_, prod_accum_29__5_, prod_accum_29__4_, prod_accum_29__3_, prod_accum_29__2_, prod_accum_29__1_, prod_accum_29__0_ })
  );


  bsg_mul_array_row_128_30_0
  genblk1_30__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[3839:3712]),
    .b_i(b_r[3839:3712]),
    .s_i({ s_r_29__127_, s_r_29__126_, s_r_29__125_, s_r_29__124_, s_r_29__123_, s_r_29__122_, s_r_29__121_, s_r_29__120_, s_r_29__119_, s_r_29__118_, s_r_29__117_, s_r_29__116_, s_r_29__115_, s_r_29__114_, s_r_29__113_, s_r_29__112_, s_r_29__111_, s_r_29__110_, s_r_29__109_, s_r_29__108_, s_r_29__107_, s_r_29__106_, s_r_29__105_, s_r_29__104_, s_r_29__103_, s_r_29__102_, s_r_29__101_, s_r_29__100_, s_r_29__99_, s_r_29__98_, s_r_29__97_, s_r_29__96_, s_r_29__95_, s_r_29__94_, s_r_29__93_, s_r_29__92_, s_r_29__91_, s_r_29__90_, s_r_29__89_, s_r_29__88_, s_r_29__87_, s_r_29__86_, s_r_29__85_, s_r_29__84_, s_r_29__83_, s_r_29__82_, s_r_29__81_, s_r_29__80_, s_r_29__79_, s_r_29__78_, s_r_29__77_, s_r_29__76_, s_r_29__75_, s_r_29__74_, s_r_29__73_, s_r_29__72_, s_r_29__71_, s_r_29__70_, s_r_29__69_, s_r_29__68_, s_r_29__67_, s_r_29__66_, s_r_29__65_, s_r_29__64_, s_r_29__63_, s_r_29__62_, s_r_29__61_, s_r_29__60_, s_r_29__59_, s_r_29__58_, s_r_29__57_, s_r_29__56_, s_r_29__55_, s_r_29__54_, s_r_29__53_, s_r_29__52_, s_r_29__51_, s_r_29__50_, s_r_29__49_, s_r_29__48_, s_r_29__47_, s_r_29__46_, s_r_29__45_, s_r_29__44_, s_r_29__43_, s_r_29__42_, s_r_29__41_, s_r_29__40_, s_r_29__39_, s_r_29__38_, s_r_29__37_, s_r_29__36_, s_r_29__35_, s_r_29__34_, s_r_29__33_, s_r_29__32_, s_r_29__31_, s_r_29__30_, s_r_29__29_, s_r_29__28_, s_r_29__27_, s_r_29__26_, s_r_29__25_, s_r_29__24_, s_r_29__23_, s_r_29__22_, s_r_29__21_, s_r_29__20_, s_r_29__19_, s_r_29__18_, s_r_29__17_, s_r_29__16_, s_r_29__15_, s_r_29__14_, s_r_29__13_, s_r_29__12_, s_r_29__11_, s_r_29__10_, s_r_29__9_, s_r_29__8_, s_r_29__7_, s_r_29__6_, s_r_29__5_, s_r_29__4_, s_r_29__3_, s_r_29__2_, s_r_29__1_, s_r_29__0_ }),
    .c_i(c_r[29]),
    .prod_accum_i({ prod_accum_29__30_, prod_accum_29__29_, prod_accum_29__28_, prod_accum_29__27_, prod_accum_29__26_, prod_accum_29__25_, prod_accum_29__24_, prod_accum_29__23_, prod_accum_29__22_, prod_accum_29__21_, prod_accum_29__20_, prod_accum_29__19_, prod_accum_29__18_, prod_accum_29__17_, prod_accum_29__16_, prod_accum_29__15_, prod_accum_29__14_, prod_accum_29__13_, prod_accum_29__12_, prod_accum_29__11_, prod_accum_29__10_, prod_accum_29__9_, prod_accum_29__8_, prod_accum_29__7_, prod_accum_29__6_, prod_accum_29__5_, prod_accum_29__4_, prod_accum_29__3_, prod_accum_29__2_, prod_accum_29__1_, prod_accum_29__0_ }),
    .a_o(a_r[3967:3840]),
    .b_o(b_r[3967:3840]),
    .s_o({ s_r_30__127_, s_r_30__126_, s_r_30__125_, s_r_30__124_, s_r_30__123_, s_r_30__122_, s_r_30__121_, s_r_30__120_, s_r_30__119_, s_r_30__118_, s_r_30__117_, s_r_30__116_, s_r_30__115_, s_r_30__114_, s_r_30__113_, s_r_30__112_, s_r_30__111_, s_r_30__110_, s_r_30__109_, s_r_30__108_, s_r_30__107_, s_r_30__106_, s_r_30__105_, s_r_30__104_, s_r_30__103_, s_r_30__102_, s_r_30__101_, s_r_30__100_, s_r_30__99_, s_r_30__98_, s_r_30__97_, s_r_30__96_, s_r_30__95_, s_r_30__94_, s_r_30__93_, s_r_30__92_, s_r_30__91_, s_r_30__90_, s_r_30__89_, s_r_30__88_, s_r_30__87_, s_r_30__86_, s_r_30__85_, s_r_30__84_, s_r_30__83_, s_r_30__82_, s_r_30__81_, s_r_30__80_, s_r_30__79_, s_r_30__78_, s_r_30__77_, s_r_30__76_, s_r_30__75_, s_r_30__74_, s_r_30__73_, s_r_30__72_, s_r_30__71_, s_r_30__70_, s_r_30__69_, s_r_30__68_, s_r_30__67_, s_r_30__66_, s_r_30__65_, s_r_30__64_, s_r_30__63_, s_r_30__62_, s_r_30__61_, s_r_30__60_, s_r_30__59_, s_r_30__58_, s_r_30__57_, s_r_30__56_, s_r_30__55_, s_r_30__54_, s_r_30__53_, s_r_30__52_, s_r_30__51_, s_r_30__50_, s_r_30__49_, s_r_30__48_, s_r_30__47_, s_r_30__46_, s_r_30__45_, s_r_30__44_, s_r_30__43_, s_r_30__42_, s_r_30__41_, s_r_30__40_, s_r_30__39_, s_r_30__38_, s_r_30__37_, s_r_30__36_, s_r_30__35_, s_r_30__34_, s_r_30__33_, s_r_30__32_, s_r_30__31_, s_r_30__30_, s_r_30__29_, s_r_30__28_, s_r_30__27_, s_r_30__26_, s_r_30__25_, s_r_30__24_, s_r_30__23_, s_r_30__22_, s_r_30__21_, s_r_30__20_, s_r_30__19_, s_r_30__18_, s_r_30__17_, s_r_30__16_, s_r_30__15_, s_r_30__14_, s_r_30__13_, s_r_30__12_, s_r_30__11_, s_r_30__10_, s_r_30__9_, s_r_30__8_, s_r_30__7_, s_r_30__6_, s_r_30__5_, s_r_30__4_, s_r_30__3_, s_r_30__2_, s_r_30__1_, s_r_30__0_ }),
    .c_o(c_r[30]),
    .prod_accum_o({ prod_accum_30__31_, prod_accum_30__30_, prod_accum_30__29_, prod_accum_30__28_, prod_accum_30__27_, prod_accum_30__26_, prod_accum_30__25_, prod_accum_30__24_, prod_accum_30__23_, prod_accum_30__22_, prod_accum_30__21_, prod_accum_30__20_, prod_accum_30__19_, prod_accum_30__18_, prod_accum_30__17_, prod_accum_30__16_, prod_accum_30__15_, prod_accum_30__14_, prod_accum_30__13_, prod_accum_30__12_, prod_accum_30__11_, prod_accum_30__10_, prod_accum_30__9_, prod_accum_30__8_, prod_accum_30__7_, prod_accum_30__6_, prod_accum_30__5_, prod_accum_30__4_, prod_accum_30__3_, prod_accum_30__2_, prod_accum_30__1_, prod_accum_30__0_ })
  );


  bsg_mul_array_row_128_31_1
  genblk1_31__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[3967:3840]),
    .b_i(b_r[3967:3840]),
    .s_i({ s_r_30__127_, s_r_30__126_, s_r_30__125_, s_r_30__124_, s_r_30__123_, s_r_30__122_, s_r_30__121_, s_r_30__120_, s_r_30__119_, s_r_30__118_, s_r_30__117_, s_r_30__116_, s_r_30__115_, s_r_30__114_, s_r_30__113_, s_r_30__112_, s_r_30__111_, s_r_30__110_, s_r_30__109_, s_r_30__108_, s_r_30__107_, s_r_30__106_, s_r_30__105_, s_r_30__104_, s_r_30__103_, s_r_30__102_, s_r_30__101_, s_r_30__100_, s_r_30__99_, s_r_30__98_, s_r_30__97_, s_r_30__96_, s_r_30__95_, s_r_30__94_, s_r_30__93_, s_r_30__92_, s_r_30__91_, s_r_30__90_, s_r_30__89_, s_r_30__88_, s_r_30__87_, s_r_30__86_, s_r_30__85_, s_r_30__84_, s_r_30__83_, s_r_30__82_, s_r_30__81_, s_r_30__80_, s_r_30__79_, s_r_30__78_, s_r_30__77_, s_r_30__76_, s_r_30__75_, s_r_30__74_, s_r_30__73_, s_r_30__72_, s_r_30__71_, s_r_30__70_, s_r_30__69_, s_r_30__68_, s_r_30__67_, s_r_30__66_, s_r_30__65_, s_r_30__64_, s_r_30__63_, s_r_30__62_, s_r_30__61_, s_r_30__60_, s_r_30__59_, s_r_30__58_, s_r_30__57_, s_r_30__56_, s_r_30__55_, s_r_30__54_, s_r_30__53_, s_r_30__52_, s_r_30__51_, s_r_30__50_, s_r_30__49_, s_r_30__48_, s_r_30__47_, s_r_30__46_, s_r_30__45_, s_r_30__44_, s_r_30__43_, s_r_30__42_, s_r_30__41_, s_r_30__40_, s_r_30__39_, s_r_30__38_, s_r_30__37_, s_r_30__36_, s_r_30__35_, s_r_30__34_, s_r_30__33_, s_r_30__32_, s_r_30__31_, s_r_30__30_, s_r_30__29_, s_r_30__28_, s_r_30__27_, s_r_30__26_, s_r_30__25_, s_r_30__24_, s_r_30__23_, s_r_30__22_, s_r_30__21_, s_r_30__20_, s_r_30__19_, s_r_30__18_, s_r_30__17_, s_r_30__16_, s_r_30__15_, s_r_30__14_, s_r_30__13_, s_r_30__12_, s_r_30__11_, s_r_30__10_, s_r_30__9_, s_r_30__8_, s_r_30__7_, s_r_30__6_, s_r_30__5_, s_r_30__4_, s_r_30__3_, s_r_30__2_, s_r_30__1_, s_r_30__0_ }),
    .c_i(c_r[30]),
    .prod_accum_i({ prod_accum_30__31_, prod_accum_30__30_, prod_accum_30__29_, prod_accum_30__28_, prod_accum_30__27_, prod_accum_30__26_, prod_accum_30__25_, prod_accum_30__24_, prod_accum_30__23_, prod_accum_30__22_, prod_accum_30__21_, prod_accum_30__20_, prod_accum_30__19_, prod_accum_30__18_, prod_accum_30__17_, prod_accum_30__16_, prod_accum_30__15_, prod_accum_30__14_, prod_accum_30__13_, prod_accum_30__12_, prod_accum_30__11_, prod_accum_30__10_, prod_accum_30__9_, prod_accum_30__8_, prod_accum_30__7_, prod_accum_30__6_, prod_accum_30__5_, prod_accum_30__4_, prod_accum_30__3_, prod_accum_30__2_, prod_accum_30__1_, prod_accum_30__0_ }),
    .a_o(a_r[4095:3968]),
    .b_o(b_r[4095:3968]),
    .s_o({ s_r_31__127_, s_r_31__126_, s_r_31__125_, s_r_31__124_, s_r_31__123_, s_r_31__122_, s_r_31__121_, s_r_31__120_, s_r_31__119_, s_r_31__118_, s_r_31__117_, s_r_31__116_, s_r_31__115_, s_r_31__114_, s_r_31__113_, s_r_31__112_, s_r_31__111_, s_r_31__110_, s_r_31__109_, s_r_31__108_, s_r_31__107_, s_r_31__106_, s_r_31__105_, s_r_31__104_, s_r_31__103_, s_r_31__102_, s_r_31__101_, s_r_31__100_, s_r_31__99_, s_r_31__98_, s_r_31__97_, s_r_31__96_, s_r_31__95_, s_r_31__94_, s_r_31__93_, s_r_31__92_, s_r_31__91_, s_r_31__90_, s_r_31__89_, s_r_31__88_, s_r_31__87_, s_r_31__86_, s_r_31__85_, s_r_31__84_, s_r_31__83_, s_r_31__82_, s_r_31__81_, s_r_31__80_, s_r_31__79_, s_r_31__78_, s_r_31__77_, s_r_31__76_, s_r_31__75_, s_r_31__74_, s_r_31__73_, s_r_31__72_, s_r_31__71_, s_r_31__70_, s_r_31__69_, s_r_31__68_, s_r_31__67_, s_r_31__66_, s_r_31__65_, s_r_31__64_, s_r_31__63_, s_r_31__62_, s_r_31__61_, s_r_31__60_, s_r_31__59_, s_r_31__58_, s_r_31__57_, s_r_31__56_, s_r_31__55_, s_r_31__54_, s_r_31__53_, s_r_31__52_, s_r_31__51_, s_r_31__50_, s_r_31__49_, s_r_31__48_, s_r_31__47_, s_r_31__46_, s_r_31__45_, s_r_31__44_, s_r_31__43_, s_r_31__42_, s_r_31__41_, s_r_31__40_, s_r_31__39_, s_r_31__38_, s_r_31__37_, s_r_31__36_, s_r_31__35_, s_r_31__34_, s_r_31__33_, s_r_31__32_, s_r_31__31_, s_r_31__30_, s_r_31__29_, s_r_31__28_, s_r_31__27_, s_r_31__26_, s_r_31__25_, s_r_31__24_, s_r_31__23_, s_r_31__22_, s_r_31__21_, s_r_31__20_, s_r_31__19_, s_r_31__18_, s_r_31__17_, s_r_31__16_, s_r_31__15_, s_r_31__14_, s_r_31__13_, s_r_31__12_, s_r_31__11_, s_r_31__10_, s_r_31__9_, s_r_31__8_, s_r_31__7_, s_r_31__6_, s_r_31__5_, s_r_31__4_, s_r_31__3_, s_r_31__2_, s_r_31__1_, s_r_31__0_ }),
    .c_o(c_r[31]),
    .prod_accum_o({ prod_accum_31__32_, prod_accum_31__31_, prod_accum_31__30_, prod_accum_31__29_, prod_accum_31__28_, prod_accum_31__27_, prod_accum_31__26_, prod_accum_31__25_, prod_accum_31__24_, prod_accum_31__23_, prod_accum_31__22_, prod_accum_31__21_, prod_accum_31__20_, prod_accum_31__19_, prod_accum_31__18_, prod_accum_31__17_, prod_accum_31__16_, prod_accum_31__15_, prod_accum_31__14_, prod_accum_31__13_, prod_accum_31__12_, prod_accum_31__11_, prod_accum_31__10_, prod_accum_31__9_, prod_accum_31__8_, prod_accum_31__7_, prod_accum_31__6_, prod_accum_31__5_, prod_accum_31__4_, prod_accum_31__3_, prod_accum_31__2_, prod_accum_31__1_, prod_accum_31__0_ })
  );


  bsg_mul_array_row_128_32_x
  genblk1_32__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[4095:3968]),
    .b_i(b_r[4095:3968]),
    .s_i({ s_r_31__127_, s_r_31__126_, s_r_31__125_, s_r_31__124_, s_r_31__123_, s_r_31__122_, s_r_31__121_, s_r_31__120_, s_r_31__119_, s_r_31__118_, s_r_31__117_, s_r_31__116_, s_r_31__115_, s_r_31__114_, s_r_31__113_, s_r_31__112_, s_r_31__111_, s_r_31__110_, s_r_31__109_, s_r_31__108_, s_r_31__107_, s_r_31__106_, s_r_31__105_, s_r_31__104_, s_r_31__103_, s_r_31__102_, s_r_31__101_, s_r_31__100_, s_r_31__99_, s_r_31__98_, s_r_31__97_, s_r_31__96_, s_r_31__95_, s_r_31__94_, s_r_31__93_, s_r_31__92_, s_r_31__91_, s_r_31__90_, s_r_31__89_, s_r_31__88_, s_r_31__87_, s_r_31__86_, s_r_31__85_, s_r_31__84_, s_r_31__83_, s_r_31__82_, s_r_31__81_, s_r_31__80_, s_r_31__79_, s_r_31__78_, s_r_31__77_, s_r_31__76_, s_r_31__75_, s_r_31__74_, s_r_31__73_, s_r_31__72_, s_r_31__71_, s_r_31__70_, s_r_31__69_, s_r_31__68_, s_r_31__67_, s_r_31__66_, s_r_31__65_, s_r_31__64_, s_r_31__63_, s_r_31__62_, s_r_31__61_, s_r_31__60_, s_r_31__59_, s_r_31__58_, s_r_31__57_, s_r_31__56_, s_r_31__55_, s_r_31__54_, s_r_31__53_, s_r_31__52_, s_r_31__51_, s_r_31__50_, s_r_31__49_, s_r_31__48_, s_r_31__47_, s_r_31__46_, s_r_31__45_, s_r_31__44_, s_r_31__43_, s_r_31__42_, s_r_31__41_, s_r_31__40_, s_r_31__39_, s_r_31__38_, s_r_31__37_, s_r_31__36_, s_r_31__35_, s_r_31__34_, s_r_31__33_, s_r_31__32_, s_r_31__31_, s_r_31__30_, s_r_31__29_, s_r_31__28_, s_r_31__27_, s_r_31__26_, s_r_31__25_, s_r_31__24_, s_r_31__23_, s_r_31__22_, s_r_31__21_, s_r_31__20_, s_r_31__19_, s_r_31__18_, s_r_31__17_, s_r_31__16_, s_r_31__15_, s_r_31__14_, s_r_31__13_, s_r_31__12_, s_r_31__11_, s_r_31__10_, s_r_31__9_, s_r_31__8_, s_r_31__7_, s_r_31__6_, s_r_31__5_, s_r_31__4_, s_r_31__3_, s_r_31__2_, s_r_31__1_, s_r_31__0_ }),
    .c_i(c_r[31]),
    .prod_accum_i({ prod_accum_31__32_, prod_accum_31__31_, prod_accum_31__30_, prod_accum_31__29_, prod_accum_31__28_, prod_accum_31__27_, prod_accum_31__26_, prod_accum_31__25_, prod_accum_31__24_, prod_accum_31__23_, prod_accum_31__22_, prod_accum_31__21_, prod_accum_31__20_, prod_accum_31__19_, prod_accum_31__18_, prod_accum_31__17_, prod_accum_31__16_, prod_accum_31__15_, prod_accum_31__14_, prod_accum_31__13_, prod_accum_31__12_, prod_accum_31__11_, prod_accum_31__10_, prod_accum_31__9_, prod_accum_31__8_, prod_accum_31__7_, prod_accum_31__6_, prod_accum_31__5_, prod_accum_31__4_, prod_accum_31__3_, prod_accum_31__2_, prod_accum_31__1_, prod_accum_31__0_ }),
    .a_o(a_r[4223:4096]),
    .b_o(b_r[4223:4096]),
    .s_o({ s_r_32__127_, s_r_32__126_, s_r_32__125_, s_r_32__124_, s_r_32__123_, s_r_32__122_, s_r_32__121_, s_r_32__120_, s_r_32__119_, s_r_32__118_, s_r_32__117_, s_r_32__116_, s_r_32__115_, s_r_32__114_, s_r_32__113_, s_r_32__112_, s_r_32__111_, s_r_32__110_, s_r_32__109_, s_r_32__108_, s_r_32__107_, s_r_32__106_, s_r_32__105_, s_r_32__104_, s_r_32__103_, s_r_32__102_, s_r_32__101_, s_r_32__100_, s_r_32__99_, s_r_32__98_, s_r_32__97_, s_r_32__96_, s_r_32__95_, s_r_32__94_, s_r_32__93_, s_r_32__92_, s_r_32__91_, s_r_32__90_, s_r_32__89_, s_r_32__88_, s_r_32__87_, s_r_32__86_, s_r_32__85_, s_r_32__84_, s_r_32__83_, s_r_32__82_, s_r_32__81_, s_r_32__80_, s_r_32__79_, s_r_32__78_, s_r_32__77_, s_r_32__76_, s_r_32__75_, s_r_32__74_, s_r_32__73_, s_r_32__72_, s_r_32__71_, s_r_32__70_, s_r_32__69_, s_r_32__68_, s_r_32__67_, s_r_32__66_, s_r_32__65_, s_r_32__64_, s_r_32__63_, s_r_32__62_, s_r_32__61_, s_r_32__60_, s_r_32__59_, s_r_32__58_, s_r_32__57_, s_r_32__56_, s_r_32__55_, s_r_32__54_, s_r_32__53_, s_r_32__52_, s_r_32__51_, s_r_32__50_, s_r_32__49_, s_r_32__48_, s_r_32__47_, s_r_32__46_, s_r_32__45_, s_r_32__44_, s_r_32__43_, s_r_32__42_, s_r_32__41_, s_r_32__40_, s_r_32__39_, s_r_32__38_, s_r_32__37_, s_r_32__36_, s_r_32__35_, s_r_32__34_, s_r_32__33_, s_r_32__32_, s_r_32__31_, s_r_32__30_, s_r_32__29_, s_r_32__28_, s_r_32__27_, s_r_32__26_, s_r_32__25_, s_r_32__24_, s_r_32__23_, s_r_32__22_, s_r_32__21_, s_r_32__20_, s_r_32__19_, s_r_32__18_, s_r_32__17_, s_r_32__16_, s_r_32__15_, s_r_32__14_, s_r_32__13_, s_r_32__12_, s_r_32__11_, s_r_32__10_, s_r_32__9_, s_r_32__8_, s_r_32__7_, s_r_32__6_, s_r_32__5_, s_r_32__4_, s_r_32__3_, s_r_32__2_, s_r_32__1_, s_r_32__0_ }),
    .c_o(c_r[32]),
    .prod_accum_o({ prod_accum_32__33_, prod_accum_32__32_, prod_accum_32__31_, prod_accum_32__30_, prod_accum_32__29_, prod_accum_32__28_, prod_accum_32__27_, prod_accum_32__26_, prod_accum_32__25_, prod_accum_32__24_, prod_accum_32__23_, prod_accum_32__22_, prod_accum_32__21_, prod_accum_32__20_, prod_accum_32__19_, prod_accum_32__18_, prod_accum_32__17_, prod_accum_32__16_, prod_accum_32__15_, prod_accum_32__14_, prod_accum_32__13_, prod_accum_32__12_, prod_accum_32__11_, prod_accum_32__10_, prod_accum_32__9_, prod_accum_32__8_, prod_accum_32__7_, prod_accum_32__6_, prod_accum_32__5_, prod_accum_32__4_, prod_accum_32__3_, prod_accum_32__2_, prod_accum_32__1_, prod_accum_32__0_ })
  );


  bsg_mul_array_row_128_33_x
  genblk1_33__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[4223:4096]),
    .b_i(b_r[4223:4096]),
    .s_i({ s_r_32__127_, s_r_32__126_, s_r_32__125_, s_r_32__124_, s_r_32__123_, s_r_32__122_, s_r_32__121_, s_r_32__120_, s_r_32__119_, s_r_32__118_, s_r_32__117_, s_r_32__116_, s_r_32__115_, s_r_32__114_, s_r_32__113_, s_r_32__112_, s_r_32__111_, s_r_32__110_, s_r_32__109_, s_r_32__108_, s_r_32__107_, s_r_32__106_, s_r_32__105_, s_r_32__104_, s_r_32__103_, s_r_32__102_, s_r_32__101_, s_r_32__100_, s_r_32__99_, s_r_32__98_, s_r_32__97_, s_r_32__96_, s_r_32__95_, s_r_32__94_, s_r_32__93_, s_r_32__92_, s_r_32__91_, s_r_32__90_, s_r_32__89_, s_r_32__88_, s_r_32__87_, s_r_32__86_, s_r_32__85_, s_r_32__84_, s_r_32__83_, s_r_32__82_, s_r_32__81_, s_r_32__80_, s_r_32__79_, s_r_32__78_, s_r_32__77_, s_r_32__76_, s_r_32__75_, s_r_32__74_, s_r_32__73_, s_r_32__72_, s_r_32__71_, s_r_32__70_, s_r_32__69_, s_r_32__68_, s_r_32__67_, s_r_32__66_, s_r_32__65_, s_r_32__64_, s_r_32__63_, s_r_32__62_, s_r_32__61_, s_r_32__60_, s_r_32__59_, s_r_32__58_, s_r_32__57_, s_r_32__56_, s_r_32__55_, s_r_32__54_, s_r_32__53_, s_r_32__52_, s_r_32__51_, s_r_32__50_, s_r_32__49_, s_r_32__48_, s_r_32__47_, s_r_32__46_, s_r_32__45_, s_r_32__44_, s_r_32__43_, s_r_32__42_, s_r_32__41_, s_r_32__40_, s_r_32__39_, s_r_32__38_, s_r_32__37_, s_r_32__36_, s_r_32__35_, s_r_32__34_, s_r_32__33_, s_r_32__32_, s_r_32__31_, s_r_32__30_, s_r_32__29_, s_r_32__28_, s_r_32__27_, s_r_32__26_, s_r_32__25_, s_r_32__24_, s_r_32__23_, s_r_32__22_, s_r_32__21_, s_r_32__20_, s_r_32__19_, s_r_32__18_, s_r_32__17_, s_r_32__16_, s_r_32__15_, s_r_32__14_, s_r_32__13_, s_r_32__12_, s_r_32__11_, s_r_32__10_, s_r_32__9_, s_r_32__8_, s_r_32__7_, s_r_32__6_, s_r_32__5_, s_r_32__4_, s_r_32__3_, s_r_32__2_, s_r_32__1_, s_r_32__0_ }),
    .c_i(c_r[32]),
    .prod_accum_i({ prod_accum_32__33_, prod_accum_32__32_, prod_accum_32__31_, prod_accum_32__30_, prod_accum_32__29_, prod_accum_32__28_, prod_accum_32__27_, prod_accum_32__26_, prod_accum_32__25_, prod_accum_32__24_, prod_accum_32__23_, prod_accum_32__22_, prod_accum_32__21_, prod_accum_32__20_, prod_accum_32__19_, prod_accum_32__18_, prod_accum_32__17_, prod_accum_32__16_, prod_accum_32__15_, prod_accum_32__14_, prod_accum_32__13_, prod_accum_32__12_, prod_accum_32__11_, prod_accum_32__10_, prod_accum_32__9_, prod_accum_32__8_, prod_accum_32__7_, prod_accum_32__6_, prod_accum_32__5_, prod_accum_32__4_, prod_accum_32__3_, prod_accum_32__2_, prod_accum_32__1_, prod_accum_32__0_ }),
    .a_o(a_r[4351:4224]),
    .b_o(b_r[4351:4224]),
    .s_o({ s_r_33__127_, s_r_33__126_, s_r_33__125_, s_r_33__124_, s_r_33__123_, s_r_33__122_, s_r_33__121_, s_r_33__120_, s_r_33__119_, s_r_33__118_, s_r_33__117_, s_r_33__116_, s_r_33__115_, s_r_33__114_, s_r_33__113_, s_r_33__112_, s_r_33__111_, s_r_33__110_, s_r_33__109_, s_r_33__108_, s_r_33__107_, s_r_33__106_, s_r_33__105_, s_r_33__104_, s_r_33__103_, s_r_33__102_, s_r_33__101_, s_r_33__100_, s_r_33__99_, s_r_33__98_, s_r_33__97_, s_r_33__96_, s_r_33__95_, s_r_33__94_, s_r_33__93_, s_r_33__92_, s_r_33__91_, s_r_33__90_, s_r_33__89_, s_r_33__88_, s_r_33__87_, s_r_33__86_, s_r_33__85_, s_r_33__84_, s_r_33__83_, s_r_33__82_, s_r_33__81_, s_r_33__80_, s_r_33__79_, s_r_33__78_, s_r_33__77_, s_r_33__76_, s_r_33__75_, s_r_33__74_, s_r_33__73_, s_r_33__72_, s_r_33__71_, s_r_33__70_, s_r_33__69_, s_r_33__68_, s_r_33__67_, s_r_33__66_, s_r_33__65_, s_r_33__64_, s_r_33__63_, s_r_33__62_, s_r_33__61_, s_r_33__60_, s_r_33__59_, s_r_33__58_, s_r_33__57_, s_r_33__56_, s_r_33__55_, s_r_33__54_, s_r_33__53_, s_r_33__52_, s_r_33__51_, s_r_33__50_, s_r_33__49_, s_r_33__48_, s_r_33__47_, s_r_33__46_, s_r_33__45_, s_r_33__44_, s_r_33__43_, s_r_33__42_, s_r_33__41_, s_r_33__40_, s_r_33__39_, s_r_33__38_, s_r_33__37_, s_r_33__36_, s_r_33__35_, s_r_33__34_, s_r_33__33_, s_r_33__32_, s_r_33__31_, s_r_33__30_, s_r_33__29_, s_r_33__28_, s_r_33__27_, s_r_33__26_, s_r_33__25_, s_r_33__24_, s_r_33__23_, s_r_33__22_, s_r_33__21_, s_r_33__20_, s_r_33__19_, s_r_33__18_, s_r_33__17_, s_r_33__16_, s_r_33__15_, s_r_33__14_, s_r_33__13_, s_r_33__12_, s_r_33__11_, s_r_33__10_, s_r_33__9_, s_r_33__8_, s_r_33__7_, s_r_33__6_, s_r_33__5_, s_r_33__4_, s_r_33__3_, s_r_33__2_, s_r_33__1_, s_r_33__0_ }),
    .c_o(c_r[33]),
    .prod_accum_o({ prod_accum_33__34_, prod_accum_33__33_, prod_accum_33__32_, prod_accum_33__31_, prod_accum_33__30_, prod_accum_33__29_, prod_accum_33__28_, prod_accum_33__27_, prod_accum_33__26_, prod_accum_33__25_, prod_accum_33__24_, prod_accum_33__23_, prod_accum_33__22_, prod_accum_33__21_, prod_accum_33__20_, prod_accum_33__19_, prod_accum_33__18_, prod_accum_33__17_, prod_accum_33__16_, prod_accum_33__15_, prod_accum_33__14_, prod_accum_33__13_, prod_accum_33__12_, prod_accum_33__11_, prod_accum_33__10_, prod_accum_33__9_, prod_accum_33__8_, prod_accum_33__7_, prod_accum_33__6_, prod_accum_33__5_, prod_accum_33__4_, prod_accum_33__3_, prod_accum_33__2_, prod_accum_33__1_, prod_accum_33__0_ })
  );


  bsg_mul_array_row_128_34_x
  genblk1_34__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[4351:4224]),
    .b_i(b_r[4351:4224]),
    .s_i({ s_r_33__127_, s_r_33__126_, s_r_33__125_, s_r_33__124_, s_r_33__123_, s_r_33__122_, s_r_33__121_, s_r_33__120_, s_r_33__119_, s_r_33__118_, s_r_33__117_, s_r_33__116_, s_r_33__115_, s_r_33__114_, s_r_33__113_, s_r_33__112_, s_r_33__111_, s_r_33__110_, s_r_33__109_, s_r_33__108_, s_r_33__107_, s_r_33__106_, s_r_33__105_, s_r_33__104_, s_r_33__103_, s_r_33__102_, s_r_33__101_, s_r_33__100_, s_r_33__99_, s_r_33__98_, s_r_33__97_, s_r_33__96_, s_r_33__95_, s_r_33__94_, s_r_33__93_, s_r_33__92_, s_r_33__91_, s_r_33__90_, s_r_33__89_, s_r_33__88_, s_r_33__87_, s_r_33__86_, s_r_33__85_, s_r_33__84_, s_r_33__83_, s_r_33__82_, s_r_33__81_, s_r_33__80_, s_r_33__79_, s_r_33__78_, s_r_33__77_, s_r_33__76_, s_r_33__75_, s_r_33__74_, s_r_33__73_, s_r_33__72_, s_r_33__71_, s_r_33__70_, s_r_33__69_, s_r_33__68_, s_r_33__67_, s_r_33__66_, s_r_33__65_, s_r_33__64_, s_r_33__63_, s_r_33__62_, s_r_33__61_, s_r_33__60_, s_r_33__59_, s_r_33__58_, s_r_33__57_, s_r_33__56_, s_r_33__55_, s_r_33__54_, s_r_33__53_, s_r_33__52_, s_r_33__51_, s_r_33__50_, s_r_33__49_, s_r_33__48_, s_r_33__47_, s_r_33__46_, s_r_33__45_, s_r_33__44_, s_r_33__43_, s_r_33__42_, s_r_33__41_, s_r_33__40_, s_r_33__39_, s_r_33__38_, s_r_33__37_, s_r_33__36_, s_r_33__35_, s_r_33__34_, s_r_33__33_, s_r_33__32_, s_r_33__31_, s_r_33__30_, s_r_33__29_, s_r_33__28_, s_r_33__27_, s_r_33__26_, s_r_33__25_, s_r_33__24_, s_r_33__23_, s_r_33__22_, s_r_33__21_, s_r_33__20_, s_r_33__19_, s_r_33__18_, s_r_33__17_, s_r_33__16_, s_r_33__15_, s_r_33__14_, s_r_33__13_, s_r_33__12_, s_r_33__11_, s_r_33__10_, s_r_33__9_, s_r_33__8_, s_r_33__7_, s_r_33__6_, s_r_33__5_, s_r_33__4_, s_r_33__3_, s_r_33__2_, s_r_33__1_, s_r_33__0_ }),
    .c_i(c_r[33]),
    .prod_accum_i({ prod_accum_33__34_, prod_accum_33__33_, prod_accum_33__32_, prod_accum_33__31_, prod_accum_33__30_, prod_accum_33__29_, prod_accum_33__28_, prod_accum_33__27_, prod_accum_33__26_, prod_accum_33__25_, prod_accum_33__24_, prod_accum_33__23_, prod_accum_33__22_, prod_accum_33__21_, prod_accum_33__20_, prod_accum_33__19_, prod_accum_33__18_, prod_accum_33__17_, prod_accum_33__16_, prod_accum_33__15_, prod_accum_33__14_, prod_accum_33__13_, prod_accum_33__12_, prod_accum_33__11_, prod_accum_33__10_, prod_accum_33__9_, prod_accum_33__8_, prod_accum_33__7_, prod_accum_33__6_, prod_accum_33__5_, prod_accum_33__4_, prod_accum_33__3_, prod_accum_33__2_, prod_accum_33__1_, prod_accum_33__0_ }),
    .a_o(a_r[4479:4352]),
    .b_o(b_r[4479:4352]),
    .s_o({ s_r_34__127_, s_r_34__126_, s_r_34__125_, s_r_34__124_, s_r_34__123_, s_r_34__122_, s_r_34__121_, s_r_34__120_, s_r_34__119_, s_r_34__118_, s_r_34__117_, s_r_34__116_, s_r_34__115_, s_r_34__114_, s_r_34__113_, s_r_34__112_, s_r_34__111_, s_r_34__110_, s_r_34__109_, s_r_34__108_, s_r_34__107_, s_r_34__106_, s_r_34__105_, s_r_34__104_, s_r_34__103_, s_r_34__102_, s_r_34__101_, s_r_34__100_, s_r_34__99_, s_r_34__98_, s_r_34__97_, s_r_34__96_, s_r_34__95_, s_r_34__94_, s_r_34__93_, s_r_34__92_, s_r_34__91_, s_r_34__90_, s_r_34__89_, s_r_34__88_, s_r_34__87_, s_r_34__86_, s_r_34__85_, s_r_34__84_, s_r_34__83_, s_r_34__82_, s_r_34__81_, s_r_34__80_, s_r_34__79_, s_r_34__78_, s_r_34__77_, s_r_34__76_, s_r_34__75_, s_r_34__74_, s_r_34__73_, s_r_34__72_, s_r_34__71_, s_r_34__70_, s_r_34__69_, s_r_34__68_, s_r_34__67_, s_r_34__66_, s_r_34__65_, s_r_34__64_, s_r_34__63_, s_r_34__62_, s_r_34__61_, s_r_34__60_, s_r_34__59_, s_r_34__58_, s_r_34__57_, s_r_34__56_, s_r_34__55_, s_r_34__54_, s_r_34__53_, s_r_34__52_, s_r_34__51_, s_r_34__50_, s_r_34__49_, s_r_34__48_, s_r_34__47_, s_r_34__46_, s_r_34__45_, s_r_34__44_, s_r_34__43_, s_r_34__42_, s_r_34__41_, s_r_34__40_, s_r_34__39_, s_r_34__38_, s_r_34__37_, s_r_34__36_, s_r_34__35_, s_r_34__34_, s_r_34__33_, s_r_34__32_, s_r_34__31_, s_r_34__30_, s_r_34__29_, s_r_34__28_, s_r_34__27_, s_r_34__26_, s_r_34__25_, s_r_34__24_, s_r_34__23_, s_r_34__22_, s_r_34__21_, s_r_34__20_, s_r_34__19_, s_r_34__18_, s_r_34__17_, s_r_34__16_, s_r_34__15_, s_r_34__14_, s_r_34__13_, s_r_34__12_, s_r_34__11_, s_r_34__10_, s_r_34__9_, s_r_34__8_, s_r_34__7_, s_r_34__6_, s_r_34__5_, s_r_34__4_, s_r_34__3_, s_r_34__2_, s_r_34__1_, s_r_34__0_ }),
    .c_o(c_r[34]),
    .prod_accum_o({ prod_accum_34__35_, prod_accum_34__34_, prod_accum_34__33_, prod_accum_34__32_, prod_accum_34__31_, prod_accum_34__30_, prod_accum_34__29_, prod_accum_34__28_, prod_accum_34__27_, prod_accum_34__26_, prod_accum_34__25_, prod_accum_34__24_, prod_accum_34__23_, prod_accum_34__22_, prod_accum_34__21_, prod_accum_34__20_, prod_accum_34__19_, prod_accum_34__18_, prod_accum_34__17_, prod_accum_34__16_, prod_accum_34__15_, prod_accum_34__14_, prod_accum_34__13_, prod_accum_34__12_, prod_accum_34__11_, prod_accum_34__10_, prod_accum_34__9_, prod_accum_34__8_, prod_accum_34__7_, prod_accum_34__6_, prod_accum_34__5_, prod_accum_34__4_, prod_accum_34__3_, prod_accum_34__2_, prod_accum_34__1_, prod_accum_34__0_ })
  );


  bsg_mul_array_row_128_35_x
  genblk1_35__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[4479:4352]),
    .b_i(b_r[4479:4352]),
    .s_i({ s_r_34__127_, s_r_34__126_, s_r_34__125_, s_r_34__124_, s_r_34__123_, s_r_34__122_, s_r_34__121_, s_r_34__120_, s_r_34__119_, s_r_34__118_, s_r_34__117_, s_r_34__116_, s_r_34__115_, s_r_34__114_, s_r_34__113_, s_r_34__112_, s_r_34__111_, s_r_34__110_, s_r_34__109_, s_r_34__108_, s_r_34__107_, s_r_34__106_, s_r_34__105_, s_r_34__104_, s_r_34__103_, s_r_34__102_, s_r_34__101_, s_r_34__100_, s_r_34__99_, s_r_34__98_, s_r_34__97_, s_r_34__96_, s_r_34__95_, s_r_34__94_, s_r_34__93_, s_r_34__92_, s_r_34__91_, s_r_34__90_, s_r_34__89_, s_r_34__88_, s_r_34__87_, s_r_34__86_, s_r_34__85_, s_r_34__84_, s_r_34__83_, s_r_34__82_, s_r_34__81_, s_r_34__80_, s_r_34__79_, s_r_34__78_, s_r_34__77_, s_r_34__76_, s_r_34__75_, s_r_34__74_, s_r_34__73_, s_r_34__72_, s_r_34__71_, s_r_34__70_, s_r_34__69_, s_r_34__68_, s_r_34__67_, s_r_34__66_, s_r_34__65_, s_r_34__64_, s_r_34__63_, s_r_34__62_, s_r_34__61_, s_r_34__60_, s_r_34__59_, s_r_34__58_, s_r_34__57_, s_r_34__56_, s_r_34__55_, s_r_34__54_, s_r_34__53_, s_r_34__52_, s_r_34__51_, s_r_34__50_, s_r_34__49_, s_r_34__48_, s_r_34__47_, s_r_34__46_, s_r_34__45_, s_r_34__44_, s_r_34__43_, s_r_34__42_, s_r_34__41_, s_r_34__40_, s_r_34__39_, s_r_34__38_, s_r_34__37_, s_r_34__36_, s_r_34__35_, s_r_34__34_, s_r_34__33_, s_r_34__32_, s_r_34__31_, s_r_34__30_, s_r_34__29_, s_r_34__28_, s_r_34__27_, s_r_34__26_, s_r_34__25_, s_r_34__24_, s_r_34__23_, s_r_34__22_, s_r_34__21_, s_r_34__20_, s_r_34__19_, s_r_34__18_, s_r_34__17_, s_r_34__16_, s_r_34__15_, s_r_34__14_, s_r_34__13_, s_r_34__12_, s_r_34__11_, s_r_34__10_, s_r_34__9_, s_r_34__8_, s_r_34__7_, s_r_34__6_, s_r_34__5_, s_r_34__4_, s_r_34__3_, s_r_34__2_, s_r_34__1_, s_r_34__0_ }),
    .c_i(c_r[34]),
    .prod_accum_i({ prod_accum_34__35_, prod_accum_34__34_, prod_accum_34__33_, prod_accum_34__32_, prod_accum_34__31_, prod_accum_34__30_, prod_accum_34__29_, prod_accum_34__28_, prod_accum_34__27_, prod_accum_34__26_, prod_accum_34__25_, prod_accum_34__24_, prod_accum_34__23_, prod_accum_34__22_, prod_accum_34__21_, prod_accum_34__20_, prod_accum_34__19_, prod_accum_34__18_, prod_accum_34__17_, prod_accum_34__16_, prod_accum_34__15_, prod_accum_34__14_, prod_accum_34__13_, prod_accum_34__12_, prod_accum_34__11_, prod_accum_34__10_, prod_accum_34__9_, prod_accum_34__8_, prod_accum_34__7_, prod_accum_34__6_, prod_accum_34__5_, prod_accum_34__4_, prod_accum_34__3_, prod_accum_34__2_, prod_accum_34__1_, prod_accum_34__0_ }),
    .a_o(a_r[4607:4480]),
    .b_o(b_r[4607:4480]),
    .s_o({ s_r_35__127_, s_r_35__126_, s_r_35__125_, s_r_35__124_, s_r_35__123_, s_r_35__122_, s_r_35__121_, s_r_35__120_, s_r_35__119_, s_r_35__118_, s_r_35__117_, s_r_35__116_, s_r_35__115_, s_r_35__114_, s_r_35__113_, s_r_35__112_, s_r_35__111_, s_r_35__110_, s_r_35__109_, s_r_35__108_, s_r_35__107_, s_r_35__106_, s_r_35__105_, s_r_35__104_, s_r_35__103_, s_r_35__102_, s_r_35__101_, s_r_35__100_, s_r_35__99_, s_r_35__98_, s_r_35__97_, s_r_35__96_, s_r_35__95_, s_r_35__94_, s_r_35__93_, s_r_35__92_, s_r_35__91_, s_r_35__90_, s_r_35__89_, s_r_35__88_, s_r_35__87_, s_r_35__86_, s_r_35__85_, s_r_35__84_, s_r_35__83_, s_r_35__82_, s_r_35__81_, s_r_35__80_, s_r_35__79_, s_r_35__78_, s_r_35__77_, s_r_35__76_, s_r_35__75_, s_r_35__74_, s_r_35__73_, s_r_35__72_, s_r_35__71_, s_r_35__70_, s_r_35__69_, s_r_35__68_, s_r_35__67_, s_r_35__66_, s_r_35__65_, s_r_35__64_, s_r_35__63_, s_r_35__62_, s_r_35__61_, s_r_35__60_, s_r_35__59_, s_r_35__58_, s_r_35__57_, s_r_35__56_, s_r_35__55_, s_r_35__54_, s_r_35__53_, s_r_35__52_, s_r_35__51_, s_r_35__50_, s_r_35__49_, s_r_35__48_, s_r_35__47_, s_r_35__46_, s_r_35__45_, s_r_35__44_, s_r_35__43_, s_r_35__42_, s_r_35__41_, s_r_35__40_, s_r_35__39_, s_r_35__38_, s_r_35__37_, s_r_35__36_, s_r_35__35_, s_r_35__34_, s_r_35__33_, s_r_35__32_, s_r_35__31_, s_r_35__30_, s_r_35__29_, s_r_35__28_, s_r_35__27_, s_r_35__26_, s_r_35__25_, s_r_35__24_, s_r_35__23_, s_r_35__22_, s_r_35__21_, s_r_35__20_, s_r_35__19_, s_r_35__18_, s_r_35__17_, s_r_35__16_, s_r_35__15_, s_r_35__14_, s_r_35__13_, s_r_35__12_, s_r_35__11_, s_r_35__10_, s_r_35__9_, s_r_35__8_, s_r_35__7_, s_r_35__6_, s_r_35__5_, s_r_35__4_, s_r_35__3_, s_r_35__2_, s_r_35__1_, s_r_35__0_ }),
    .c_o(c_r[35]),
    .prod_accum_o({ prod_accum_35__36_, prod_accum_35__35_, prod_accum_35__34_, prod_accum_35__33_, prod_accum_35__32_, prod_accum_35__31_, prod_accum_35__30_, prod_accum_35__29_, prod_accum_35__28_, prod_accum_35__27_, prod_accum_35__26_, prod_accum_35__25_, prod_accum_35__24_, prod_accum_35__23_, prod_accum_35__22_, prod_accum_35__21_, prod_accum_35__20_, prod_accum_35__19_, prod_accum_35__18_, prod_accum_35__17_, prod_accum_35__16_, prod_accum_35__15_, prod_accum_35__14_, prod_accum_35__13_, prod_accum_35__12_, prod_accum_35__11_, prod_accum_35__10_, prod_accum_35__9_, prod_accum_35__8_, prod_accum_35__7_, prod_accum_35__6_, prod_accum_35__5_, prod_accum_35__4_, prod_accum_35__3_, prod_accum_35__2_, prod_accum_35__1_, prod_accum_35__0_ })
  );


  bsg_mul_array_row_128_36_x
  genblk1_36__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[4607:4480]),
    .b_i(b_r[4607:4480]),
    .s_i({ s_r_35__127_, s_r_35__126_, s_r_35__125_, s_r_35__124_, s_r_35__123_, s_r_35__122_, s_r_35__121_, s_r_35__120_, s_r_35__119_, s_r_35__118_, s_r_35__117_, s_r_35__116_, s_r_35__115_, s_r_35__114_, s_r_35__113_, s_r_35__112_, s_r_35__111_, s_r_35__110_, s_r_35__109_, s_r_35__108_, s_r_35__107_, s_r_35__106_, s_r_35__105_, s_r_35__104_, s_r_35__103_, s_r_35__102_, s_r_35__101_, s_r_35__100_, s_r_35__99_, s_r_35__98_, s_r_35__97_, s_r_35__96_, s_r_35__95_, s_r_35__94_, s_r_35__93_, s_r_35__92_, s_r_35__91_, s_r_35__90_, s_r_35__89_, s_r_35__88_, s_r_35__87_, s_r_35__86_, s_r_35__85_, s_r_35__84_, s_r_35__83_, s_r_35__82_, s_r_35__81_, s_r_35__80_, s_r_35__79_, s_r_35__78_, s_r_35__77_, s_r_35__76_, s_r_35__75_, s_r_35__74_, s_r_35__73_, s_r_35__72_, s_r_35__71_, s_r_35__70_, s_r_35__69_, s_r_35__68_, s_r_35__67_, s_r_35__66_, s_r_35__65_, s_r_35__64_, s_r_35__63_, s_r_35__62_, s_r_35__61_, s_r_35__60_, s_r_35__59_, s_r_35__58_, s_r_35__57_, s_r_35__56_, s_r_35__55_, s_r_35__54_, s_r_35__53_, s_r_35__52_, s_r_35__51_, s_r_35__50_, s_r_35__49_, s_r_35__48_, s_r_35__47_, s_r_35__46_, s_r_35__45_, s_r_35__44_, s_r_35__43_, s_r_35__42_, s_r_35__41_, s_r_35__40_, s_r_35__39_, s_r_35__38_, s_r_35__37_, s_r_35__36_, s_r_35__35_, s_r_35__34_, s_r_35__33_, s_r_35__32_, s_r_35__31_, s_r_35__30_, s_r_35__29_, s_r_35__28_, s_r_35__27_, s_r_35__26_, s_r_35__25_, s_r_35__24_, s_r_35__23_, s_r_35__22_, s_r_35__21_, s_r_35__20_, s_r_35__19_, s_r_35__18_, s_r_35__17_, s_r_35__16_, s_r_35__15_, s_r_35__14_, s_r_35__13_, s_r_35__12_, s_r_35__11_, s_r_35__10_, s_r_35__9_, s_r_35__8_, s_r_35__7_, s_r_35__6_, s_r_35__5_, s_r_35__4_, s_r_35__3_, s_r_35__2_, s_r_35__1_, s_r_35__0_ }),
    .c_i(c_r[35]),
    .prod_accum_i({ prod_accum_35__36_, prod_accum_35__35_, prod_accum_35__34_, prod_accum_35__33_, prod_accum_35__32_, prod_accum_35__31_, prod_accum_35__30_, prod_accum_35__29_, prod_accum_35__28_, prod_accum_35__27_, prod_accum_35__26_, prod_accum_35__25_, prod_accum_35__24_, prod_accum_35__23_, prod_accum_35__22_, prod_accum_35__21_, prod_accum_35__20_, prod_accum_35__19_, prod_accum_35__18_, prod_accum_35__17_, prod_accum_35__16_, prod_accum_35__15_, prod_accum_35__14_, prod_accum_35__13_, prod_accum_35__12_, prod_accum_35__11_, prod_accum_35__10_, prod_accum_35__9_, prod_accum_35__8_, prod_accum_35__7_, prod_accum_35__6_, prod_accum_35__5_, prod_accum_35__4_, prod_accum_35__3_, prod_accum_35__2_, prod_accum_35__1_, prod_accum_35__0_ }),
    .a_o(a_r[4735:4608]),
    .b_o(b_r[4735:4608]),
    .s_o({ s_r_36__127_, s_r_36__126_, s_r_36__125_, s_r_36__124_, s_r_36__123_, s_r_36__122_, s_r_36__121_, s_r_36__120_, s_r_36__119_, s_r_36__118_, s_r_36__117_, s_r_36__116_, s_r_36__115_, s_r_36__114_, s_r_36__113_, s_r_36__112_, s_r_36__111_, s_r_36__110_, s_r_36__109_, s_r_36__108_, s_r_36__107_, s_r_36__106_, s_r_36__105_, s_r_36__104_, s_r_36__103_, s_r_36__102_, s_r_36__101_, s_r_36__100_, s_r_36__99_, s_r_36__98_, s_r_36__97_, s_r_36__96_, s_r_36__95_, s_r_36__94_, s_r_36__93_, s_r_36__92_, s_r_36__91_, s_r_36__90_, s_r_36__89_, s_r_36__88_, s_r_36__87_, s_r_36__86_, s_r_36__85_, s_r_36__84_, s_r_36__83_, s_r_36__82_, s_r_36__81_, s_r_36__80_, s_r_36__79_, s_r_36__78_, s_r_36__77_, s_r_36__76_, s_r_36__75_, s_r_36__74_, s_r_36__73_, s_r_36__72_, s_r_36__71_, s_r_36__70_, s_r_36__69_, s_r_36__68_, s_r_36__67_, s_r_36__66_, s_r_36__65_, s_r_36__64_, s_r_36__63_, s_r_36__62_, s_r_36__61_, s_r_36__60_, s_r_36__59_, s_r_36__58_, s_r_36__57_, s_r_36__56_, s_r_36__55_, s_r_36__54_, s_r_36__53_, s_r_36__52_, s_r_36__51_, s_r_36__50_, s_r_36__49_, s_r_36__48_, s_r_36__47_, s_r_36__46_, s_r_36__45_, s_r_36__44_, s_r_36__43_, s_r_36__42_, s_r_36__41_, s_r_36__40_, s_r_36__39_, s_r_36__38_, s_r_36__37_, s_r_36__36_, s_r_36__35_, s_r_36__34_, s_r_36__33_, s_r_36__32_, s_r_36__31_, s_r_36__30_, s_r_36__29_, s_r_36__28_, s_r_36__27_, s_r_36__26_, s_r_36__25_, s_r_36__24_, s_r_36__23_, s_r_36__22_, s_r_36__21_, s_r_36__20_, s_r_36__19_, s_r_36__18_, s_r_36__17_, s_r_36__16_, s_r_36__15_, s_r_36__14_, s_r_36__13_, s_r_36__12_, s_r_36__11_, s_r_36__10_, s_r_36__9_, s_r_36__8_, s_r_36__7_, s_r_36__6_, s_r_36__5_, s_r_36__4_, s_r_36__3_, s_r_36__2_, s_r_36__1_, s_r_36__0_ }),
    .c_o(c_r[36]),
    .prod_accum_o({ prod_accum_36__37_, prod_accum_36__36_, prod_accum_36__35_, prod_accum_36__34_, prod_accum_36__33_, prod_accum_36__32_, prod_accum_36__31_, prod_accum_36__30_, prod_accum_36__29_, prod_accum_36__28_, prod_accum_36__27_, prod_accum_36__26_, prod_accum_36__25_, prod_accum_36__24_, prod_accum_36__23_, prod_accum_36__22_, prod_accum_36__21_, prod_accum_36__20_, prod_accum_36__19_, prod_accum_36__18_, prod_accum_36__17_, prod_accum_36__16_, prod_accum_36__15_, prod_accum_36__14_, prod_accum_36__13_, prod_accum_36__12_, prod_accum_36__11_, prod_accum_36__10_, prod_accum_36__9_, prod_accum_36__8_, prod_accum_36__7_, prod_accum_36__6_, prod_accum_36__5_, prod_accum_36__4_, prod_accum_36__3_, prod_accum_36__2_, prod_accum_36__1_, prod_accum_36__0_ })
  );


  bsg_mul_array_row_128_37_x
  genblk1_37__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[4735:4608]),
    .b_i(b_r[4735:4608]),
    .s_i({ s_r_36__127_, s_r_36__126_, s_r_36__125_, s_r_36__124_, s_r_36__123_, s_r_36__122_, s_r_36__121_, s_r_36__120_, s_r_36__119_, s_r_36__118_, s_r_36__117_, s_r_36__116_, s_r_36__115_, s_r_36__114_, s_r_36__113_, s_r_36__112_, s_r_36__111_, s_r_36__110_, s_r_36__109_, s_r_36__108_, s_r_36__107_, s_r_36__106_, s_r_36__105_, s_r_36__104_, s_r_36__103_, s_r_36__102_, s_r_36__101_, s_r_36__100_, s_r_36__99_, s_r_36__98_, s_r_36__97_, s_r_36__96_, s_r_36__95_, s_r_36__94_, s_r_36__93_, s_r_36__92_, s_r_36__91_, s_r_36__90_, s_r_36__89_, s_r_36__88_, s_r_36__87_, s_r_36__86_, s_r_36__85_, s_r_36__84_, s_r_36__83_, s_r_36__82_, s_r_36__81_, s_r_36__80_, s_r_36__79_, s_r_36__78_, s_r_36__77_, s_r_36__76_, s_r_36__75_, s_r_36__74_, s_r_36__73_, s_r_36__72_, s_r_36__71_, s_r_36__70_, s_r_36__69_, s_r_36__68_, s_r_36__67_, s_r_36__66_, s_r_36__65_, s_r_36__64_, s_r_36__63_, s_r_36__62_, s_r_36__61_, s_r_36__60_, s_r_36__59_, s_r_36__58_, s_r_36__57_, s_r_36__56_, s_r_36__55_, s_r_36__54_, s_r_36__53_, s_r_36__52_, s_r_36__51_, s_r_36__50_, s_r_36__49_, s_r_36__48_, s_r_36__47_, s_r_36__46_, s_r_36__45_, s_r_36__44_, s_r_36__43_, s_r_36__42_, s_r_36__41_, s_r_36__40_, s_r_36__39_, s_r_36__38_, s_r_36__37_, s_r_36__36_, s_r_36__35_, s_r_36__34_, s_r_36__33_, s_r_36__32_, s_r_36__31_, s_r_36__30_, s_r_36__29_, s_r_36__28_, s_r_36__27_, s_r_36__26_, s_r_36__25_, s_r_36__24_, s_r_36__23_, s_r_36__22_, s_r_36__21_, s_r_36__20_, s_r_36__19_, s_r_36__18_, s_r_36__17_, s_r_36__16_, s_r_36__15_, s_r_36__14_, s_r_36__13_, s_r_36__12_, s_r_36__11_, s_r_36__10_, s_r_36__9_, s_r_36__8_, s_r_36__7_, s_r_36__6_, s_r_36__5_, s_r_36__4_, s_r_36__3_, s_r_36__2_, s_r_36__1_, s_r_36__0_ }),
    .c_i(c_r[36]),
    .prod_accum_i({ prod_accum_36__37_, prod_accum_36__36_, prod_accum_36__35_, prod_accum_36__34_, prod_accum_36__33_, prod_accum_36__32_, prod_accum_36__31_, prod_accum_36__30_, prod_accum_36__29_, prod_accum_36__28_, prod_accum_36__27_, prod_accum_36__26_, prod_accum_36__25_, prod_accum_36__24_, prod_accum_36__23_, prod_accum_36__22_, prod_accum_36__21_, prod_accum_36__20_, prod_accum_36__19_, prod_accum_36__18_, prod_accum_36__17_, prod_accum_36__16_, prod_accum_36__15_, prod_accum_36__14_, prod_accum_36__13_, prod_accum_36__12_, prod_accum_36__11_, prod_accum_36__10_, prod_accum_36__9_, prod_accum_36__8_, prod_accum_36__7_, prod_accum_36__6_, prod_accum_36__5_, prod_accum_36__4_, prod_accum_36__3_, prod_accum_36__2_, prod_accum_36__1_, prod_accum_36__0_ }),
    .a_o(a_r[4863:4736]),
    .b_o(b_r[4863:4736]),
    .s_o({ s_r_37__127_, s_r_37__126_, s_r_37__125_, s_r_37__124_, s_r_37__123_, s_r_37__122_, s_r_37__121_, s_r_37__120_, s_r_37__119_, s_r_37__118_, s_r_37__117_, s_r_37__116_, s_r_37__115_, s_r_37__114_, s_r_37__113_, s_r_37__112_, s_r_37__111_, s_r_37__110_, s_r_37__109_, s_r_37__108_, s_r_37__107_, s_r_37__106_, s_r_37__105_, s_r_37__104_, s_r_37__103_, s_r_37__102_, s_r_37__101_, s_r_37__100_, s_r_37__99_, s_r_37__98_, s_r_37__97_, s_r_37__96_, s_r_37__95_, s_r_37__94_, s_r_37__93_, s_r_37__92_, s_r_37__91_, s_r_37__90_, s_r_37__89_, s_r_37__88_, s_r_37__87_, s_r_37__86_, s_r_37__85_, s_r_37__84_, s_r_37__83_, s_r_37__82_, s_r_37__81_, s_r_37__80_, s_r_37__79_, s_r_37__78_, s_r_37__77_, s_r_37__76_, s_r_37__75_, s_r_37__74_, s_r_37__73_, s_r_37__72_, s_r_37__71_, s_r_37__70_, s_r_37__69_, s_r_37__68_, s_r_37__67_, s_r_37__66_, s_r_37__65_, s_r_37__64_, s_r_37__63_, s_r_37__62_, s_r_37__61_, s_r_37__60_, s_r_37__59_, s_r_37__58_, s_r_37__57_, s_r_37__56_, s_r_37__55_, s_r_37__54_, s_r_37__53_, s_r_37__52_, s_r_37__51_, s_r_37__50_, s_r_37__49_, s_r_37__48_, s_r_37__47_, s_r_37__46_, s_r_37__45_, s_r_37__44_, s_r_37__43_, s_r_37__42_, s_r_37__41_, s_r_37__40_, s_r_37__39_, s_r_37__38_, s_r_37__37_, s_r_37__36_, s_r_37__35_, s_r_37__34_, s_r_37__33_, s_r_37__32_, s_r_37__31_, s_r_37__30_, s_r_37__29_, s_r_37__28_, s_r_37__27_, s_r_37__26_, s_r_37__25_, s_r_37__24_, s_r_37__23_, s_r_37__22_, s_r_37__21_, s_r_37__20_, s_r_37__19_, s_r_37__18_, s_r_37__17_, s_r_37__16_, s_r_37__15_, s_r_37__14_, s_r_37__13_, s_r_37__12_, s_r_37__11_, s_r_37__10_, s_r_37__9_, s_r_37__8_, s_r_37__7_, s_r_37__6_, s_r_37__5_, s_r_37__4_, s_r_37__3_, s_r_37__2_, s_r_37__1_, s_r_37__0_ }),
    .c_o(c_r[37]),
    .prod_accum_o({ prod_accum_37__38_, prod_accum_37__37_, prod_accum_37__36_, prod_accum_37__35_, prod_accum_37__34_, prod_accum_37__33_, prod_accum_37__32_, prod_accum_37__31_, prod_accum_37__30_, prod_accum_37__29_, prod_accum_37__28_, prod_accum_37__27_, prod_accum_37__26_, prod_accum_37__25_, prod_accum_37__24_, prod_accum_37__23_, prod_accum_37__22_, prod_accum_37__21_, prod_accum_37__20_, prod_accum_37__19_, prod_accum_37__18_, prod_accum_37__17_, prod_accum_37__16_, prod_accum_37__15_, prod_accum_37__14_, prod_accum_37__13_, prod_accum_37__12_, prod_accum_37__11_, prod_accum_37__10_, prod_accum_37__9_, prod_accum_37__8_, prod_accum_37__7_, prod_accum_37__6_, prod_accum_37__5_, prod_accum_37__4_, prod_accum_37__3_, prod_accum_37__2_, prod_accum_37__1_, prod_accum_37__0_ })
  );


  bsg_mul_array_row_128_38_x
  genblk1_38__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[4863:4736]),
    .b_i(b_r[4863:4736]),
    .s_i({ s_r_37__127_, s_r_37__126_, s_r_37__125_, s_r_37__124_, s_r_37__123_, s_r_37__122_, s_r_37__121_, s_r_37__120_, s_r_37__119_, s_r_37__118_, s_r_37__117_, s_r_37__116_, s_r_37__115_, s_r_37__114_, s_r_37__113_, s_r_37__112_, s_r_37__111_, s_r_37__110_, s_r_37__109_, s_r_37__108_, s_r_37__107_, s_r_37__106_, s_r_37__105_, s_r_37__104_, s_r_37__103_, s_r_37__102_, s_r_37__101_, s_r_37__100_, s_r_37__99_, s_r_37__98_, s_r_37__97_, s_r_37__96_, s_r_37__95_, s_r_37__94_, s_r_37__93_, s_r_37__92_, s_r_37__91_, s_r_37__90_, s_r_37__89_, s_r_37__88_, s_r_37__87_, s_r_37__86_, s_r_37__85_, s_r_37__84_, s_r_37__83_, s_r_37__82_, s_r_37__81_, s_r_37__80_, s_r_37__79_, s_r_37__78_, s_r_37__77_, s_r_37__76_, s_r_37__75_, s_r_37__74_, s_r_37__73_, s_r_37__72_, s_r_37__71_, s_r_37__70_, s_r_37__69_, s_r_37__68_, s_r_37__67_, s_r_37__66_, s_r_37__65_, s_r_37__64_, s_r_37__63_, s_r_37__62_, s_r_37__61_, s_r_37__60_, s_r_37__59_, s_r_37__58_, s_r_37__57_, s_r_37__56_, s_r_37__55_, s_r_37__54_, s_r_37__53_, s_r_37__52_, s_r_37__51_, s_r_37__50_, s_r_37__49_, s_r_37__48_, s_r_37__47_, s_r_37__46_, s_r_37__45_, s_r_37__44_, s_r_37__43_, s_r_37__42_, s_r_37__41_, s_r_37__40_, s_r_37__39_, s_r_37__38_, s_r_37__37_, s_r_37__36_, s_r_37__35_, s_r_37__34_, s_r_37__33_, s_r_37__32_, s_r_37__31_, s_r_37__30_, s_r_37__29_, s_r_37__28_, s_r_37__27_, s_r_37__26_, s_r_37__25_, s_r_37__24_, s_r_37__23_, s_r_37__22_, s_r_37__21_, s_r_37__20_, s_r_37__19_, s_r_37__18_, s_r_37__17_, s_r_37__16_, s_r_37__15_, s_r_37__14_, s_r_37__13_, s_r_37__12_, s_r_37__11_, s_r_37__10_, s_r_37__9_, s_r_37__8_, s_r_37__7_, s_r_37__6_, s_r_37__5_, s_r_37__4_, s_r_37__3_, s_r_37__2_, s_r_37__1_, s_r_37__0_ }),
    .c_i(c_r[37]),
    .prod_accum_i({ prod_accum_37__38_, prod_accum_37__37_, prod_accum_37__36_, prod_accum_37__35_, prod_accum_37__34_, prod_accum_37__33_, prod_accum_37__32_, prod_accum_37__31_, prod_accum_37__30_, prod_accum_37__29_, prod_accum_37__28_, prod_accum_37__27_, prod_accum_37__26_, prod_accum_37__25_, prod_accum_37__24_, prod_accum_37__23_, prod_accum_37__22_, prod_accum_37__21_, prod_accum_37__20_, prod_accum_37__19_, prod_accum_37__18_, prod_accum_37__17_, prod_accum_37__16_, prod_accum_37__15_, prod_accum_37__14_, prod_accum_37__13_, prod_accum_37__12_, prod_accum_37__11_, prod_accum_37__10_, prod_accum_37__9_, prod_accum_37__8_, prod_accum_37__7_, prod_accum_37__6_, prod_accum_37__5_, prod_accum_37__4_, prod_accum_37__3_, prod_accum_37__2_, prod_accum_37__1_, prod_accum_37__0_ }),
    .a_o(a_r[4991:4864]),
    .b_o(b_r[4991:4864]),
    .s_o({ s_r_38__127_, s_r_38__126_, s_r_38__125_, s_r_38__124_, s_r_38__123_, s_r_38__122_, s_r_38__121_, s_r_38__120_, s_r_38__119_, s_r_38__118_, s_r_38__117_, s_r_38__116_, s_r_38__115_, s_r_38__114_, s_r_38__113_, s_r_38__112_, s_r_38__111_, s_r_38__110_, s_r_38__109_, s_r_38__108_, s_r_38__107_, s_r_38__106_, s_r_38__105_, s_r_38__104_, s_r_38__103_, s_r_38__102_, s_r_38__101_, s_r_38__100_, s_r_38__99_, s_r_38__98_, s_r_38__97_, s_r_38__96_, s_r_38__95_, s_r_38__94_, s_r_38__93_, s_r_38__92_, s_r_38__91_, s_r_38__90_, s_r_38__89_, s_r_38__88_, s_r_38__87_, s_r_38__86_, s_r_38__85_, s_r_38__84_, s_r_38__83_, s_r_38__82_, s_r_38__81_, s_r_38__80_, s_r_38__79_, s_r_38__78_, s_r_38__77_, s_r_38__76_, s_r_38__75_, s_r_38__74_, s_r_38__73_, s_r_38__72_, s_r_38__71_, s_r_38__70_, s_r_38__69_, s_r_38__68_, s_r_38__67_, s_r_38__66_, s_r_38__65_, s_r_38__64_, s_r_38__63_, s_r_38__62_, s_r_38__61_, s_r_38__60_, s_r_38__59_, s_r_38__58_, s_r_38__57_, s_r_38__56_, s_r_38__55_, s_r_38__54_, s_r_38__53_, s_r_38__52_, s_r_38__51_, s_r_38__50_, s_r_38__49_, s_r_38__48_, s_r_38__47_, s_r_38__46_, s_r_38__45_, s_r_38__44_, s_r_38__43_, s_r_38__42_, s_r_38__41_, s_r_38__40_, s_r_38__39_, s_r_38__38_, s_r_38__37_, s_r_38__36_, s_r_38__35_, s_r_38__34_, s_r_38__33_, s_r_38__32_, s_r_38__31_, s_r_38__30_, s_r_38__29_, s_r_38__28_, s_r_38__27_, s_r_38__26_, s_r_38__25_, s_r_38__24_, s_r_38__23_, s_r_38__22_, s_r_38__21_, s_r_38__20_, s_r_38__19_, s_r_38__18_, s_r_38__17_, s_r_38__16_, s_r_38__15_, s_r_38__14_, s_r_38__13_, s_r_38__12_, s_r_38__11_, s_r_38__10_, s_r_38__9_, s_r_38__8_, s_r_38__7_, s_r_38__6_, s_r_38__5_, s_r_38__4_, s_r_38__3_, s_r_38__2_, s_r_38__1_, s_r_38__0_ }),
    .c_o(c_r[38]),
    .prod_accum_o({ prod_accum_38__39_, prod_accum_38__38_, prod_accum_38__37_, prod_accum_38__36_, prod_accum_38__35_, prod_accum_38__34_, prod_accum_38__33_, prod_accum_38__32_, prod_accum_38__31_, prod_accum_38__30_, prod_accum_38__29_, prod_accum_38__28_, prod_accum_38__27_, prod_accum_38__26_, prod_accum_38__25_, prod_accum_38__24_, prod_accum_38__23_, prod_accum_38__22_, prod_accum_38__21_, prod_accum_38__20_, prod_accum_38__19_, prod_accum_38__18_, prod_accum_38__17_, prod_accum_38__16_, prod_accum_38__15_, prod_accum_38__14_, prod_accum_38__13_, prod_accum_38__12_, prod_accum_38__11_, prod_accum_38__10_, prod_accum_38__9_, prod_accum_38__8_, prod_accum_38__7_, prod_accum_38__6_, prod_accum_38__5_, prod_accum_38__4_, prod_accum_38__3_, prod_accum_38__2_, prod_accum_38__1_, prod_accum_38__0_ })
  );


  bsg_mul_array_row_128_39_x
  genblk1_39__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[4991:4864]),
    .b_i(b_r[4991:4864]),
    .s_i({ s_r_38__127_, s_r_38__126_, s_r_38__125_, s_r_38__124_, s_r_38__123_, s_r_38__122_, s_r_38__121_, s_r_38__120_, s_r_38__119_, s_r_38__118_, s_r_38__117_, s_r_38__116_, s_r_38__115_, s_r_38__114_, s_r_38__113_, s_r_38__112_, s_r_38__111_, s_r_38__110_, s_r_38__109_, s_r_38__108_, s_r_38__107_, s_r_38__106_, s_r_38__105_, s_r_38__104_, s_r_38__103_, s_r_38__102_, s_r_38__101_, s_r_38__100_, s_r_38__99_, s_r_38__98_, s_r_38__97_, s_r_38__96_, s_r_38__95_, s_r_38__94_, s_r_38__93_, s_r_38__92_, s_r_38__91_, s_r_38__90_, s_r_38__89_, s_r_38__88_, s_r_38__87_, s_r_38__86_, s_r_38__85_, s_r_38__84_, s_r_38__83_, s_r_38__82_, s_r_38__81_, s_r_38__80_, s_r_38__79_, s_r_38__78_, s_r_38__77_, s_r_38__76_, s_r_38__75_, s_r_38__74_, s_r_38__73_, s_r_38__72_, s_r_38__71_, s_r_38__70_, s_r_38__69_, s_r_38__68_, s_r_38__67_, s_r_38__66_, s_r_38__65_, s_r_38__64_, s_r_38__63_, s_r_38__62_, s_r_38__61_, s_r_38__60_, s_r_38__59_, s_r_38__58_, s_r_38__57_, s_r_38__56_, s_r_38__55_, s_r_38__54_, s_r_38__53_, s_r_38__52_, s_r_38__51_, s_r_38__50_, s_r_38__49_, s_r_38__48_, s_r_38__47_, s_r_38__46_, s_r_38__45_, s_r_38__44_, s_r_38__43_, s_r_38__42_, s_r_38__41_, s_r_38__40_, s_r_38__39_, s_r_38__38_, s_r_38__37_, s_r_38__36_, s_r_38__35_, s_r_38__34_, s_r_38__33_, s_r_38__32_, s_r_38__31_, s_r_38__30_, s_r_38__29_, s_r_38__28_, s_r_38__27_, s_r_38__26_, s_r_38__25_, s_r_38__24_, s_r_38__23_, s_r_38__22_, s_r_38__21_, s_r_38__20_, s_r_38__19_, s_r_38__18_, s_r_38__17_, s_r_38__16_, s_r_38__15_, s_r_38__14_, s_r_38__13_, s_r_38__12_, s_r_38__11_, s_r_38__10_, s_r_38__9_, s_r_38__8_, s_r_38__7_, s_r_38__6_, s_r_38__5_, s_r_38__4_, s_r_38__3_, s_r_38__2_, s_r_38__1_, s_r_38__0_ }),
    .c_i(c_r[38]),
    .prod_accum_i({ prod_accum_38__39_, prod_accum_38__38_, prod_accum_38__37_, prod_accum_38__36_, prod_accum_38__35_, prod_accum_38__34_, prod_accum_38__33_, prod_accum_38__32_, prod_accum_38__31_, prod_accum_38__30_, prod_accum_38__29_, prod_accum_38__28_, prod_accum_38__27_, prod_accum_38__26_, prod_accum_38__25_, prod_accum_38__24_, prod_accum_38__23_, prod_accum_38__22_, prod_accum_38__21_, prod_accum_38__20_, prod_accum_38__19_, prod_accum_38__18_, prod_accum_38__17_, prod_accum_38__16_, prod_accum_38__15_, prod_accum_38__14_, prod_accum_38__13_, prod_accum_38__12_, prod_accum_38__11_, prod_accum_38__10_, prod_accum_38__9_, prod_accum_38__8_, prod_accum_38__7_, prod_accum_38__6_, prod_accum_38__5_, prod_accum_38__4_, prod_accum_38__3_, prod_accum_38__2_, prod_accum_38__1_, prod_accum_38__0_ }),
    .a_o(a_r[5119:4992]),
    .b_o(b_r[5119:4992]),
    .s_o({ s_r_39__127_, s_r_39__126_, s_r_39__125_, s_r_39__124_, s_r_39__123_, s_r_39__122_, s_r_39__121_, s_r_39__120_, s_r_39__119_, s_r_39__118_, s_r_39__117_, s_r_39__116_, s_r_39__115_, s_r_39__114_, s_r_39__113_, s_r_39__112_, s_r_39__111_, s_r_39__110_, s_r_39__109_, s_r_39__108_, s_r_39__107_, s_r_39__106_, s_r_39__105_, s_r_39__104_, s_r_39__103_, s_r_39__102_, s_r_39__101_, s_r_39__100_, s_r_39__99_, s_r_39__98_, s_r_39__97_, s_r_39__96_, s_r_39__95_, s_r_39__94_, s_r_39__93_, s_r_39__92_, s_r_39__91_, s_r_39__90_, s_r_39__89_, s_r_39__88_, s_r_39__87_, s_r_39__86_, s_r_39__85_, s_r_39__84_, s_r_39__83_, s_r_39__82_, s_r_39__81_, s_r_39__80_, s_r_39__79_, s_r_39__78_, s_r_39__77_, s_r_39__76_, s_r_39__75_, s_r_39__74_, s_r_39__73_, s_r_39__72_, s_r_39__71_, s_r_39__70_, s_r_39__69_, s_r_39__68_, s_r_39__67_, s_r_39__66_, s_r_39__65_, s_r_39__64_, s_r_39__63_, s_r_39__62_, s_r_39__61_, s_r_39__60_, s_r_39__59_, s_r_39__58_, s_r_39__57_, s_r_39__56_, s_r_39__55_, s_r_39__54_, s_r_39__53_, s_r_39__52_, s_r_39__51_, s_r_39__50_, s_r_39__49_, s_r_39__48_, s_r_39__47_, s_r_39__46_, s_r_39__45_, s_r_39__44_, s_r_39__43_, s_r_39__42_, s_r_39__41_, s_r_39__40_, s_r_39__39_, s_r_39__38_, s_r_39__37_, s_r_39__36_, s_r_39__35_, s_r_39__34_, s_r_39__33_, s_r_39__32_, s_r_39__31_, s_r_39__30_, s_r_39__29_, s_r_39__28_, s_r_39__27_, s_r_39__26_, s_r_39__25_, s_r_39__24_, s_r_39__23_, s_r_39__22_, s_r_39__21_, s_r_39__20_, s_r_39__19_, s_r_39__18_, s_r_39__17_, s_r_39__16_, s_r_39__15_, s_r_39__14_, s_r_39__13_, s_r_39__12_, s_r_39__11_, s_r_39__10_, s_r_39__9_, s_r_39__8_, s_r_39__7_, s_r_39__6_, s_r_39__5_, s_r_39__4_, s_r_39__3_, s_r_39__2_, s_r_39__1_, s_r_39__0_ }),
    .c_o(c_r[39]),
    .prod_accum_o({ prod_accum_39__40_, prod_accum_39__39_, prod_accum_39__38_, prod_accum_39__37_, prod_accum_39__36_, prod_accum_39__35_, prod_accum_39__34_, prod_accum_39__33_, prod_accum_39__32_, prod_accum_39__31_, prod_accum_39__30_, prod_accum_39__29_, prod_accum_39__28_, prod_accum_39__27_, prod_accum_39__26_, prod_accum_39__25_, prod_accum_39__24_, prod_accum_39__23_, prod_accum_39__22_, prod_accum_39__21_, prod_accum_39__20_, prod_accum_39__19_, prod_accum_39__18_, prod_accum_39__17_, prod_accum_39__16_, prod_accum_39__15_, prod_accum_39__14_, prod_accum_39__13_, prod_accum_39__12_, prod_accum_39__11_, prod_accum_39__10_, prod_accum_39__9_, prod_accum_39__8_, prod_accum_39__7_, prod_accum_39__6_, prod_accum_39__5_, prod_accum_39__4_, prod_accum_39__3_, prod_accum_39__2_, prod_accum_39__1_, prod_accum_39__0_ })
  );


  bsg_mul_array_row_128_40_x
  genblk1_40__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[5119:4992]),
    .b_i(b_r[5119:4992]),
    .s_i({ s_r_39__127_, s_r_39__126_, s_r_39__125_, s_r_39__124_, s_r_39__123_, s_r_39__122_, s_r_39__121_, s_r_39__120_, s_r_39__119_, s_r_39__118_, s_r_39__117_, s_r_39__116_, s_r_39__115_, s_r_39__114_, s_r_39__113_, s_r_39__112_, s_r_39__111_, s_r_39__110_, s_r_39__109_, s_r_39__108_, s_r_39__107_, s_r_39__106_, s_r_39__105_, s_r_39__104_, s_r_39__103_, s_r_39__102_, s_r_39__101_, s_r_39__100_, s_r_39__99_, s_r_39__98_, s_r_39__97_, s_r_39__96_, s_r_39__95_, s_r_39__94_, s_r_39__93_, s_r_39__92_, s_r_39__91_, s_r_39__90_, s_r_39__89_, s_r_39__88_, s_r_39__87_, s_r_39__86_, s_r_39__85_, s_r_39__84_, s_r_39__83_, s_r_39__82_, s_r_39__81_, s_r_39__80_, s_r_39__79_, s_r_39__78_, s_r_39__77_, s_r_39__76_, s_r_39__75_, s_r_39__74_, s_r_39__73_, s_r_39__72_, s_r_39__71_, s_r_39__70_, s_r_39__69_, s_r_39__68_, s_r_39__67_, s_r_39__66_, s_r_39__65_, s_r_39__64_, s_r_39__63_, s_r_39__62_, s_r_39__61_, s_r_39__60_, s_r_39__59_, s_r_39__58_, s_r_39__57_, s_r_39__56_, s_r_39__55_, s_r_39__54_, s_r_39__53_, s_r_39__52_, s_r_39__51_, s_r_39__50_, s_r_39__49_, s_r_39__48_, s_r_39__47_, s_r_39__46_, s_r_39__45_, s_r_39__44_, s_r_39__43_, s_r_39__42_, s_r_39__41_, s_r_39__40_, s_r_39__39_, s_r_39__38_, s_r_39__37_, s_r_39__36_, s_r_39__35_, s_r_39__34_, s_r_39__33_, s_r_39__32_, s_r_39__31_, s_r_39__30_, s_r_39__29_, s_r_39__28_, s_r_39__27_, s_r_39__26_, s_r_39__25_, s_r_39__24_, s_r_39__23_, s_r_39__22_, s_r_39__21_, s_r_39__20_, s_r_39__19_, s_r_39__18_, s_r_39__17_, s_r_39__16_, s_r_39__15_, s_r_39__14_, s_r_39__13_, s_r_39__12_, s_r_39__11_, s_r_39__10_, s_r_39__9_, s_r_39__8_, s_r_39__7_, s_r_39__6_, s_r_39__5_, s_r_39__4_, s_r_39__3_, s_r_39__2_, s_r_39__1_, s_r_39__0_ }),
    .c_i(c_r[39]),
    .prod_accum_i({ prod_accum_39__40_, prod_accum_39__39_, prod_accum_39__38_, prod_accum_39__37_, prod_accum_39__36_, prod_accum_39__35_, prod_accum_39__34_, prod_accum_39__33_, prod_accum_39__32_, prod_accum_39__31_, prod_accum_39__30_, prod_accum_39__29_, prod_accum_39__28_, prod_accum_39__27_, prod_accum_39__26_, prod_accum_39__25_, prod_accum_39__24_, prod_accum_39__23_, prod_accum_39__22_, prod_accum_39__21_, prod_accum_39__20_, prod_accum_39__19_, prod_accum_39__18_, prod_accum_39__17_, prod_accum_39__16_, prod_accum_39__15_, prod_accum_39__14_, prod_accum_39__13_, prod_accum_39__12_, prod_accum_39__11_, prod_accum_39__10_, prod_accum_39__9_, prod_accum_39__8_, prod_accum_39__7_, prod_accum_39__6_, prod_accum_39__5_, prod_accum_39__4_, prod_accum_39__3_, prod_accum_39__2_, prod_accum_39__1_, prod_accum_39__0_ }),
    .a_o(a_r[5247:5120]),
    .b_o(b_r[5247:5120]),
    .s_o({ s_r_40__127_, s_r_40__126_, s_r_40__125_, s_r_40__124_, s_r_40__123_, s_r_40__122_, s_r_40__121_, s_r_40__120_, s_r_40__119_, s_r_40__118_, s_r_40__117_, s_r_40__116_, s_r_40__115_, s_r_40__114_, s_r_40__113_, s_r_40__112_, s_r_40__111_, s_r_40__110_, s_r_40__109_, s_r_40__108_, s_r_40__107_, s_r_40__106_, s_r_40__105_, s_r_40__104_, s_r_40__103_, s_r_40__102_, s_r_40__101_, s_r_40__100_, s_r_40__99_, s_r_40__98_, s_r_40__97_, s_r_40__96_, s_r_40__95_, s_r_40__94_, s_r_40__93_, s_r_40__92_, s_r_40__91_, s_r_40__90_, s_r_40__89_, s_r_40__88_, s_r_40__87_, s_r_40__86_, s_r_40__85_, s_r_40__84_, s_r_40__83_, s_r_40__82_, s_r_40__81_, s_r_40__80_, s_r_40__79_, s_r_40__78_, s_r_40__77_, s_r_40__76_, s_r_40__75_, s_r_40__74_, s_r_40__73_, s_r_40__72_, s_r_40__71_, s_r_40__70_, s_r_40__69_, s_r_40__68_, s_r_40__67_, s_r_40__66_, s_r_40__65_, s_r_40__64_, s_r_40__63_, s_r_40__62_, s_r_40__61_, s_r_40__60_, s_r_40__59_, s_r_40__58_, s_r_40__57_, s_r_40__56_, s_r_40__55_, s_r_40__54_, s_r_40__53_, s_r_40__52_, s_r_40__51_, s_r_40__50_, s_r_40__49_, s_r_40__48_, s_r_40__47_, s_r_40__46_, s_r_40__45_, s_r_40__44_, s_r_40__43_, s_r_40__42_, s_r_40__41_, s_r_40__40_, s_r_40__39_, s_r_40__38_, s_r_40__37_, s_r_40__36_, s_r_40__35_, s_r_40__34_, s_r_40__33_, s_r_40__32_, s_r_40__31_, s_r_40__30_, s_r_40__29_, s_r_40__28_, s_r_40__27_, s_r_40__26_, s_r_40__25_, s_r_40__24_, s_r_40__23_, s_r_40__22_, s_r_40__21_, s_r_40__20_, s_r_40__19_, s_r_40__18_, s_r_40__17_, s_r_40__16_, s_r_40__15_, s_r_40__14_, s_r_40__13_, s_r_40__12_, s_r_40__11_, s_r_40__10_, s_r_40__9_, s_r_40__8_, s_r_40__7_, s_r_40__6_, s_r_40__5_, s_r_40__4_, s_r_40__3_, s_r_40__2_, s_r_40__1_, s_r_40__0_ }),
    .c_o(c_r[40]),
    .prod_accum_o({ prod_accum_40__41_, prod_accum_40__40_, prod_accum_40__39_, prod_accum_40__38_, prod_accum_40__37_, prod_accum_40__36_, prod_accum_40__35_, prod_accum_40__34_, prod_accum_40__33_, prod_accum_40__32_, prod_accum_40__31_, prod_accum_40__30_, prod_accum_40__29_, prod_accum_40__28_, prod_accum_40__27_, prod_accum_40__26_, prod_accum_40__25_, prod_accum_40__24_, prod_accum_40__23_, prod_accum_40__22_, prod_accum_40__21_, prod_accum_40__20_, prod_accum_40__19_, prod_accum_40__18_, prod_accum_40__17_, prod_accum_40__16_, prod_accum_40__15_, prod_accum_40__14_, prod_accum_40__13_, prod_accum_40__12_, prod_accum_40__11_, prod_accum_40__10_, prod_accum_40__9_, prod_accum_40__8_, prod_accum_40__7_, prod_accum_40__6_, prod_accum_40__5_, prod_accum_40__4_, prod_accum_40__3_, prod_accum_40__2_, prod_accum_40__1_, prod_accum_40__0_ })
  );


  bsg_mul_array_row_128_41_x
  genblk1_41__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[5247:5120]),
    .b_i(b_r[5247:5120]),
    .s_i({ s_r_40__127_, s_r_40__126_, s_r_40__125_, s_r_40__124_, s_r_40__123_, s_r_40__122_, s_r_40__121_, s_r_40__120_, s_r_40__119_, s_r_40__118_, s_r_40__117_, s_r_40__116_, s_r_40__115_, s_r_40__114_, s_r_40__113_, s_r_40__112_, s_r_40__111_, s_r_40__110_, s_r_40__109_, s_r_40__108_, s_r_40__107_, s_r_40__106_, s_r_40__105_, s_r_40__104_, s_r_40__103_, s_r_40__102_, s_r_40__101_, s_r_40__100_, s_r_40__99_, s_r_40__98_, s_r_40__97_, s_r_40__96_, s_r_40__95_, s_r_40__94_, s_r_40__93_, s_r_40__92_, s_r_40__91_, s_r_40__90_, s_r_40__89_, s_r_40__88_, s_r_40__87_, s_r_40__86_, s_r_40__85_, s_r_40__84_, s_r_40__83_, s_r_40__82_, s_r_40__81_, s_r_40__80_, s_r_40__79_, s_r_40__78_, s_r_40__77_, s_r_40__76_, s_r_40__75_, s_r_40__74_, s_r_40__73_, s_r_40__72_, s_r_40__71_, s_r_40__70_, s_r_40__69_, s_r_40__68_, s_r_40__67_, s_r_40__66_, s_r_40__65_, s_r_40__64_, s_r_40__63_, s_r_40__62_, s_r_40__61_, s_r_40__60_, s_r_40__59_, s_r_40__58_, s_r_40__57_, s_r_40__56_, s_r_40__55_, s_r_40__54_, s_r_40__53_, s_r_40__52_, s_r_40__51_, s_r_40__50_, s_r_40__49_, s_r_40__48_, s_r_40__47_, s_r_40__46_, s_r_40__45_, s_r_40__44_, s_r_40__43_, s_r_40__42_, s_r_40__41_, s_r_40__40_, s_r_40__39_, s_r_40__38_, s_r_40__37_, s_r_40__36_, s_r_40__35_, s_r_40__34_, s_r_40__33_, s_r_40__32_, s_r_40__31_, s_r_40__30_, s_r_40__29_, s_r_40__28_, s_r_40__27_, s_r_40__26_, s_r_40__25_, s_r_40__24_, s_r_40__23_, s_r_40__22_, s_r_40__21_, s_r_40__20_, s_r_40__19_, s_r_40__18_, s_r_40__17_, s_r_40__16_, s_r_40__15_, s_r_40__14_, s_r_40__13_, s_r_40__12_, s_r_40__11_, s_r_40__10_, s_r_40__9_, s_r_40__8_, s_r_40__7_, s_r_40__6_, s_r_40__5_, s_r_40__4_, s_r_40__3_, s_r_40__2_, s_r_40__1_, s_r_40__0_ }),
    .c_i(c_r[40]),
    .prod_accum_i({ prod_accum_40__41_, prod_accum_40__40_, prod_accum_40__39_, prod_accum_40__38_, prod_accum_40__37_, prod_accum_40__36_, prod_accum_40__35_, prod_accum_40__34_, prod_accum_40__33_, prod_accum_40__32_, prod_accum_40__31_, prod_accum_40__30_, prod_accum_40__29_, prod_accum_40__28_, prod_accum_40__27_, prod_accum_40__26_, prod_accum_40__25_, prod_accum_40__24_, prod_accum_40__23_, prod_accum_40__22_, prod_accum_40__21_, prod_accum_40__20_, prod_accum_40__19_, prod_accum_40__18_, prod_accum_40__17_, prod_accum_40__16_, prod_accum_40__15_, prod_accum_40__14_, prod_accum_40__13_, prod_accum_40__12_, prod_accum_40__11_, prod_accum_40__10_, prod_accum_40__9_, prod_accum_40__8_, prod_accum_40__7_, prod_accum_40__6_, prod_accum_40__5_, prod_accum_40__4_, prod_accum_40__3_, prod_accum_40__2_, prod_accum_40__1_, prod_accum_40__0_ }),
    .a_o(a_r[5375:5248]),
    .b_o(b_r[5375:5248]),
    .s_o({ s_r_41__127_, s_r_41__126_, s_r_41__125_, s_r_41__124_, s_r_41__123_, s_r_41__122_, s_r_41__121_, s_r_41__120_, s_r_41__119_, s_r_41__118_, s_r_41__117_, s_r_41__116_, s_r_41__115_, s_r_41__114_, s_r_41__113_, s_r_41__112_, s_r_41__111_, s_r_41__110_, s_r_41__109_, s_r_41__108_, s_r_41__107_, s_r_41__106_, s_r_41__105_, s_r_41__104_, s_r_41__103_, s_r_41__102_, s_r_41__101_, s_r_41__100_, s_r_41__99_, s_r_41__98_, s_r_41__97_, s_r_41__96_, s_r_41__95_, s_r_41__94_, s_r_41__93_, s_r_41__92_, s_r_41__91_, s_r_41__90_, s_r_41__89_, s_r_41__88_, s_r_41__87_, s_r_41__86_, s_r_41__85_, s_r_41__84_, s_r_41__83_, s_r_41__82_, s_r_41__81_, s_r_41__80_, s_r_41__79_, s_r_41__78_, s_r_41__77_, s_r_41__76_, s_r_41__75_, s_r_41__74_, s_r_41__73_, s_r_41__72_, s_r_41__71_, s_r_41__70_, s_r_41__69_, s_r_41__68_, s_r_41__67_, s_r_41__66_, s_r_41__65_, s_r_41__64_, s_r_41__63_, s_r_41__62_, s_r_41__61_, s_r_41__60_, s_r_41__59_, s_r_41__58_, s_r_41__57_, s_r_41__56_, s_r_41__55_, s_r_41__54_, s_r_41__53_, s_r_41__52_, s_r_41__51_, s_r_41__50_, s_r_41__49_, s_r_41__48_, s_r_41__47_, s_r_41__46_, s_r_41__45_, s_r_41__44_, s_r_41__43_, s_r_41__42_, s_r_41__41_, s_r_41__40_, s_r_41__39_, s_r_41__38_, s_r_41__37_, s_r_41__36_, s_r_41__35_, s_r_41__34_, s_r_41__33_, s_r_41__32_, s_r_41__31_, s_r_41__30_, s_r_41__29_, s_r_41__28_, s_r_41__27_, s_r_41__26_, s_r_41__25_, s_r_41__24_, s_r_41__23_, s_r_41__22_, s_r_41__21_, s_r_41__20_, s_r_41__19_, s_r_41__18_, s_r_41__17_, s_r_41__16_, s_r_41__15_, s_r_41__14_, s_r_41__13_, s_r_41__12_, s_r_41__11_, s_r_41__10_, s_r_41__9_, s_r_41__8_, s_r_41__7_, s_r_41__6_, s_r_41__5_, s_r_41__4_, s_r_41__3_, s_r_41__2_, s_r_41__1_, s_r_41__0_ }),
    .c_o(c_r[41]),
    .prod_accum_o({ prod_accum_41__42_, prod_accum_41__41_, prod_accum_41__40_, prod_accum_41__39_, prod_accum_41__38_, prod_accum_41__37_, prod_accum_41__36_, prod_accum_41__35_, prod_accum_41__34_, prod_accum_41__33_, prod_accum_41__32_, prod_accum_41__31_, prod_accum_41__30_, prod_accum_41__29_, prod_accum_41__28_, prod_accum_41__27_, prod_accum_41__26_, prod_accum_41__25_, prod_accum_41__24_, prod_accum_41__23_, prod_accum_41__22_, prod_accum_41__21_, prod_accum_41__20_, prod_accum_41__19_, prod_accum_41__18_, prod_accum_41__17_, prod_accum_41__16_, prod_accum_41__15_, prod_accum_41__14_, prod_accum_41__13_, prod_accum_41__12_, prod_accum_41__11_, prod_accum_41__10_, prod_accum_41__9_, prod_accum_41__8_, prod_accum_41__7_, prod_accum_41__6_, prod_accum_41__5_, prod_accum_41__4_, prod_accum_41__3_, prod_accum_41__2_, prod_accum_41__1_, prod_accum_41__0_ })
  );


  bsg_mul_array_row_128_42_x
  genblk1_42__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[5375:5248]),
    .b_i(b_r[5375:5248]),
    .s_i({ s_r_41__127_, s_r_41__126_, s_r_41__125_, s_r_41__124_, s_r_41__123_, s_r_41__122_, s_r_41__121_, s_r_41__120_, s_r_41__119_, s_r_41__118_, s_r_41__117_, s_r_41__116_, s_r_41__115_, s_r_41__114_, s_r_41__113_, s_r_41__112_, s_r_41__111_, s_r_41__110_, s_r_41__109_, s_r_41__108_, s_r_41__107_, s_r_41__106_, s_r_41__105_, s_r_41__104_, s_r_41__103_, s_r_41__102_, s_r_41__101_, s_r_41__100_, s_r_41__99_, s_r_41__98_, s_r_41__97_, s_r_41__96_, s_r_41__95_, s_r_41__94_, s_r_41__93_, s_r_41__92_, s_r_41__91_, s_r_41__90_, s_r_41__89_, s_r_41__88_, s_r_41__87_, s_r_41__86_, s_r_41__85_, s_r_41__84_, s_r_41__83_, s_r_41__82_, s_r_41__81_, s_r_41__80_, s_r_41__79_, s_r_41__78_, s_r_41__77_, s_r_41__76_, s_r_41__75_, s_r_41__74_, s_r_41__73_, s_r_41__72_, s_r_41__71_, s_r_41__70_, s_r_41__69_, s_r_41__68_, s_r_41__67_, s_r_41__66_, s_r_41__65_, s_r_41__64_, s_r_41__63_, s_r_41__62_, s_r_41__61_, s_r_41__60_, s_r_41__59_, s_r_41__58_, s_r_41__57_, s_r_41__56_, s_r_41__55_, s_r_41__54_, s_r_41__53_, s_r_41__52_, s_r_41__51_, s_r_41__50_, s_r_41__49_, s_r_41__48_, s_r_41__47_, s_r_41__46_, s_r_41__45_, s_r_41__44_, s_r_41__43_, s_r_41__42_, s_r_41__41_, s_r_41__40_, s_r_41__39_, s_r_41__38_, s_r_41__37_, s_r_41__36_, s_r_41__35_, s_r_41__34_, s_r_41__33_, s_r_41__32_, s_r_41__31_, s_r_41__30_, s_r_41__29_, s_r_41__28_, s_r_41__27_, s_r_41__26_, s_r_41__25_, s_r_41__24_, s_r_41__23_, s_r_41__22_, s_r_41__21_, s_r_41__20_, s_r_41__19_, s_r_41__18_, s_r_41__17_, s_r_41__16_, s_r_41__15_, s_r_41__14_, s_r_41__13_, s_r_41__12_, s_r_41__11_, s_r_41__10_, s_r_41__9_, s_r_41__8_, s_r_41__7_, s_r_41__6_, s_r_41__5_, s_r_41__4_, s_r_41__3_, s_r_41__2_, s_r_41__1_, s_r_41__0_ }),
    .c_i(c_r[41]),
    .prod_accum_i({ prod_accum_41__42_, prod_accum_41__41_, prod_accum_41__40_, prod_accum_41__39_, prod_accum_41__38_, prod_accum_41__37_, prod_accum_41__36_, prod_accum_41__35_, prod_accum_41__34_, prod_accum_41__33_, prod_accum_41__32_, prod_accum_41__31_, prod_accum_41__30_, prod_accum_41__29_, prod_accum_41__28_, prod_accum_41__27_, prod_accum_41__26_, prod_accum_41__25_, prod_accum_41__24_, prod_accum_41__23_, prod_accum_41__22_, prod_accum_41__21_, prod_accum_41__20_, prod_accum_41__19_, prod_accum_41__18_, prod_accum_41__17_, prod_accum_41__16_, prod_accum_41__15_, prod_accum_41__14_, prod_accum_41__13_, prod_accum_41__12_, prod_accum_41__11_, prod_accum_41__10_, prod_accum_41__9_, prod_accum_41__8_, prod_accum_41__7_, prod_accum_41__6_, prod_accum_41__5_, prod_accum_41__4_, prod_accum_41__3_, prod_accum_41__2_, prod_accum_41__1_, prod_accum_41__0_ }),
    .a_o(a_r[5503:5376]),
    .b_o(b_r[5503:5376]),
    .s_o({ s_r_42__127_, s_r_42__126_, s_r_42__125_, s_r_42__124_, s_r_42__123_, s_r_42__122_, s_r_42__121_, s_r_42__120_, s_r_42__119_, s_r_42__118_, s_r_42__117_, s_r_42__116_, s_r_42__115_, s_r_42__114_, s_r_42__113_, s_r_42__112_, s_r_42__111_, s_r_42__110_, s_r_42__109_, s_r_42__108_, s_r_42__107_, s_r_42__106_, s_r_42__105_, s_r_42__104_, s_r_42__103_, s_r_42__102_, s_r_42__101_, s_r_42__100_, s_r_42__99_, s_r_42__98_, s_r_42__97_, s_r_42__96_, s_r_42__95_, s_r_42__94_, s_r_42__93_, s_r_42__92_, s_r_42__91_, s_r_42__90_, s_r_42__89_, s_r_42__88_, s_r_42__87_, s_r_42__86_, s_r_42__85_, s_r_42__84_, s_r_42__83_, s_r_42__82_, s_r_42__81_, s_r_42__80_, s_r_42__79_, s_r_42__78_, s_r_42__77_, s_r_42__76_, s_r_42__75_, s_r_42__74_, s_r_42__73_, s_r_42__72_, s_r_42__71_, s_r_42__70_, s_r_42__69_, s_r_42__68_, s_r_42__67_, s_r_42__66_, s_r_42__65_, s_r_42__64_, s_r_42__63_, s_r_42__62_, s_r_42__61_, s_r_42__60_, s_r_42__59_, s_r_42__58_, s_r_42__57_, s_r_42__56_, s_r_42__55_, s_r_42__54_, s_r_42__53_, s_r_42__52_, s_r_42__51_, s_r_42__50_, s_r_42__49_, s_r_42__48_, s_r_42__47_, s_r_42__46_, s_r_42__45_, s_r_42__44_, s_r_42__43_, s_r_42__42_, s_r_42__41_, s_r_42__40_, s_r_42__39_, s_r_42__38_, s_r_42__37_, s_r_42__36_, s_r_42__35_, s_r_42__34_, s_r_42__33_, s_r_42__32_, s_r_42__31_, s_r_42__30_, s_r_42__29_, s_r_42__28_, s_r_42__27_, s_r_42__26_, s_r_42__25_, s_r_42__24_, s_r_42__23_, s_r_42__22_, s_r_42__21_, s_r_42__20_, s_r_42__19_, s_r_42__18_, s_r_42__17_, s_r_42__16_, s_r_42__15_, s_r_42__14_, s_r_42__13_, s_r_42__12_, s_r_42__11_, s_r_42__10_, s_r_42__9_, s_r_42__8_, s_r_42__7_, s_r_42__6_, s_r_42__5_, s_r_42__4_, s_r_42__3_, s_r_42__2_, s_r_42__1_, s_r_42__0_ }),
    .c_o(c_r[42]),
    .prod_accum_o({ prod_accum_42__43_, prod_accum_42__42_, prod_accum_42__41_, prod_accum_42__40_, prod_accum_42__39_, prod_accum_42__38_, prod_accum_42__37_, prod_accum_42__36_, prod_accum_42__35_, prod_accum_42__34_, prod_accum_42__33_, prod_accum_42__32_, prod_accum_42__31_, prod_accum_42__30_, prod_accum_42__29_, prod_accum_42__28_, prod_accum_42__27_, prod_accum_42__26_, prod_accum_42__25_, prod_accum_42__24_, prod_accum_42__23_, prod_accum_42__22_, prod_accum_42__21_, prod_accum_42__20_, prod_accum_42__19_, prod_accum_42__18_, prod_accum_42__17_, prod_accum_42__16_, prod_accum_42__15_, prod_accum_42__14_, prod_accum_42__13_, prod_accum_42__12_, prod_accum_42__11_, prod_accum_42__10_, prod_accum_42__9_, prod_accum_42__8_, prod_accum_42__7_, prod_accum_42__6_, prod_accum_42__5_, prod_accum_42__4_, prod_accum_42__3_, prod_accum_42__2_, prod_accum_42__1_, prod_accum_42__0_ })
  );


  bsg_mul_array_row_128_43_x
  genblk1_43__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[5503:5376]),
    .b_i(b_r[5503:5376]),
    .s_i({ s_r_42__127_, s_r_42__126_, s_r_42__125_, s_r_42__124_, s_r_42__123_, s_r_42__122_, s_r_42__121_, s_r_42__120_, s_r_42__119_, s_r_42__118_, s_r_42__117_, s_r_42__116_, s_r_42__115_, s_r_42__114_, s_r_42__113_, s_r_42__112_, s_r_42__111_, s_r_42__110_, s_r_42__109_, s_r_42__108_, s_r_42__107_, s_r_42__106_, s_r_42__105_, s_r_42__104_, s_r_42__103_, s_r_42__102_, s_r_42__101_, s_r_42__100_, s_r_42__99_, s_r_42__98_, s_r_42__97_, s_r_42__96_, s_r_42__95_, s_r_42__94_, s_r_42__93_, s_r_42__92_, s_r_42__91_, s_r_42__90_, s_r_42__89_, s_r_42__88_, s_r_42__87_, s_r_42__86_, s_r_42__85_, s_r_42__84_, s_r_42__83_, s_r_42__82_, s_r_42__81_, s_r_42__80_, s_r_42__79_, s_r_42__78_, s_r_42__77_, s_r_42__76_, s_r_42__75_, s_r_42__74_, s_r_42__73_, s_r_42__72_, s_r_42__71_, s_r_42__70_, s_r_42__69_, s_r_42__68_, s_r_42__67_, s_r_42__66_, s_r_42__65_, s_r_42__64_, s_r_42__63_, s_r_42__62_, s_r_42__61_, s_r_42__60_, s_r_42__59_, s_r_42__58_, s_r_42__57_, s_r_42__56_, s_r_42__55_, s_r_42__54_, s_r_42__53_, s_r_42__52_, s_r_42__51_, s_r_42__50_, s_r_42__49_, s_r_42__48_, s_r_42__47_, s_r_42__46_, s_r_42__45_, s_r_42__44_, s_r_42__43_, s_r_42__42_, s_r_42__41_, s_r_42__40_, s_r_42__39_, s_r_42__38_, s_r_42__37_, s_r_42__36_, s_r_42__35_, s_r_42__34_, s_r_42__33_, s_r_42__32_, s_r_42__31_, s_r_42__30_, s_r_42__29_, s_r_42__28_, s_r_42__27_, s_r_42__26_, s_r_42__25_, s_r_42__24_, s_r_42__23_, s_r_42__22_, s_r_42__21_, s_r_42__20_, s_r_42__19_, s_r_42__18_, s_r_42__17_, s_r_42__16_, s_r_42__15_, s_r_42__14_, s_r_42__13_, s_r_42__12_, s_r_42__11_, s_r_42__10_, s_r_42__9_, s_r_42__8_, s_r_42__7_, s_r_42__6_, s_r_42__5_, s_r_42__4_, s_r_42__3_, s_r_42__2_, s_r_42__1_, s_r_42__0_ }),
    .c_i(c_r[42]),
    .prod_accum_i({ prod_accum_42__43_, prod_accum_42__42_, prod_accum_42__41_, prod_accum_42__40_, prod_accum_42__39_, prod_accum_42__38_, prod_accum_42__37_, prod_accum_42__36_, prod_accum_42__35_, prod_accum_42__34_, prod_accum_42__33_, prod_accum_42__32_, prod_accum_42__31_, prod_accum_42__30_, prod_accum_42__29_, prod_accum_42__28_, prod_accum_42__27_, prod_accum_42__26_, prod_accum_42__25_, prod_accum_42__24_, prod_accum_42__23_, prod_accum_42__22_, prod_accum_42__21_, prod_accum_42__20_, prod_accum_42__19_, prod_accum_42__18_, prod_accum_42__17_, prod_accum_42__16_, prod_accum_42__15_, prod_accum_42__14_, prod_accum_42__13_, prod_accum_42__12_, prod_accum_42__11_, prod_accum_42__10_, prod_accum_42__9_, prod_accum_42__8_, prod_accum_42__7_, prod_accum_42__6_, prod_accum_42__5_, prod_accum_42__4_, prod_accum_42__3_, prod_accum_42__2_, prod_accum_42__1_, prod_accum_42__0_ }),
    .a_o(a_r[5631:5504]),
    .b_o(b_r[5631:5504]),
    .s_o({ s_r_43__127_, s_r_43__126_, s_r_43__125_, s_r_43__124_, s_r_43__123_, s_r_43__122_, s_r_43__121_, s_r_43__120_, s_r_43__119_, s_r_43__118_, s_r_43__117_, s_r_43__116_, s_r_43__115_, s_r_43__114_, s_r_43__113_, s_r_43__112_, s_r_43__111_, s_r_43__110_, s_r_43__109_, s_r_43__108_, s_r_43__107_, s_r_43__106_, s_r_43__105_, s_r_43__104_, s_r_43__103_, s_r_43__102_, s_r_43__101_, s_r_43__100_, s_r_43__99_, s_r_43__98_, s_r_43__97_, s_r_43__96_, s_r_43__95_, s_r_43__94_, s_r_43__93_, s_r_43__92_, s_r_43__91_, s_r_43__90_, s_r_43__89_, s_r_43__88_, s_r_43__87_, s_r_43__86_, s_r_43__85_, s_r_43__84_, s_r_43__83_, s_r_43__82_, s_r_43__81_, s_r_43__80_, s_r_43__79_, s_r_43__78_, s_r_43__77_, s_r_43__76_, s_r_43__75_, s_r_43__74_, s_r_43__73_, s_r_43__72_, s_r_43__71_, s_r_43__70_, s_r_43__69_, s_r_43__68_, s_r_43__67_, s_r_43__66_, s_r_43__65_, s_r_43__64_, s_r_43__63_, s_r_43__62_, s_r_43__61_, s_r_43__60_, s_r_43__59_, s_r_43__58_, s_r_43__57_, s_r_43__56_, s_r_43__55_, s_r_43__54_, s_r_43__53_, s_r_43__52_, s_r_43__51_, s_r_43__50_, s_r_43__49_, s_r_43__48_, s_r_43__47_, s_r_43__46_, s_r_43__45_, s_r_43__44_, s_r_43__43_, s_r_43__42_, s_r_43__41_, s_r_43__40_, s_r_43__39_, s_r_43__38_, s_r_43__37_, s_r_43__36_, s_r_43__35_, s_r_43__34_, s_r_43__33_, s_r_43__32_, s_r_43__31_, s_r_43__30_, s_r_43__29_, s_r_43__28_, s_r_43__27_, s_r_43__26_, s_r_43__25_, s_r_43__24_, s_r_43__23_, s_r_43__22_, s_r_43__21_, s_r_43__20_, s_r_43__19_, s_r_43__18_, s_r_43__17_, s_r_43__16_, s_r_43__15_, s_r_43__14_, s_r_43__13_, s_r_43__12_, s_r_43__11_, s_r_43__10_, s_r_43__9_, s_r_43__8_, s_r_43__7_, s_r_43__6_, s_r_43__5_, s_r_43__4_, s_r_43__3_, s_r_43__2_, s_r_43__1_, s_r_43__0_ }),
    .c_o(c_r[43]),
    .prod_accum_o({ prod_accum_43__44_, prod_accum_43__43_, prod_accum_43__42_, prod_accum_43__41_, prod_accum_43__40_, prod_accum_43__39_, prod_accum_43__38_, prod_accum_43__37_, prod_accum_43__36_, prod_accum_43__35_, prod_accum_43__34_, prod_accum_43__33_, prod_accum_43__32_, prod_accum_43__31_, prod_accum_43__30_, prod_accum_43__29_, prod_accum_43__28_, prod_accum_43__27_, prod_accum_43__26_, prod_accum_43__25_, prod_accum_43__24_, prod_accum_43__23_, prod_accum_43__22_, prod_accum_43__21_, prod_accum_43__20_, prod_accum_43__19_, prod_accum_43__18_, prod_accum_43__17_, prod_accum_43__16_, prod_accum_43__15_, prod_accum_43__14_, prod_accum_43__13_, prod_accum_43__12_, prod_accum_43__11_, prod_accum_43__10_, prod_accum_43__9_, prod_accum_43__8_, prod_accum_43__7_, prod_accum_43__6_, prod_accum_43__5_, prod_accum_43__4_, prod_accum_43__3_, prod_accum_43__2_, prod_accum_43__1_, prod_accum_43__0_ })
  );


  bsg_mul_array_row_128_44_x
  genblk1_44__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[5631:5504]),
    .b_i(b_r[5631:5504]),
    .s_i({ s_r_43__127_, s_r_43__126_, s_r_43__125_, s_r_43__124_, s_r_43__123_, s_r_43__122_, s_r_43__121_, s_r_43__120_, s_r_43__119_, s_r_43__118_, s_r_43__117_, s_r_43__116_, s_r_43__115_, s_r_43__114_, s_r_43__113_, s_r_43__112_, s_r_43__111_, s_r_43__110_, s_r_43__109_, s_r_43__108_, s_r_43__107_, s_r_43__106_, s_r_43__105_, s_r_43__104_, s_r_43__103_, s_r_43__102_, s_r_43__101_, s_r_43__100_, s_r_43__99_, s_r_43__98_, s_r_43__97_, s_r_43__96_, s_r_43__95_, s_r_43__94_, s_r_43__93_, s_r_43__92_, s_r_43__91_, s_r_43__90_, s_r_43__89_, s_r_43__88_, s_r_43__87_, s_r_43__86_, s_r_43__85_, s_r_43__84_, s_r_43__83_, s_r_43__82_, s_r_43__81_, s_r_43__80_, s_r_43__79_, s_r_43__78_, s_r_43__77_, s_r_43__76_, s_r_43__75_, s_r_43__74_, s_r_43__73_, s_r_43__72_, s_r_43__71_, s_r_43__70_, s_r_43__69_, s_r_43__68_, s_r_43__67_, s_r_43__66_, s_r_43__65_, s_r_43__64_, s_r_43__63_, s_r_43__62_, s_r_43__61_, s_r_43__60_, s_r_43__59_, s_r_43__58_, s_r_43__57_, s_r_43__56_, s_r_43__55_, s_r_43__54_, s_r_43__53_, s_r_43__52_, s_r_43__51_, s_r_43__50_, s_r_43__49_, s_r_43__48_, s_r_43__47_, s_r_43__46_, s_r_43__45_, s_r_43__44_, s_r_43__43_, s_r_43__42_, s_r_43__41_, s_r_43__40_, s_r_43__39_, s_r_43__38_, s_r_43__37_, s_r_43__36_, s_r_43__35_, s_r_43__34_, s_r_43__33_, s_r_43__32_, s_r_43__31_, s_r_43__30_, s_r_43__29_, s_r_43__28_, s_r_43__27_, s_r_43__26_, s_r_43__25_, s_r_43__24_, s_r_43__23_, s_r_43__22_, s_r_43__21_, s_r_43__20_, s_r_43__19_, s_r_43__18_, s_r_43__17_, s_r_43__16_, s_r_43__15_, s_r_43__14_, s_r_43__13_, s_r_43__12_, s_r_43__11_, s_r_43__10_, s_r_43__9_, s_r_43__8_, s_r_43__7_, s_r_43__6_, s_r_43__5_, s_r_43__4_, s_r_43__3_, s_r_43__2_, s_r_43__1_, s_r_43__0_ }),
    .c_i(c_r[43]),
    .prod_accum_i({ prod_accum_43__44_, prod_accum_43__43_, prod_accum_43__42_, prod_accum_43__41_, prod_accum_43__40_, prod_accum_43__39_, prod_accum_43__38_, prod_accum_43__37_, prod_accum_43__36_, prod_accum_43__35_, prod_accum_43__34_, prod_accum_43__33_, prod_accum_43__32_, prod_accum_43__31_, prod_accum_43__30_, prod_accum_43__29_, prod_accum_43__28_, prod_accum_43__27_, prod_accum_43__26_, prod_accum_43__25_, prod_accum_43__24_, prod_accum_43__23_, prod_accum_43__22_, prod_accum_43__21_, prod_accum_43__20_, prod_accum_43__19_, prod_accum_43__18_, prod_accum_43__17_, prod_accum_43__16_, prod_accum_43__15_, prod_accum_43__14_, prod_accum_43__13_, prod_accum_43__12_, prod_accum_43__11_, prod_accum_43__10_, prod_accum_43__9_, prod_accum_43__8_, prod_accum_43__7_, prod_accum_43__6_, prod_accum_43__5_, prod_accum_43__4_, prod_accum_43__3_, prod_accum_43__2_, prod_accum_43__1_, prod_accum_43__0_ }),
    .a_o(a_r[5759:5632]),
    .b_o(b_r[5759:5632]),
    .s_o({ s_r_44__127_, s_r_44__126_, s_r_44__125_, s_r_44__124_, s_r_44__123_, s_r_44__122_, s_r_44__121_, s_r_44__120_, s_r_44__119_, s_r_44__118_, s_r_44__117_, s_r_44__116_, s_r_44__115_, s_r_44__114_, s_r_44__113_, s_r_44__112_, s_r_44__111_, s_r_44__110_, s_r_44__109_, s_r_44__108_, s_r_44__107_, s_r_44__106_, s_r_44__105_, s_r_44__104_, s_r_44__103_, s_r_44__102_, s_r_44__101_, s_r_44__100_, s_r_44__99_, s_r_44__98_, s_r_44__97_, s_r_44__96_, s_r_44__95_, s_r_44__94_, s_r_44__93_, s_r_44__92_, s_r_44__91_, s_r_44__90_, s_r_44__89_, s_r_44__88_, s_r_44__87_, s_r_44__86_, s_r_44__85_, s_r_44__84_, s_r_44__83_, s_r_44__82_, s_r_44__81_, s_r_44__80_, s_r_44__79_, s_r_44__78_, s_r_44__77_, s_r_44__76_, s_r_44__75_, s_r_44__74_, s_r_44__73_, s_r_44__72_, s_r_44__71_, s_r_44__70_, s_r_44__69_, s_r_44__68_, s_r_44__67_, s_r_44__66_, s_r_44__65_, s_r_44__64_, s_r_44__63_, s_r_44__62_, s_r_44__61_, s_r_44__60_, s_r_44__59_, s_r_44__58_, s_r_44__57_, s_r_44__56_, s_r_44__55_, s_r_44__54_, s_r_44__53_, s_r_44__52_, s_r_44__51_, s_r_44__50_, s_r_44__49_, s_r_44__48_, s_r_44__47_, s_r_44__46_, s_r_44__45_, s_r_44__44_, s_r_44__43_, s_r_44__42_, s_r_44__41_, s_r_44__40_, s_r_44__39_, s_r_44__38_, s_r_44__37_, s_r_44__36_, s_r_44__35_, s_r_44__34_, s_r_44__33_, s_r_44__32_, s_r_44__31_, s_r_44__30_, s_r_44__29_, s_r_44__28_, s_r_44__27_, s_r_44__26_, s_r_44__25_, s_r_44__24_, s_r_44__23_, s_r_44__22_, s_r_44__21_, s_r_44__20_, s_r_44__19_, s_r_44__18_, s_r_44__17_, s_r_44__16_, s_r_44__15_, s_r_44__14_, s_r_44__13_, s_r_44__12_, s_r_44__11_, s_r_44__10_, s_r_44__9_, s_r_44__8_, s_r_44__7_, s_r_44__6_, s_r_44__5_, s_r_44__4_, s_r_44__3_, s_r_44__2_, s_r_44__1_, s_r_44__0_ }),
    .c_o(c_r[44]),
    .prod_accum_o({ prod_accum_44__45_, prod_accum_44__44_, prod_accum_44__43_, prod_accum_44__42_, prod_accum_44__41_, prod_accum_44__40_, prod_accum_44__39_, prod_accum_44__38_, prod_accum_44__37_, prod_accum_44__36_, prod_accum_44__35_, prod_accum_44__34_, prod_accum_44__33_, prod_accum_44__32_, prod_accum_44__31_, prod_accum_44__30_, prod_accum_44__29_, prod_accum_44__28_, prod_accum_44__27_, prod_accum_44__26_, prod_accum_44__25_, prod_accum_44__24_, prod_accum_44__23_, prod_accum_44__22_, prod_accum_44__21_, prod_accum_44__20_, prod_accum_44__19_, prod_accum_44__18_, prod_accum_44__17_, prod_accum_44__16_, prod_accum_44__15_, prod_accum_44__14_, prod_accum_44__13_, prod_accum_44__12_, prod_accum_44__11_, prod_accum_44__10_, prod_accum_44__9_, prod_accum_44__8_, prod_accum_44__7_, prod_accum_44__6_, prod_accum_44__5_, prod_accum_44__4_, prod_accum_44__3_, prod_accum_44__2_, prod_accum_44__1_, prod_accum_44__0_ })
  );


  bsg_mul_array_row_128_45_x
  genblk1_45__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[5759:5632]),
    .b_i(b_r[5759:5632]),
    .s_i({ s_r_44__127_, s_r_44__126_, s_r_44__125_, s_r_44__124_, s_r_44__123_, s_r_44__122_, s_r_44__121_, s_r_44__120_, s_r_44__119_, s_r_44__118_, s_r_44__117_, s_r_44__116_, s_r_44__115_, s_r_44__114_, s_r_44__113_, s_r_44__112_, s_r_44__111_, s_r_44__110_, s_r_44__109_, s_r_44__108_, s_r_44__107_, s_r_44__106_, s_r_44__105_, s_r_44__104_, s_r_44__103_, s_r_44__102_, s_r_44__101_, s_r_44__100_, s_r_44__99_, s_r_44__98_, s_r_44__97_, s_r_44__96_, s_r_44__95_, s_r_44__94_, s_r_44__93_, s_r_44__92_, s_r_44__91_, s_r_44__90_, s_r_44__89_, s_r_44__88_, s_r_44__87_, s_r_44__86_, s_r_44__85_, s_r_44__84_, s_r_44__83_, s_r_44__82_, s_r_44__81_, s_r_44__80_, s_r_44__79_, s_r_44__78_, s_r_44__77_, s_r_44__76_, s_r_44__75_, s_r_44__74_, s_r_44__73_, s_r_44__72_, s_r_44__71_, s_r_44__70_, s_r_44__69_, s_r_44__68_, s_r_44__67_, s_r_44__66_, s_r_44__65_, s_r_44__64_, s_r_44__63_, s_r_44__62_, s_r_44__61_, s_r_44__60_, s_r_44__59_, s_r_44__58_, s_r_44__57_, s_r_44__56_, s_r_44__55_, s_r_44__54_, s_r_44__53_, s_r_44__52_, s_r_44__51_, s_r_44__50_, s_r_44__49_, s_r_44__48_, s_r_44__47_, s_r_44__46_, s_r_44__45_, s_r_44__44_, s_r_44__43_, s_r_44__42_, s_r_44__41_, s_r_44__40_, s_r_44__39_, s_r_44__38_, s_r_44__37_, s_r_44__36_, s_r_44__35_, s_r_44__34_, s_r_44__33_, s_r_44__32_, s_r_44__31_, s_r_44__30_, s_r_44__29_, s_r_44__28_, s_r_44__27_, s_r_44__26_, s_r_44__25_, s_r_44__24_, s_r_44__23_, s_r_44__22_, s_r_44__21_, s_r_44__20_, s_r_44__19_, s_r_44__18_, s_r_44__17_, s_r_44__16_, s_r_44__15_, s_r_44__14_, s_r_44__13_, s_r_44__12_, s_r_44__11_, s_r_44__10_, s_r_44__9_, s_r_44__8_, s_r_44__7_, s_r_44__6_, s_r_44__5_, s_r_44__4_, s_r_44__3_, s_r_44__2_, s_r_44__1_, s_r_44__0_ }),
    .c_i(c_r[44]),
    .prod_accum_i({ prod_accum_44__45_, prod_accum_44__44_, prod_accum_44__43_, prod_accum_44__42_, prod_accum_44__41_, prod_accum_44__40_, prod_accum_44__39_, prod_accum_44__38_, prod_accum_44__37_, prod_accum_44__36_, prod_accum_44__35_, prod_accum_44__34_, prod_accum_44__33_, prod_accum_44__32_, prod_accum_44__31_, prod_accum_44__30_, prod_accum_44__29_, prod_accum_44__28_, prod_accum_44__27_, prod_accum_44__26_, prod_accum_44__25_, prod_accum_44__24_, prod_accum_44__23_, prod_accum_44__22_, prod_accum_44__21_, prod_accum_44__20_, prod_accum_44__19_, prod_accum_44__18_, prod_accum_44__17_, prod_accum_44__16_, prod_accum_44__15_, prod_accum_44__14_, prod_accum_44__13_, prod_accum_44__12_, prod_accum_44__11_, prod_accum_44__10_, prod_accum_44__9_, prod_accum_44__8_, prod_accum_44__7_, prod_accum_44__6_, prod_accum_44__5_, prod_accum_44__4_, prod_accum_44__3_, prod_accum_44__2_, prod_accum_44__1_, prod_accum_44__0_ }),
    .a_o(a_r[5887:5760]),
    .b_o(b_r[5887:5760]),
    .s_o({ s_r_45__127_, s_r_45__126_, s_r_45__125_, s_r_45__124_, s_r_45__123_, s_r_45__122_, s_r_45__121_, s_r_45__120_, s_r_45__119_, s_r_45__118_, s_r_45__117_, s_r_45__116_, s_r_45__115_, s_r_45__114_, s_r_45__113_, s_r_45__112_, s_r_45__111_, s_r_45__110_, s_r_45__109_, s_r_45__108_, s_r_45__107_, s_r_45__106_, s_r_45__105_, s_r_45__104_, s_r_45__103_, s_r_45__102_, s_r_45__101_, s_r_45__100_, s_r_45__99_, s_r_45__98_, s_r_45__97_, s_r_45__96_, s_r_45__95_, s_r_45__94_, s_r_45__93_, s_r_45__92_, s_r_45__91_, s_r_45__90_, s_r_45__89_, s_r_45__88_, s_r_45__87_, s_r_45__86_, s_r_45__85_, s_r_45__84_, s_r_45__83_, s_r_45__82_, s_r_45__81_, s_r_45__80_, s_r_45__79_, s_r_45__78_, s_r_45__77_, s_r_45__76_, s_r_45__75_, s_r_45__74_, s_r_45__73_, s_r_45__72_, s_r_45__71_, s_r_45__70_, s_r_45__69_, s_r_45__68_, s_r_45__67_, s_r_45__66_, s_r_45__65_, s_r_45__64_, s_r_45__63_, s_r_45__62_, s_r_45__61_, s_r_45__60_, s_r_45__59_, s_r_45__58_, s_r_45__57_, s_r_45__56_, s_r_45__55_, s_r_45__54_, s_r_45__53_, s_r_45__52_, s_r_45__51_, s_r_45__50_, s_r_45__49_, s_r_45__48_, s_r_45__47_, s_r_45__46_, s_r_45__45_, s_r_45__44_, s_r_45__43_, s_r_45__42_, s_r_45__41_, s_r_45__40_, s_r_45__39_, s_r_45__38_, s_r_45__37_, s_r_45__36_, s_r_45__35_, s_r_45__34_, s_r_45__33_, s_r_45__32_, s_r_45__31_, s_r_45__30_, s_r_45__29_, s_r_45__28_, s_r_45__27_, s_r_45__26_, s_r_45__25_, s_r_45__24_, s_r_45__23_, s_r_45__22_, s_r_45__21_, s_r_45__20_, s_r_45__19_, s_r_45__18_, s_r_45__17_, s_r_45__16_, s_r_45__15_, s_r_45__14_, s_r_45__13_, s_r_45__12_, s_r_45__11_, s_r_45__10_, s_r_45__9_, s_r_45__8_, s_r_45__7_, s_r_45__6_, s_r_45__5_, s_r_45__4_, s_r_45__3_, s_r_45__2_, s_r_45__1_, s_r_45__0_ }),
    .c_o(c_r[45]),
    .prod_accum_o({ prod_accum_45__46_, prod_accum_45__45_, prod_accum_45__44_, prod_accum_45__43_, prod_accum_45__42_, prod_accum_45__41_, prod_accum_45__40_, prod_accum_45__39_, prod_accum_45__38_, prod_accum_45__37_, prod_accum_45__36_, prod_accum_45__35_, prod_accum_45__34_, prod_accum_45__33_, prod_accum_45__32_, prod_accum_45__31_, prod_accum_45__30_, prod_accum_45__29_, prod_accum_45__28_, prod_accum_45__27_, prod_accum_45__26_, prod_accum_45__25_, prod_accum_45__24_, prod_accum_45__23_, prod_accum_45__22_, prod_accum_45__21_, prod_accum_45__20_, prod_accum_45__19_, prod_accum_45__18_, prod_accum_45__17_, prod_accum_45__16_, prod_accum_45__15_, prod_accum_45__14_, prod_accum_45__13_, prod_accum_45__12_, prod_accum_45__11_, prod_accum_45__10_, prod_accum_45__9_, prod_accum_45__8_, prod_accum_45__7_, prod_accum_45__6_, prod_accum_45__5_, prod_accum_45__4_, prod_accum_45__3_, prod_accum_45__2_, prod_accum_45__1_, prod_accum_45__0_ })
  );


  bsg_mul_array_row_128_46_x
  genblk1_46__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[5887:5760]),
    .b_i(b_r[5887:5760]),
    .s_i({ s_r_45__127_, s_r_45__126_, s_r_45__125_, s_r_45__124_, s_r_45__123_, s_r_45__122_, s_r_45__121_, s_r_45__120_, s_r_45__119_, s_r_45__118_, s_r_45__117_, s_r_45__116_, s_r_45__115_, s_r_45__114_, s_r_45__113_, s_r_45__112_, s_r_45__111_, s_r_45__110_, s_r_45__109_, s_r_45__108_, s_r_45__107_, s_r_45__106_, s_r_45__105_, s_r_45__104_, s_r_45__103_, s_r_45__102_, s_r_45__101_, s_r_45__100_, s_r_45__99_, s_r_45__98_, s_r_45__97_, s_r_45__96_, s_r_45__95_, s_r_45__94_, s_r_45__93_, s_r_45__92_, s_r_45__91_, s_r_45__90_, s_r_45__89_, s_r_45__88_, s_r_45__87_, s_r_45__86_, s_r_45__85_, s_r_45__84_, s_r_45__83_, s_r_45__82_, s_r_45__81_, s_r_45__80_, s_r_45__79_, s_r_45__78_, s_r_45__77_, s_r_45__76_, s_r_45__75_, s_r_45__74_, s_r_45__73_, s_r_45__72_, s_r_45__71_, s_r_45__70_, s_r_45__69_, s_r_45__68_, s_r_45__67_, s_r_45__66_, s_r_45__65_, s_r_45__64_, s_r_45__63_, s_r_45__62_, s_r_45__61_, s_r_45__60_, s_r_45__59_, s_r_45__58_, s_r_45__57_, s_r_45__56_, s_r_45__55_, s_r_45__54_, s_r_45__53_, s_r_45__52_, s_r_45__51_, s_r_45__50_, s_r_45__49_, s_r_45__48_, s_r_45__47_, s_r_45__46_, s_r_45__45_, s_r_45__44_, s_r_45__43_, s_r_45__42_, s_r_45__41_, s_r_45__40_, s_r_45__39_, s_r_45__38_, s_r_45__37_, s_r_45__36_, s_r_45__35_, s_r_45__34_, s_r_45__33_, s_r_45__32_, s_r_45__31_, s_r_45__30_, s_r_45__29_, s_r_45__28_, s_r_45__27_, s_r_45__26_, s_r_45__25_, s_r_45__24_, s_r_45__23_, s_r_45__22_, s_r_45__21_, s_r_45__20_, s_r_45__19_, s_r_45__18_, s_r_45__17_, s_r_45__16_, s_r_45__15_, s_r_45__14_, s_r_45__13_, s_r_45__12_, s_r_45__11_, s_r_45__10_, s_r_45__9_, s_r_45__8_, s_r_45__7_, s_r_45__6_, s_r_45__5_, s_r_45__4_, s_r_45__3_, s_r_45__2_, s_r_45__1_, s_r_45__0_ }),
    .c_i(c_r[45]),
    .prod_accum_i({ prod_accum_45__46_, prod_accum_45__45_, prod_accum_45__44_, prod_accum_45__43_, prod_accum_45__42_, prod_accum_45__41_, prod_accum_45__40_, prod_accum_45__39_, prod_accum_45__38_, prod_accum_45__37_, prod_accum_45__36_, prod_accum_45__35_, prod_accum_45__34_, prod_accum_45__33_, prod_accum_45__32_, prod_accum_45__31_, prod_accum_45__30_, prod_accum_45__29_, prod_accum_45__28_, prod_accum_45__27_, prod_accum_45__26_, prod_accum_45__25_, prod_accum_45__24_, prod_accum_45__23_, prod_accum_45__22_, prod_accum_45__21_, prod_accum_45__20_, prod_accum_45__19_, prod_accum_45__18_, prod_accum_45__17_, prod_accum_45__16_, prod_accum_45__15_, prod_accum_45__14_, prod_accum_45__13_, prod_accum_45__12_, prod_accum_45__11_, prod_accum_45__10_, prod_accum_45__9_, prod_accum_45__8_, prod_accum_45__7_, prod_accum_45__6_, prod_accum_45__5_, prod_accum_45__4_, prod_accum_45__3_, prod_accum_45__2_, prod_accum_45__1_, prod_accum_45__0_ }),
    .a_o(a_r[6015:5888]),
    .b_o(b_r[6015:5888]),
    .s_o({ s_r_46__127_, s_r_46__126_, s_r_46__125_, s_r_46__124_, s_r_46__123_, s_r_46__122_, s_r_46__121_, s_r_46__120_, s_r_46__119_, s_r_46__118_, s_r_46__117_, s_r_46__116_, s_r_46__115_, s_r_46__114_, s_r_46__113_, s_r_46__112_, s_r_46__111_, s_r_46__110_, s_r_46__109_, s_r_46__108_, s_r_46__107_, s_r_46__106_, s_r_46__105_, s_r_46__104_, s_r_46__103_, s_r_46__102_, s_r_46__101_, s_r_46__100_, s_r_46__99_, s_r_46__98_, s_r_46__97_, s_r_46__96_, s_r_46__95_, s_r_46__94_, s_r_46__93_, s_r_46__92_, s_r_46__91_, s_r_46__90_, s_r_46__89_, s_r_46__88_, s_r_46__87_, s_r_46__86_, s_r_46__85_, s_r_46__84_, s_r_46__83_, s_r_46__82_, s_r_46__81_, s_r_46__80_, s_r_46__79_, s_r_46__78_, s_r_46__77_, s_r_46__76_, s_r_46__75_, s_r_46__74_, s_r_46__73_, s_r_46__72_, s_r_46__71_, s_r_46__70_, s_r_46__69_, s_r_46__68_, s_r_46__67_, s_r_46__66_, s_r_46__65_, s_r_46__64_, s_r_46__63_, s_r_46__62_, s_r_46__61_, s_r_46__60_, s_r_46__59_, s_r_46__58_, s_r_46__57_, s_r_46__56_, s_r_46__55_, s_r_46__54_, s_r_46__53_, s_r_46__52_, s_r_46__51_, s_r_46__50_, s_r_46__49_, s_r_46__48_, s_r_46__47_, s_r_46__46_, s_r_46__45_, s_r_46__44_, s_r_46__43_, s_r_46__42_, s_r_46__41_, s_r_46__40_, s_r_46__39_, s_r_46__38_, s_r_46__37_, s_r_46__36_, s_r_46__35_, s_r_46__34_, s_r_46__33_, s_r_46__32_, s_r_46__31_, s_r_46__30_, s_r_46__29_, s_r_46__28_, s_r_46__27_, s_r_46__26_, s_r_46__25_, s_r_46__24_, s_r_46__23_, s_r_46__22_, s_r_46__21_, s_r_46__20_, s_r_46__19_, s_r_46__18_, s_r_46__17_, s_r_46__16_, s_r_46__15_, s_r_46__14_, s_r_46__13_, s_r_46__12_, s_r_46__11_, s_r_46__10_, s_r_46__9_, s_r_46__8_, s_r_46__7_, s_r_46__6_, s_r_46__5_, s_r_46__4_, s_r_46__3_, s_r_46__2_, s_r_46__1_, s_r_46__0_ }),
    .c_o(c_r[46]),
    .prod_accum_o({ prod_accum_46__47_, prod_accum_46__46_, prod_accum_46__45_, prod_accum_46__44_, prod_accum_46__43_, prod_accum_46__42_, prod_accum_46__41_, prod_accum_46__40_, prod_accum_46__39_, prod_accum_46__38_, prod_accum_46__37_, prod_accum_46__36_, prod_accum_46__35_, prod_accum_46__34_, prod_accum_46__33_, prod_accum_46__32_, prod_accum_46__31_, prod_accum_46__30_, prod_accum_46__29_, prod_accum_46__28_, prod_accum_46__27_, prod_accum_46__26_, prod_accum_46__25_, prod_accum_46__24_, prod_accum_46__23_, prod_accum_46__22_, prod_accum_46__21_, prod_accum_46__20_, prod_accum_46__19_, prod_accum_46__18_, prod_accum_46__17_, prod_accum_46__16_, prod_accum_46__15_, prod_accum_46__14_, prod_accum_46__13_, prod_accum_46__12_, prod_accum_46__11_, prod_accum_46__10_, prod_accum_46__9_, prod_accum_46__8_, prod_accum_46__7_, prod_accum_46__6_, prod_accum_46__5_, prod_accum_46__4_, prod_accum_46__3_, prod_accum_46__2_, prod_accum_46__1_, prod_accum_46__0_ })
  );


  bsg_mul_array_row_128_47_x
  genblk1_47__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[6015:5888]),
    .b_i(b_r[6015:5888]),
    .s_i({ s_r_46__127_, s_r_46__126_, s_r_46__125_, s_r_46__124_, s_r_46__123_, s_r_46__122_, s_r_46__121_, s_r_46__120_, s_r_46__119_, s_r_46__118_, s_r_46__117_, s_r_46__116_, s_r_46__115_, s_r_46__114_, s_r_46__113_, s_r_46__112_, s_r_46__111_, s_r_46__110_, s_r_46__109_, s_r_46__108_, s_r_46__107_, s_r_46__106_, s_r_46__105_, s_r_46__104_, s_r_46__103_, s_r_46__102_, s_r_46__101_, s_r_46__100_, s_r_46__99_, s_r_46__98_, s_r_46__97_, s_r_46__96_, s_r_46__95_, s_r_46__94_, s_r_46__93_, s_r_46__92_, s_r_46__91_, s_r_46__90_, s_r_46__89_, s_r_46__88_, s_r_46__87_, s_r_46__86_, s_r_46__85_, s_r_46__84_, s_r_46__83_, s_r_46__82_, s_r_46__81_, s_r_46__80_, s_r_46__79_, s_r_46__78_, s_r_46__77_, s_r_46__76_, s_r_46__75_, s_r_46__74_, s_r_46__73_, s_r_46__72_, s_r_46__71_, s_r_46__70_, s_r_46__69_, s_r_46__68_, s_r_46__67_, s_r_46__66_, s_r_46__65_, s_r_46__64_, s_r_46__63_, s_r_46__62_, s_r_46__61_, s_r_46__60_, s_r_46__59_, s_r_46__58_, s_r_46__57_, s_r_46__56_, s_r_46__55_, s_r_46__54_, s_r_46__53_, s_r_46__52_, s_r_46__51_, s_r_46__50_, s_r_46__49_, s_r_46__48_, s_r_46__47_, s_r_46__46_, s_r_46__45_, s_r_46__44_, s_r_46__43_, s_r_46__42_, s_r_46__41_, s_r_46__40_, s_r_46__39_, s_r_46__38_, s_r_46__37_, s_r_46__36_, s_r_46__35_, s_r_46__34_, s_r_46__33_, s_r_46__32_, s_r_46__31_, s_r_46__30_, s_r_46__29_, s_r_46__28_, s_r_46__27_, s_r_46__26_, s_r_46__25_, s_r_46__24_, s_r_46__23_, s_r_46__22_, s_r_46__21_, s_r_46__20_, s_r_46__19_, s_r_46__18_, s_r_46__17_, s_r_46__16_, s_r_46__15_, s_r_46__14_, s_r_46__13_, s_r_46__12_, s_r_46__11_, s_r_46__10_, s_r_46__9_, s_r_46__8_, s_r_46__7_, s_r_46__6_, s_r_46__5_, s_r_46__4_, s_r_46__3_, s_r_46__2_, s_r_46__1_, s_r_46__0_ }),
    .c_i(c_r[46]),
    .prod_accum_i({ prod_accum_46__47_, prod_accum_46__46_, prod_accum_46__45_, prod_accum_46__44_, prod_accum_46__43_, prod_accum_46__42_, prod_accum_46__41_, prod_accum_46__40_, prod_accum_46__39_, prod_accum_46__38_, prod_accum_46__37_, prod_accum_46__36_, prod_accum_46__35_, prod_accum_46__34_, prod_accum_46__33_, prod_accum_46__32_, prod_accum_46__31_, prod_accum_46__30_, prod_accum_46__29_, prod_accum_46__28_, prod_accum_46__27_, prod_accum_46__26_, prod_accum_46__25_, prod_accum_46__24_, prod_accum_46__23_, prod_accum_46__22_, prod_accum_46__21_, prod_accum_46__20_, prod_accum_46__19_, prod_accum_46__18_, prod_accum_46__17_, prod_accum_46__16_, prod_accum_46__15_, prod_accum_46__14_, prod_accum_46__13_, prod_accum_46__12_, prod_accum_46__11_, prod_accum_46__10_, prod_accum_46__9_, prod_accum_46__8_, prod_accum_46__7_, prod_accum_46__6_, prod_accum_46__5_, prod_accum_46__4_, prod_accum_46__3_, prod_accum_46__2_, prod_accum_46__1_, prod_accum_46__0_ }),
    .a_o(a_r[6143:6016]),
    .b_o(b_r[6143:6016]),
    .s_o({ s_r_47__127_, s_r_47__126_, s_r_47__125_, s_r_47__124_, s_r_47__123_, s_r_47__122_, s_r_47__121_, s_r_47__120_, s_r_47__119_, s_r_47__118_, s_r_47__117_, s_r_47__116_, s_r_47__115_, s_r_47__114_, s_r_47__113_, s_r_47__112_, s_r_47__111_, s_r_47__110_, s_r_47__109_, s_r_47__108_, s_r_47__107_, s_r_47__106_, s_r_47__105_, s_r_47__104_, s_r_47__103_, s_r_47__102_, s_r_47__101_, s_r_47__100_, s_r_47__99_, s_r_47__98_, s_r_47__97_, s_r_47__96_, s_r_47__95_, s_r_47__94_, s_r_47__93_, s_r_47__92_, s_r_47__91_, s_r_47__90_, s_r_47__89_, s_r_47__88_, s_r_47__87_, s_r_47__86_, s_r_47__85_, s_r_47__84_, s_r_47__83_, s_r_47__82_, s_r_47__81_, s_r_47__80_, s_r_47__79_, s_r_47__78_, s_r_47__77_, s_r_47__76_, s_r_47__75_, s_r_47__74_, s_r_47__73_, s_r_47__72_, s_r_47__71_, s_r_47__70_, s_r_47__69_, s_r_47__68_, s_r_47__67_, s_r_47__66_, s_r_47__65_, s_r_47__64_, s_r_47__63_, s_r_47__62_, s_r_47__61_, s_r_47__60_, s_r_47__59_, s_r_47__58_, s_r_47__57_, s_r_47__56_, s_r_47__55_, s_r_47__54_, s_r_47__53_, s_r_47__52_, s_r_47__51_, s_r_47__50_, s_r_47__49_, s_r_47__48_, s_r_47__47_, s_r_47__46_, s_r_47__45_, s_r_47__44_, s_r_47__43_, s_r_47__42_, s_r_47__41_, s_r_47__40_, s_r_47__39_, s_r_47__38_, s_r_47__37_, s_r_47__36_, s_r_47__35_, s_r_47__34_, s_r_47__33_, s_r_47__32_, s_r_47__31_, s_r_47__30_, s_r_47__29_, s_r_47__28_, s_r_47__27_, s_r_47__26_, s_r_47__25_, s_r_47__24_, s_r_47__23_, s_r_47__22_, s_r_47__21_, s_r_47__20_, s_r_47__19_, s_r_47__18_, s_r_47__17_, s_r_47__16_, s_r_47__15_, s_r_47__14_, s_r_47__13_, s_r_47__12_, s_r_47__11_, s_r_47__10_, s_r_47__9_, s_r_47__8_, s_r_47__7_, s_r_47__6_, s_r_47__5_, s_r_47__4_, s_r_47__3_, s_r_47__2_, s_r_47__1_, s_r_47__0_ }),
    .c_o(c_r[47]),
    .prod_accum_o({ prod_accum_47__48_, prod_accum_47__47_, prod_accum_47__46_, prod_accum_47__45_, prod_accum_47__44_, prod_accum_47__43_, prod_accum_47__42_, prod_accum_47__41_, prod_accum_47__40_, prod_accum_47__39_, prod_accum_47__38_, prod_accum_47__37_, prod_accum_47__36_, prod_accum_47__35_, prod_accum_47__34_, prod_accum_47__33_, prod_accum_47__32_, prod_accum_47__31_, prod_accum_47__30_, prod_accum_47__29_, prod_accum_47__28_, prod_accum_47__27_, prod_accum_47__26_, prod_accum_47__25_, prod_accum_47__24_, prod_accum_47__23_, prod_accum_47__22_, prod_accum_47__21_, prod_accum_47__20_, prod_accum_47__19_, prod_accum_47__18_, prod_accum_47__17_, prod_accum_47__16_, prod_accum_47__15_, prod_accum_47__14_, prod_accum_47__13_, prod_accum_47__12_, prod_accum_47__11_, prod_accum_47__10_, prod_accum_47__9_, prod_accum_47__8_, prod_accum_47__7_, prod_accum_47__6_, prod_accum_47__5_, prod_accum_47__4_, prod_accum_47__3_, prod_accum_47__2_, prod_accum_47__1_, prod_accum_47__0_ })
  );


  bsg_mul_array_row_128_48_x
  genblk1_48__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[6143:6016]),
    .b_i(b_r[6143:6016]),
    .s_i({ s_r_47__127_, s_r_47__126_, s_r_47__125_, s_r_47__124_, s_r_47__123_, s_r_47__122_, s_r_47__121_, s_r_47__120_, s_r_47__119_, s_r_47__118_, s_r_47__117_, s_r_47__116_, s_r_47__115_, s_r_47__114_, s_r_47__113_, s_r_47__112_, s_r_47__111_, s_r_47__110_, s_r_47__109_, s_r_47__108_, s_r_47__107_, s_r_47__106_, s_r_47__105_, s_r_47__104_, s_r_47__103_, s_r_47__102_, s_r_47__101_, s_r_47__100_, s_r_47__99_, s_r_47__98_, s_r_47__97_, s_r_47__96_, s_r_47__95_, s_r_47__94_, s_r_47__93_, s_r_47__92_, s_r_47__91_, s_r_47__90_, s_r_47__89_, s_r_47__88_, s_r_47__87_, s_r_47__86_, s_r_47__85_, s_r_47__84_, s_r_47__83_, s_r_47__82_, s_r_47__81_, s_r_47__80_, s_r_47__79_, s_r_47__78_, s_r_47__77_, s_r_47__76_, s_r_47__75_, s_r_47__74_, s_r_47__73_, s_r_47__72_, s_r_47__71_, s_r_47__70_, s_r_47__69_, s_r_47__68_, s_r_47__67_, s_r_47__66_, s_r_47__65_, s_r_47__64_, s_r_47__63_, s_r_47__62_, s_r_47__61_, s_r_47__60_, s_r_47__59_, s_r_47__58_, s_r_47__57_, s_r_47__56_, s_r_47__55_, s_r_47__54_, s_r_47__53_, s_r_47__52_, s_r_47__51_, s_r_47__50_, s_r_47__49_, s_r_47__48_, s_r_47__47_, s_r_47__46_, s_r_47__45_, s_r_47__44_, s_r_47__43_, s_r_47__42_, s_r_47__41_, s_r_47__40_, s_r_47__39_, s_r_47__38_, s_r_47__37_, s_r_47__36_, s_r_47__35_, s_r_47__34_, s_r_47__33_, s_r_47__32_, s_r_47__31_, s_r_47__30_, s_r_47__29_, s_r_47__28_, s_r_47__27_, s_r_47__26_, s_r_47__25_, s_r_47__24_, s_r_47__23_, s_r_47__22_, s_r_47__21_, s_r_47__20_, s_r_47__19_, s_r_47__18_, s_r_47__17_, s_r_47__16_, s_r_47__15_, s_r_47__14_, s_r_47__13_, s_r_47__12_, s_r_47__11_, s_r_47__10_, s_r_47__9_, s_r_47__8_, s_r_47__7_, s_r_47__6_, s_r_47__5_, s_r_47__4_, s_r_47__3_, s_r_47__2_, s_r_47__1_, s_r_47__0_ }),
    .c_i(c_r[47]),
    .prod_accum_i({ prod_accum_47__48_, prod_accum_47__47_, prod_accum_47__46_, prod_accum_47__45_, prod_accum_47__44_, prod_accum_47__43_, prod_accum_47__42_, prod_accum_47__41_, prod_accum_47__40_, prod_accum_47__39_, prod_accum_47__38_, prod_accum_47__37_, prod_accum_47__36_, prod_accum_47__35_, prod_accum_47__34_, prod_accum_47__33_, prod_accum_47__32_, prod_accum_47__31_, prod_accum_47__30_, prod_accum_47__29_, prod_accum_47__28_, prod_accum_47__27_, prod_accum_47__26_, prod_accum_47__25_, prod_accum_47__24_, prod_accum_47__23_, prod_accum_47__22_, prod_accum_47__21_, prod_accum_47__20_, prod_accum_47__19_, prod_accum_47__18_, prod_accum_47__17_, prod_accum_47__16_, prod_accum_47__15_, prod_accum_47__14_, prod_accum_47__13_, prod_accum_47__12_, prod_accum_47__11_, prod_accum_47__10_, prod_accum_47__9_, prod_accum_47__8_, prod_accum_47__7_, prod_accum_47__6_, prod_accum_47__5_, prod_accum_47__4_, prod_accum_47__3_, prod_accum_47__2_, prod_accum_47__1_, prod_accum_47__0_ }),
    .a_o(a_r[6271:6144]),
    .b_o(b_r[6271:6144]),
    .s_o({ s_r_48__127_, s_r_48__126_, s_r_48__125_, s_r_48__124_, s_r_48__123_, s_r_48__122_, s_r_48__121_, s_r_48__120_, s_r_48__119_, s_r_48__118_, s_r_48__117_, s_r_48__116_, s_r_48__115_, s_r_48__114_, s_r_48__113_, s_r_48__112_, s_r_48__111_, s_r_48__110_, s_r_48__109_, s_r_48__108_, s_r_48__107_, s_r_48__106_, s_r_48__105_, s_r_48__104_, s_r_48__103_, s_r_48__102_, s_r_48__101_, s_r_48__100_, s_r_48__99_, s_r_48__98_, s_r_48__97_, s_r_48__96_, s_r_48__95_, s_r_48__94_, s_r_48__93_, s_r_48__92_, s_r_48__91_, s_r_48__90_, s_r_48__89_, s_r_48__88_, s_r_48__87_, s_r_48__86_, s_r_48__85_, s_r_48__84_, s_r_48__83_, s_r_48__82_, s_r_48__81_, s_r_48__80_, s_r_48__79_, s_r_48__78_, s_r_48__77_, s_r_48__76_, s_r_48__75_, s_r_48__74_, s_r_48__73_, s_r_48__72_, s_r_48__71_, s_r_48__70_, s_r_48__69_, s_r_48__68_, s_r_48__67_, s_r_48__66_, s_r_48__65_, s_r_48__64_, s_r_48__63_, s_r_48__62_, s_r_48__61_, s_r_48__60_, s_r_48__59_, s_r_48__58_, s_r_48__57_, s_r_48__56_, s_r_48__55_, s_r_48__54_, s_r_48__53_, s_r_48__52_, s_r_48__51_, s_r_48__50_, s_r_48__49_, s_r_48__48_, s_r_48__47_, s_r_48__46_, s_r_48__45_, s_r_48__44_, s_r_48__43_, s_r_48__42_, s_r_48__41_, s_r_48__40_, s_r_48__39_, s_r_48__38_, s_r_48__37_, s_r_48__36_, s_r_48__35_, s_r_48__34_, s_r_48__33_, s_r_48__32_, s_r_48__31_, s_r_48__30_, s_r_48__29_, s_r_48__28_, s_r_48__27_, s_r_48__26_, s_r_48__25_, s_r_48__24_, s_r_48__23_, s_r_48__22_, s_r_48__21_, s_r_48__20_, s_r_48__19_, s_r_48__18_, s_r_48__17_, s_r_48__16_, s_r_48__15_, s_r_48__14_, s_r_48__13_, s_r_48__12_, s_r_48__11_, s_r_48__10_, s_r_48__9_, s_r_48__8_, s_r_48__7_, s_r_48__6_, s_r_48__5_, s_r_48__4_, s_r_48__3_, s_r_48__2_, s_r_48__1_, s_r_48__0_ }),
    .c_o(c_r[48]),
    .prod_accum_o({ prod_accum_48__49_, prod_accum_48__48_, prod_accum_48__47_, prod_accum_48__46_, prod_accum_48__45_, prod_accum_48__44_, prod_accum_48__43_, prod_accum_48__42_, prod_accum_48__41_, prod_accum_48__40_, prod_accum_48__39_, prod_accum_48__38_, prod_accum_48__37_, prod_accum_48__36_, prod_accum_48__35_, prod_accum_48__34_, prod_accum_48__33_, prod_accum_48__32_, prod_accum_48__31_, prod_accum_48__30_, prod_accum_48__29_, prod_accum_48__28_, prod_accum_48__27_, prod_accum_48__26_, prod_accum_48__25_, prod_accum_48__24_, prod_accum_48__23_, prod_accum_48__22_, prod_accum_48__21_, prod_accum_48__20_, prod_accum_48__19_, prod_accum_48__18_, prod_accum_48__17_, prod_accum_48__16_, prod_accum_48__15_, prod_accum_48__14_, prod_accum_48__13_, prod_accum_48__12_, prod_accum_48__11_, prod_accum_48__10_, prod_accum_48__9_, prod_accum_48__8_, prod_accum_48__7_, prod_accum_48__6_, prod_accum_48__5_, prod_accum_48__4_, prod_accum_48__3_, prod_accum_48__2_, prod_accum_48__1_, prod_accum_48__0_ })
  );


  bsg_mul_array_row_128_49_x
  genblk1_49__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[6271:6144]),
    .b_i(b_r[6271:6144]),
    .s_i({ s_r_48__127_, s_r_48__126_, s_r_48__125_, s_r_48__124_, s_r_48__123_, s_r_48__122_, s_r_48__121_, s_r_48__120_, s_r_48__119_, s_r_48__118_, s_r_48__117_, s_r_48__116_, s_r_48__115_, s_r_48__114_, s_r_48__113_, s_r_48__112_, s_r_48__111_, s_r_48__110_, s_r_48__109_, s_r_48__108_, s_r_48__107_, s_r_48__106_, s_r_48__105_, s_r_48__104_, s_r_48__103_, s_r_48__102_, s_r_48__101_, s_r_48__100_, s_r_48__99_, s_r_48__98_, s_r_48__97_, s_r_48__96_, s_r_48__95_, s_r_48__94_, s_r_48__93_, s_r_48__92_, s_r_48__91_, s_r_48__90_, s_r_48__89_, s_r_48__88_, s_r_48__87_, s_r_48__86_, s_r_48__85_, s_r_48__84_, s_r_48__83_, s_r_48__82_, s_r_48__81_, s_r_48__80_, s_r_48__79_, s_r_48__78_, s_r_48__77_, s_r_48__76_, s_r_48__75_, s_r_48__74_, s_r_48__73_, s_r_48__72_, s_r_48__71_, s_r_48__70_, s_r_48__69_, s_r_48__68_, s_r_48__67_, s_r_48__66_, s_r_48__65_, s_r_48__64_, s_r_48__63_, s_r_48__62_, s_r_48__61_, s_r_48__60_, s_r_48__59_, s_r_48__58_, s_r_48__57_, s_r_48__56_, s_r_48__55_, s_r_48__54_, s_r_48__53_, s_r_48__52_, s_r_48__51_, s_r_48__50_, s_r_48__49_, s_r_48__48_, s_r_48__47_, s_r_48__46_, s_r_48__45_, s_r_48__44_, s_r_48__43_, s_r_48__42_, s_r_48__41_, s_r_48__40_, s_r_48__39_, s_r_48__38_, s_r_48__37_, s_r_48__36_, s_r_48__35_, s_r_48__34_, s_r_48__33_, s_r_48__32_, s_r_48__31_, s_r_48__30_, s_r_48__29_, s_r_48__28_, s_r_48__27_, s_r_48__26_, s_r_48__25_, s_r_48__24_, s_r_48__23_, s_r_48__22_, s_r_48__21_, s_r_48__20_, s_r_48__19_, s_r_48__18_, s_r_48__17_, s_r_48__16_, s_r_48__15_, s_r_48__14_, s_r_48__13_, s_r_48__12_, s_r_48__11_, s_r_48__10_, s_r_48__9_, s_r_48__8_, s_r_48__7_, s_r_48__6_, s_r_48__5_, s_r_48__4_, s_r_48__3_, s_r_48__2_, s_r_48__1_, s_r_48__0_ }),
    .c_i(c_r[48]),
    .prod_accum_i({ prod_accum_48__49_, prod_accum_48__48_, prod_accum_48__47_, prod_accum_48__46_, prod_accum_48__45_, prod_accum_48__44_, prod_accum_48__43_, prod_accum_48__42_, prod_accum_48__41_, prod_accum_48__40_, prod_accum_48__39_, prod_accum_48__38_, prod_accum_48__37_, prod_accum_48__36_, prod_accum_48__35_, prod_accum_48__34_, prod_accum_48__33_, prod_accum_48__32_, prod_accum_48__31_, prod_accum_48__30_, prod_accum_48__29_, prod_accum_48__28_, prod_accum_48__27_, prod_accum_48__26_, prod_accum_48__25_, prod_accum_48__24_, prod_accum_48__23_, prod_accum_48__22_, prod_accum_48__21_, prod_accum_48__20_, prod_accum_48__19_, prod_accum_48__18_, prod_accum_48__17_, prod_accum_48__16_, prod_accum_48__15_, prod_accum_48__14_, prod_accum_48__13_, prod_accum_48__12_, prod_accum_48__11_, prod_accum_48__10_, prod_accum_48__9_, prod_accum_48__8_, prod_accum_48__7_, prod_accum_48__6_, prod_accum_48__5_, prod_accum_48__4_, prod_accum_48__3_, prod_accum_48__2_, prod_accum_48__1_, prod_accum_48__0_ }),
    .a_o(a_r[6399:6272]),
    .b_o(b_r[6399:6272]),
    .s_o({ s_r_49__127_, s_r_49__126_, s_r_49__125_, s_r_49__124_, s_r_49__123_, s_r_49__122_, s_r_49__121_, s_r_49__120_, s_r_49__119_, s_r_49__118_, s_r_49__117_, s_r_49__116_, s_r_49__115_, s_r_49__114_, s_r_49__113_, s_r_49__112_, s_r_49__111_, s_r_49__110_, s_r_49__109_, s_r_49__108_, s_r_49__107_, s_r_49__106_, s_r_49__105_, s_r_49__104_, s_r_49__103_, s_r_49__102_, s_r_49__101_, s_r_49__100_, s_r_49__99_, s_r_49__98_, s_r_49__97_, s_r_49__96_, s_r_49__95_, s_r_49__94_, s_r_49__93_, s_r_49__92_, s_r_49__91_, s_r_49__90_, s_r_49__89_, s_r_49__88_, s_r_49__87_, s_r_49__86_, s_r_49__85_, s_r_49__84_, s_r_49__83_, s_r_49__82_, s_r_49__81_, s_r_49__80_, s_r_49__79_, s_r_49__78_, s_r_49__77_, s_r_49__76_, s_r_49__75_, s_r_49__74_, s_r_49__73_, s_r_49__72_, s_r_49__71_, s_r_49__70_, s_r_49__69_, s_r_49__68_, s_r_49__67_, s_r_49__66_, s_r_49__65_, s_r_49__64_, s_r_49__63_, s_r_49__62_, s_r_49__61_, s_r_49__60_, s_r_49__59_, s_r_49__58_, s_r_49__57_, s_r_49__56_, s_r_49__55_, s_r_49__54_, s_r_49__53_, s_r_49__52_, s_r_49__51_, s_r_49__50_, s_r_49__49_, s_r_49__48_, s_r_49__47_, s_r_49__46_, s_r_49__45_, s_r_49__44_, s_r_49__43_, s_r_49__42_, s_r_49__41_, s_r_49__40_, s_r_49__39_, s_r_49__38_, s_r_49__37_, s_r_49__36_, s_r_49__35_, s_r_49__34_, s_r_49__33_, s_r_49__32_, s_r_49__31_, s_r_49__30_, s_r_49__29_, s_r_49__28_, s_r_49__27_, s_r_49__26_, s_r_49__25_, s_r_49__24_, s_r_49__23_, s_r_49__22_, s_r_49__21_, s_r_49__20_, s_r_49__19_, s_r_49__18_, s_r_49__17_, s_r_49__16_, s_r_49__15_, s_r_49__14_, s_r_49__13_, s_r_49__12_, s_r_49__11_, s_r_49__10_, s_r_49__9_, s_r_49__8_, s_r_49__7_, s_r_49__6_, s_r_49__5_, s_r_49__4_, s_r_49__3_, s_r_49__2_, s_r_49__1_, s_r_49__0_ }),
    .c_o(c_r[49]),
    .prod_accum_o({ prod_accum_49__50_, prod_accum_49__49_, prod_accum_49__48_, prod_accum_49__47_, prod_accum_49__46_, prod_accum_49__45_, prod_accum_49__44_, prod_accum_49__43_, prod_accum_49__42_, prod_accum_49__41_, prod_accum_49__40_, prod_accum_49__39_, prod_accum_49__38_, prod_accum_49__37_, prod_accum_49__36_, prod_accum_49__35_, prod_accum_49__34_, prod_accum_49__33_, prod_accum_49__32_, prod_accum_49__31_, prod_accum_49__30_, prod_accum_49__29_, prod_accum_49__28_, prod_accum_49__27_, prod_accum_49__26_, prod_accum_49__25_, prod_accum_49__24_, prod_accum_49__23_, prod_accum_49__22_, prod_accum_49__21_, prod_accum_49__20_, prod_accum_49__19_, prod_accum_49__18_, prod_accum_49__17_, prod_accum_49__16_, prod_accum_49__15_, prod_accum_49__14_, prod_accum_49__13_, prod_accum_49__12_, prod_accum_49__11_, prod_accum_49__10_, prod_accum_49__9_, prod_accum_49__8_, prod_accum_49__7_, prod_accum_49__6_, prod_accum_49__5_, prod_accum_49__4_, prod_accum_49__3_, prod_accum_49__2_, prod_accum_49__1_, prod_accum_49__0_ })
  );


  bsg_mul_array_row_128_50_x
  genblk1_50__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[6399:6272]),
    .b_i(b_r[6399:6272]),
    .s_i({ s_r_49__127_, s_r_49__126_, s_r_49__125_, s_r_49__124_, s_r_49__123_, s_r_49__122_, s_r_49__121_, s_r_49__120_, s_r_49__119_, s_r_49__118_, s_r_49__117_, s_r_49__116_, s_r_49__115_, s_r_49__114_, s_r_49__113_, s_r_49__112_, s_r_49__111_, s_r_49__110_, s_r_49__109_, s_r_49__108_, s_r_49__107_, s_r_49__106_, s_r_49__105_, s_r_49__104_, s_r_49__103_, s_r_49__102_, s_r_49__101_, s_r_49__100_, s_r_49__99_, s_r_49__98_, s_r_49__97_, s_r_49__96_, s_r_49__95_, s_r_49__94_, s_r_49__93_, s_r_49__92_, s_r_49__91_, s_r_49__90_, s_r_49__89_, s_r_49__88_, s_r_49__87_, s_r_49__86_, s_r_49__85_, s_r_49__84_, s_r_49__83_, s_r_49__82_, s_r_49__81_, s_r_49__80_, s_r_49__79_, s_r_49__78_, s_r_49__77_, s_r_49__76_, s_r_49__75_, s_r_49__74_, s_r_49__73_, s_r_49__72_, s_r_49__71_, s_r_49__70_, s_r_49__69_, s_r_49__68_, s_r_49__67_, s_r_49__66_, s_r_49__65_, s_r_49__64_, s_r_49__63_, s_r_49__62_, s_r_49__61_, s_r_49__60_, s_r_49__59_, s_r_49__58_, s_r_49__57_, s_r_49__56_, s_r_49__55_, s_r_49__54_, s_r_49__53_, s_r_49__52_, s_r_49__51_, s_r_49__50_, s_r_49__49_, s_r_49__48_, s_r_49__47_, s_r_49__46_, s_r_49__45_, s_r_49__44_, s_r_49__43_, s_r_49__42_, s_r_49__41_, s_r_49__40_, s_r_49__39_, s_r_49__38_, s_r_49__37_, s_r_49__36_, s_r_49__35_, s_r_49__34_, s_r_49__33_, s_r_49__32_, s_r_49__31_, s_r_49__30_, s_r_49__29_, s_r_49__28_, s_r_49__27_, s_r_49__26_, s_r_49__25_, s_r_49__24_, s_r_49__23_, s_r_49__22_, s_r_49__21_, s_r_49__20_, s_r_49__19_, s_r_49__18_, s_r_49__17_, s_r_49__16_, s_r_49__15_, s_r_49__14_, s_r_49__13_, s_r_49__12_, s_r_49__11_, s_r_49__10_, s_r_49__9_, s_r_49__8_, s_r_49__7_, s_r_49__6_, s_r_49__5_, s_r_49__4_, s_r_49__3_, s_r_49__2_, s_r_49__1_, s_r_49__0_ }),
    .c_i(c_r[49]),
    .prod_accum_i({ prod_accum_49__50_, prod_accum_49__49_, prod_accum_49__48_, prod_accum_49__47_, prod_accum_49__46_, prod_accum_49__45_, prod_accum_49__44_, prod_accum_49__43_, prod_accum_49__42_, prod_accum_49__41_, prod_accum_49__40_, prod_accum_49__39_, prod_accum_49__38_, prod_accum_49__37_, prod_accum_49__36_, prod_accum_49__35_, prod_accum_49__34_, prod_accum_49__33_, prod_accum_49__32_, prod_accum_49__31_, prod_accum_49__30_, prod_accum_49__29_, prod_accum_49__28_, prod_accum_49__27_, prod_accum_49__26_, prod_accum_49__25_, prod_accum_49__24_, prod_accum_49__23_, prod_accum_49__22_, prod_accum_49__21_, prod_accum_49__20_, prod_accum_49__19_, prod_accum_49__18_, prod_accum_49__17_, prod_accum_49__16_, prod_accum_49__15_, prod_accum_49__14_, prod_accum_49__13_, prod_accum_49__12_, prod_accum_49__11_, prod_accum_49__10_, prod_accum_49__9_, prod_accum_49__8_, prod_accum_49__7_, prod_accum_49__6_, prod_accum_49__5_, prod_accum_49__4_, prod_accum_49__3_, prod_accum_49__2_, prod_accum_49__1_, prod_accum_49__0_ }),
    .a_o(a_r[6527:6400]),
    .b_o(b_r[6527:6400]),
    .s_o({ s_r_50__127_, s_r_50__126_, s_r_50__125_, s_r_50__124_, s_r_50__123_, s_r_50__122_, s_r_50__121_, s_r_50__120_, s_r_50__119_, s_r_50__118_, s_r_50__117_, s_r_50__116_, s_r_50__115_, s_r_50__114_, s_r_50__113_, s_r_50__112_, s_r_50__111_, s_r_50__110_, s_r_50__109_, s_r_50__108_, s_r_50__107_, s_r_50__106_, s_r_50__105_, s_r_50__104_, s_r_50__103_, s_r_50__102_, s_r_50__101_, s_r_50__100_, s_r_50__99_, s_r_50__98_, s_r_50__97_, s_r_50__96_, s_r_50__95_, s_r_50__94_, s_r_50__93_, s_r_50__92_, s_r_50__91_, s_r_50__90_, s_r_50__89_, s_r_50__88_, s_r_50__87_, s_r_50__86_, s_r_50__85_, s_r_50__84_, s_r_50__83_, s_r_50__82_, s_r_50__81_, s_r_50__80_, s_r_50__79_, s_r_50__78_, s_r_50__77_, s_r_50__76_, s_r_50__75_, s_r_50__74_, s_r_50__73_, s_r_50__72_, s_r_50__71_, s_r_50__70_, s_r_50__69_, s_r_50__68_, s_r_50__67_, s_r_50__66_, s_r_50__65_, s_r_50__64_, s_r_50__63_, s_r_50__62_, s_r_50__61_, s_r_50__60_, s_r_50__59_, s_r_50__58_, s_r_50__57_, s_r_50__56_, s_r_50__55_, s_r_50__54_, s_r_50__53_, s_r_50__52_, s_r_50__51_, s_r_50__50_, s_r_50__49_, s_r_50__48_, s_r_50__47_, s_r_50__46_, s_r_50__45_, s_r_50__44_, s_r_50__43_, s_r_50__42_, s_r_50__41_, s_r_50__40_, s_r_50__39_, s_r_50__38_, s_r_50__37_, s_r_50__36_, s_r_50__35_, s_r_50__34_, s_r_50__33_, s_r_50__32_, s_r_50__31_, s_r_50__30_, s_r_50__29_, s_r_50__28_, s_r_50__27_, s_r_50__26_, s_r_50__25_, s_r_50__24_, s_r_50__23_, s_r_50__22_, s_r_50__21_, s_r_50__20_, s_r_50__19_, s_r_50__18_, s_r_50__17_, s_r_50__16_, s_r_50__15_, s_r_50__14_, s_r_50__13_, s_r_50__12_, s_r_50__11_, s_r_50__10_, s_r_50__9_, s_r_50__8_, s_r_50__7_, s_r_50__6_, s_r_50__5_, s_r_50__4_, s_r_50__3_, s_r_50__2_, s_r_50__1_, s_r_50__0_ }),
    .c_o(c_r[50]),
    .prod_accum_o({ prod_accum_50__51_, prod_accum_50__50_, prod_accum_50__49_, prod_accum_50__48_, prod_accum_50__47_, prod_accum_50__46_, prod_accum_50__45_, prod_accum_50__44_, prod_accum_50__43_, prod_accum_50__42_, prod_accum_50__41_, prod_accum_50__40_, prod_accum_50__39_, prod_accum_50__38_, prod_accum_50__37_, prod_accum_50__36_, prod_accum_50__35_, prod_accum_50__34_, prod_accum_50__33_, prod_accum_50__32_, prod_accum_50__31_, prod_accum_50__30_, prod_accum_50__29_, prod_accum_50__28_, prod_accum_50__27_, prod_accum_50__26_, prod_accum_50__25_, prod_accum_50__24_, prod_accum_50__23_, prod_accum_50__22_, prod_accum_50__21_, prod_accum_50__20_, prod_accum_50__19_, prod_accum_50__18_, prod_accum_50__17_, prod_accum_50__16_, prod_accum_50__15_, prod_accum_50__14_, prod_accum_50__13_, prod_accum_50__12_, prod_accum_50__11_, prod_accum_50__10_, prod_accum_50__9_, prod_accum_50__8_, prod_accum_50__7_, prod_accum_50__6_, prod_accum_50__5_, prod_accum_50__4_, prod_accum_50__3_, prod_accum_50__2_, prod_accum_50__1_, prod_accum_50__0_ })
  );


  bsg_mul_array_row_128_51_x
  genblk1_51__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[6527:6400]),
    .b_i(b_r[6527:6400]),
    .s_i({ s_r_50__127_, s_r_50__126_, s_r_50__125_, s_r_50__124_, s_r_50__123_, s_r_50__122_, s_r_50__121_, s_r_50__120_, s_r_50__119_, s_r_50__118_, s_r_50__117_, s_r_50__116_, s_r_50__115_, s_r_50__114_, s_r_50__113_, s_r_50__112_, s_r_50__111_, s_r_50__110_, s_r_50__109_, s_r_50__108_, s_r_50__107_, s_r_50__106_, s_r_50__105_, s_r_50__104_, s_r_50__103_, s_r_50__102_, s_r_50__101_, s_r_50__100_, s_r_50__99_, s_r_50__98_, s_r_50__97_, s_r_50__96_, s_r_50__95_, s_r_50__94_, s_r_50__93_, s_r_50__92_, s_r_50__91_, s_r_50__90_, s_r_50__89_, s_r_50__88_, s_r_50__87_, s_r_50__86_, s_r_50__85_, s_r_50__84_, s_r_50__83_, s_r_50__82_, s_r_50__81_, s_r_50__80_, s_r_50__79_, s_r_50__78_, s_r_50__77_, s_r_50__76_, s_r_50__75_, s_r_50__74_, s_r_50__73_, s_r_50__72_, s_r_50__71_, s_r_50__70_, s_r_50__69_, s_r_50__68_, s_r_50__67_, s_r_50__66_, s_r_50__65_, s_r_50__64_, s_r_50__63_, s_r_50__62_, s_r_50__61_, s_r_50__60_, s_r_50__59_, s_r_50__58_, s_r_50__57_, s_r_50__56_, s_r_50__55_, s_r_50__54_, s_r_50__53_, s_r_50__52_, s_r_50__51_, s_r_50__50_, s_r_50__49_, s_r_50__48_, s_r_50__47_, s_r_50__46_, s_r_50__45_, s_r_50__44_, s_r_50__43_, s_r_50__42_, s_r_50__41_, s_r_50__40_, s_r_50__39_, s_r_50__38_, s_r_50__37_, s_r_50__36_, s_r_50__35_, s_r_50__34_, s_r_50__33_, s_r_50__32_, s_r_50__31_, s_r_50__30_, s_r_50__29_, s_r_50__28_, s_r_50__27_, s_r_50__26_, s_r_50__25_, s_r_50__24_, s_r_50__23_, s_r_50__22_, s_r_50__21_, s_r_50__20_, s_r_50__19_, s_r_50__18_, s_r_50__17_, s_r_50__16_, s_r_50__15_, s_r_50__14_, s_r_50__13_, s_r_50__12_, s_r_50__11_, s_r_50__10_, s_r_50__9_, s_r_50__8_, s_r_50__7_, s_r_50__6_, s_r_50__5_, s_r_50__4_, s_r_50__3_, s_r_50__2_, s_r_50__1_, s_r_50__0_ }),
    .c_i(c_r[50]),
    .prod_accum_i({ prod_accum_50__51_, prod_accum_50__50_, prod_accum_50__49_, prod_accum_50__48_, prod_accum_50__47_, prod_accum_50__46_, prod_accum_50__45_, prod_accum_50__44_, prod_accum_50__43_, prod_accum_50__42_, prod_accum_50__41_, prod_accum_50__40_, prod_accum_50__39_, prod_accum_50__38_, prod_accum_50__37_, prod_accum_50__36_, prod_accum_50__35_, prod_accum_50__34_, prod_accum_50__33_, prod_accum_50__32_, prod_accum_50__31_, prod_accum_50__30_, prod_accum_50__29_, prod_accum_50__28_, prod_accum_50__27_, prod_accum_50__26_, prod_accum_50__25_, prod_accum_50__24_, prod_accum_50__23_, prod_accum_50__22_, prod_accum_50__21_, prod_accum_50__20_, prod_accum_50__19_, prod_accum_50__18_, prod_accum_50__17_, prod_accum_50__16_, prod_accum_50__15_, prod_accum_50__14_, prod_accum_50__13_, prod_accum_50__12_, prod_accum_50__11_, prod_accum_50__10_, prod_accum_50__9_, prod_accum_50__8_, prod_accum_50__7_, prod_accum_50__6_, prod_accum_50__5_, prod_accum_50__4_, prod_accum_50__3_, prod_accum_50__2_, prod_accum_50__1_, prod_accum_50__0_ }),
    .a_o(a_r[6655:6528]),
    .b_o(b_r[6655:6528]),
    .s_o({ s_r_51__127_, s_r_51__126_, s_r_51__125_, s_r_51__124_, s_r_51__123_, s_r_51__122_, s_r_51__121_, s_r_51__120_, s_r_51__119_, s_r_51__118_, s_r_51__117_, s_r_51__116_, s_r_51__115_, s_r_51__114_, s_r_51__113_, s_r_51__112_, s_r_51__111_, s_r_51__110_, s_r_51__109_, s_r_51__108_, s_r_51__107_, s_r_51__106_, s_r_51__105_, s_r_51__104_, s_r_51__103_, s_r_51__102_, s_r_51__101_, s_r_51__100_, s_r_51__99_, s_r_51__98_, s_r_51__97_, s_r_51__96_, s_r_51__95_, s_r_51__94_, s_r_51__93_, s_r_51__92_, s_r_51__91_, s_r_51__90_, s_r_51__89_, s_r_51__88_, s_r_51__87_, s_r_51__86_, s_r_51__85_, s_r_51__84_, s_r_51__83_, s_r_51__82_, s_r_51__81_, s_r_51__80_, s_r_51__79_, s_r_51__78_, s_r_51__77_, s_r_51__76_, s_r_51__75_, s_r_51__74_, s_r_51__73_, s_r_51__72_, s_r_51__71_, s_r_51__70_, s_r_51__69_, s_r_51__68_, s_r_51__67_, s_r_51__66_, s_r_51__65_, s_r_51__64_, s_r_51__63_, s_r_51__62_, s_r_51__61_, s_r_51__60_, s_r_51__59_, s_r_51__58_, s_r_51__57_, s_r_51__56_, s_r_51__55_, s_r_51__54_, s_r_51__53_, s_r_51__52_, s_r_51__51_, s_r_51__50_, s_r_51__49_, s_r_51__48_, s_r_51__47_, s_r_51__46_, s_r_51__45_, s_r_51__44_, s_r_51__43_, s_r_51__42_, s_r_51__41_, s_r_51__40_, s_r_51__39_, s_r_51__38_, s_r_51__37_, s_r_51__36_, s_r_51__35_, s_r_51__34_, s_r_51__33_, s_r_51__32_, s_r_51__31_, s_r_51__30_, s_r_51__29_, s_r_51__28_, s_r_51__27_, s_r_51__26_, s_r_51__25_, s_r_51__24_, s_r_51__23_, s_r_51__22_, s_r_51__21_, s_r_51__20_, s_r_51__19_, s_r_51__18_, s_r_51__17_, s_r_51__16_, s_r_51__15_, s_r_51__14_, s_r_51__13_, s_r_51__12_, s_r_51__11_, s_r_51__10_, s_r_51__9_, s_r_51__8_, s_r_51__7_, s_r_51__6_, s_r_51__5_, s_r_51__4_, s_r_51__3_, s_r_51__2_, s_r_51__1_, s_r_51__0_ }),
    .c_o(c_r[51]),
    .prod_accum_o({ prod_accum_51__52_, prod_accum_51__51_, prod_accum_51__50_, prod_accum_51__49_, prod_accum_51__48_, prod_accum_51__47_, prod_accum_51__46_, prod_accum_51__45_, prod_accum_51__44_, prod_accum_51__43_, prod_accum_51__42_, prod_accum_51__41_, prod_accum_51__40_, prod_accum_51__39_, prod_accum_51__38_, prod_accum_51__37_, prod_accum_51__36_, prod_accum_51__35_, prod_accum_51__34_, prod_accum_51__33_, prod_accum_51__32_, prod_accum_51__31_, prod_accum_51__30_, prod_accum_51__29_, prod_accum_51__28_, prod_accum_51__27_, prod_accum_51__26_, prod_accum_51__25_, prod_accum_51__24_, prod_accum_51__23_, prod_accum_51__22_, prod_accum_51__21_, prod_accum_51__20_, prod_accum_51__19_, prod_accum_51__18_, prod_accum_51__17_, prod_accum_51__16_, prod_accum_51__15_, prod_accum_51__14_, prod_accum_51__13_, prod_accum_51__12_, prod_accum_51__11_, prod_accum_51__10_, prod_accum_51__9_, prod_accum_51__8_, prod_accum_51__7_, prod_accum_51__6_, prod_accum_51__5_, prod_accum_51__4_, prod_accum_51__3_, prod_accum_51__2_, prod_accum_51__1_, prod_accum_51__0_ })
  );


  bsg_mul_array_row_128_52_x
  genblk1_52__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[6655:6528]),
    .b_i(b_r[6655:6528]),
    .s_i({ s_r_51__127_, s_r_51__126_, s_r_51__125_, s_r_51__124_, s_r_51__123_, s_r_51__122_, s_r_51__121_, s_r_51__120_, s_r_51__119_, s_r_51__118_, s_r_51__117_, s_r_51__116_, s_r_51__115_, s_r_51__114_, s_r_51__113_, s_r_51__112_, s_r_51__111_, s_r_51__110_, s_r_51__109_, s_r_51__108_, s_r_51__107_, s_r_51__106_, s_r_51__105_, s_r_51__104_, s_r_51__103_, s_r_51__102_, s_r_51__101_, s_r_51__100_, s_r_51__99_, s_r_51__98_, s_r_51__97_, s_r_51__96_, s_r_51__95_, s_r_51__94_, s_r_51__93_, s_r_51__92_, s_r_51__91_, s_r_51__90_, s_r_51__89_, s_r_51__88_, s_r_51__87_, s_r_51__86_, s_r_51__85_, s_r_51__84_, s_r_51__83_, s_r_51__82_, s_r_51__81_, s_r_51__80_, s_r_51__79_, s_r_51__78_, s_r_51__77_, s_r_51__76_, s_r_51__75_, s_r_51__74_, s_r_51__73_, s_r_51__72_, s_r_51__71_, s_r_51__70_, s_r_51__69_, s_r_51__68_, s_r_51__67_, s_r_51__66_, s_r_51__65_, s_r_51__64_, s_r_51__63_, s_r_51__62_, s_r_51__61_, s_r_51__60_, s_r_51__59_, s_r_51__58_, s_r_51__57_, s_r_51__56_, s_r_51__55_, s_r_51__54_, s_r_51__53_, s_r_51__52_, s_r_51__51_, s_r_51__50_, s_r_51__49_, s_r_51__48_, s_r_51__47_, s_r_51__46_, s_r_51__45_, s_r_51__44_, s_r_51__43_, s_r_51__42_, s_r_51__41_, s_r_51__40_, s_r_51__39_, s_r_51__38_, s_r_51__37_, s_r_51__36_, s_r_51__35_, s_r_51__34_, s_r_51__33_, s_r_51__32_, s_r_51__31_, s_r_51__30_, s_r_51__29_, s_r_51__28_, s_r_51__27_, s_r_51__26_, s_r_51__25_, s_r_51__24_, s_r_51__23_, s_r_51__22_, s_r_51__21_, s_r_51__20_, s_r_51__19_, s_r_51__18_, s_r_51__17_, s_r_51__16_, s_r_51__15_, s_r_51__14_, s_r_51__13_, s_r_51__12_, s_r_51__11_, s_r_51__10_, s_r_51__9_, s_r_51__8_, s_r_51__7_, s_r_51__6_, s_r_51__5_, s_r_51__4_, s_r_51__3_, s_r_51__2_, s_r_51__1_, s_r_51__0_ }),
    .c_i(c_r[51]),
    .prod_accum_i({ prod_accum_51__52_, prod_accum_51__51_, prod_accum_51__50_, prod_accum_51__49_, prod_accum_51__48_, prod_accum_51__47_, prod_accum_51__46_, prod_accum_51__45_, prod_accum_51__44_, prod_accum_51__43_, prod_accum_51__42_, prod_accum_51__41_, prod_accum_51__40_, prod_accum_51__39_, prod_accum_51__38_, prod_accum_51__37_, prod_accum_51__36_, prod_accum_51__35_, prod_accum_51__34_, prod_accum_51__33_, prod_accum_51__32_, prod_accum_51__31_, prod_accum_51__30_, prod_accum_51__29_, prod_accum_51__28_, prod_accum_51__27_, prod_accum_51__26_, prod_accum_51__25_, prod_accum_51__24_, prod_accum_51__23_, prod_accum_51__22_, prod_accum_51__21_, prod_accum_51__20_, prod_accum_51__19_, prod_accum_51__18_, prod_accum_51__17_, prod_accum_51__16_, prod_accum_51__15_, prod_accum_51__14_, prod_accum_51__13_, prod_accum_51__12_, prod_accum_51__11_, prod_accum_51__10_, prod_accum_51__9_, prod_accum_51__8_, prod_accum_51__7_, prod_accum_51__6_, prod_accum_51__5_, prod_accum_51__4_, prod_accum_51__3_, prod_accum_51__2_, prod_accum_51__1_, prod_accum_51__0_ }),
    .a_o(a_r[6783:6656]),
    .b_o(b_r[6783:6656]),
    .s_o({ s_r_52__127_, s_r_52__126_, s_r_52__125_, s_r_52__124_, s_r_52__123_, s_r_52__122_, s_r_52__121_, s_r_52__120_, s_r_52__119_, s_r_52__118_, s_r_52__117_, s_r_52__116_, s_r_52__115_, s_r_52__114_, s_r_52__113_, s_r_52__112_, s_r_52__111_, s_r_52__110_, s_r_52__109_, s_r_52__108_, s_r_52__107_, s_r_52__106_, s_r_52__105_, s_r_52__104_, s_r_52__103_, s_r_52__102_, s_r_52__101_, s_r_52__100_, s_r_52__99_, s_r_52__98_, s_r_52__97_, s_r_52__96_, s_r_52__95_, s_r_52__94_, s_r_52__93_, s_r_52__92_, s_r_52__91_, s_r_52__90_, s_r_52__89_, s_r_52__88_, s_r_52__87_, s_r_52__86_, s_r_52__85_, s_r_52__84_, s_r_52__83_, s_r_52__82_, s_r_52__81_, s_r_52__80_, s_r_52__79_, s_r_52__78_, s_r_52__77_, s_r_52__76_, s_r_52__75_, s_r_52__74_, s_r_52__73_, s_r_52__72_, s_r_52__71_, s_r_52__70_, s_r_52__69_, s_r_52__68_, s_r_52__67_, s_r_52__66_, s_r_52__65_, s_r_52__64_, s_r_52__63_, s_r_52__62_, s_r_52__61_, s_r_52__60_, s_r_52__59_, s_r_52__58_, s_r_52__57_, s_r_52__56_, s_r_52__55_, s_r_52__54_, s_r_52__53_, s_r_52__52_, s_r_52__51_, s_r_52__50_, s_r_52__49_, s_r_52__48_, s_r_52__47_, s_r_52__46_, s_r_52__45_, s_r_52__44_, s_r_52__43_, s_r_52__42_, s_r_52__41_, s_r_52__40_, s_r_52__39_, s_r_52__38_, s_r_52__37_, s_r_52__36_, s_r_52__35_, s_r_52__34_, s_r_52__33_, s_r_52__32_, s_r_52__31_, s_r_52__30_, s_r_52__29_, s_r_52__28_, s_r_52__27_, s_r_52__26_, s_r_52__25_, s_r_52__24_, s_r_52__23_, s_r_52__22_, s_r_52__21_, s_r_52__20_, s_r_52__19_, s_r_52__18_, s_r_52__17_, s_r_52__16_, s_r_52__15_, s_r_52__14_, s_r_52__13_, s_r_52__12_, s_r_52__11_, s_r_52__10_, s_r_52__9_, s_r_52__8_, s_r_52__7_, s_r_52__6_, s_r_52__5_, s_r_52__4_, s_r_52__3_, s_r_52__2_, s_r_52__1_, s_r_52__0_ }),
    .c_o(c_r[52]),
    .prod_accum_o({ prod_accum_52__53_, prod_accum_52__52_, prod_accum_52__51_, prod_accum_52__50_, prod_accum_52__49_, prod_accum_52__48_, prod_accum_52__47_, prod_accum_52__46_, prod_accum_52__45_, prod_accum_52__44_, prod_accum_52__43_, prod_accum_52__42_, prod_accum_52__41_, prod_accum_52__40_, prod_accum_52__39_, prod_accum_52__38_, prod_accum_52__37_, prod_accum_52__36_, prod_accum_52__35_, prod_accum_52__34_, prod_accum_52__33_, prod_accum_52__32_, prod_accum_52__31_, prod_accum_52__30_, prod_accum_52__29_, prod_accum_52__28_, prod_accum_52__27_, prod_accum_52__26_, prod_accum_52__25_, prod_accum_52__24_, prod_accum_52__23_, prod_accum_52__22_, prod_accum_52__21_, prod_accum_52__20_, prod_accum_52__19_, prod_accum_52__18_, prod_accum_52__17_, prod_accum_52__16_, prod_accum_52__15_, prod_accum_52__14_, prod_accum_52__13_, prod_accum_52__12_, prod_accum_52__11_, prod_accum_52__10_, prod_accum_52__9_, prod_accum_52__8_, prod_accum_52__7_, prod_accum_52__6_, prod_accum_52__5_, prod_accum_52__4_, prod_accum_52__3_, prod_accum_52__2_, prod_accum_52__1_, prod_accum_52__0_ })
  );


  bsg_mul_array_row_128_53_x
  genblk1_53__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[6783:6656]),
    .b_i(b_r[6783:6656]),
    .s_i({ s_r_52__127_, s_r_52__126_, s_r_52__125_, s_r_52__124_, s_r_52__123_, s_r_52__122_, s_r_52__121_, s_r_52__120_, s_r_52__119_, s_r_52__118_, s_r_52__117_, s_r_52__116_, s_r_52__115_, s_r_52__114_, s_r_52__113_, s_r_52__112_, s_r_52__111_, s_r_52__110_, s_r_52__109_, s_r_52__108_, s_r_52__107_, s_r_52__106_, s_r_52__105_, s_r_52__104_, s_r_52__103_, s_r_52__102_, s_r_52__101_, s_r_52__100_, s_r_52__99_, s_r_52__98_, s_r_52__97_, s_r_52__96_, s_r_52__95_, s_r_52__94_, s_r_52__93_, s_r_52__92_, s_r_52__91_, s_r_52__90_, s_r_52__89_, s_r_52__88_, s_r_52__87_, s_r_52__86_, s_r_52__85_, s_r_52__84_, s_r_52__83_, s_r_52__82_, s_r_52__81_, s_r_52__80_, s_r_52__79_, s_r_52__78_, s_r_52__77_, s_r_52__76_, s_r_52__75_, s_r_52__74_, s_r_52__73_, s_r_52__72_, s_r_52__71_, s_r_52__70_, s_r_52__69_, s_r_52__68_, s_r_52__67_, s_r_52__66_, s_r_52__65_, s_r_52__64_, s_r_52__63_, s_r_52__62_, s_r_52__61_, s_r_52__60_, s_r_52__59_, s_r_52__58_, s_r_52__57_, s_r_52__56_, s_r_52__55_, s_r_52__54_, s_r_52__53_, s_r_52__52_, s_r_52__51_, s_r_52__50_, s_r_52__49_, s_r_52__48_, s_r_52__47_, s_r_52__46_, s_r_52__45_, s_r_52__44_, s_r_52__43_, s_r_52__42_, s_r_52__41_, s_r_52__40_, s_r_52__39_, s_r_52__38_, s_r_52__37_, s_r_52__36_, s_r_52__35_, s_r_52__34_, s_r_52__33_, s_r_52__32_, s_r_52__31_, s_r_52__30_, s_r_52__29_, s_r_52__28_, s_r_52__27_, s_r_52__26_, s_r_52__25_, s_r_52__24_, s_r_52__23_, s_r_52__22_, s_r_52__21_, s_r_52__20_, s_r_52__19_, s_r_52__18_, s_r_52__17_, s_r_52__16_, s_r_52__15_, s_r_52__14_, s_r_52__13_, s_r_52__12_, s_r_52__11_, s_r_52__10_, s_r_52__9_, s_r_52__8_, s_r_52__7_, s_r_52__6_, s_r_52__5_, s_r_52__4_, s_r_52__3_, s_r_52__2_, s_r_52__1_, s_r_52__0_ }),
    .c_i(c_r[52]),
    .prod_accum_i({ prod_accum_52__53_, prod_accum_52__52_, prod_accum_52__51_, prod_accum_52__50_, prod_accum_52__49_, prod_accum_52__48_, prod_accum_52__47_, prod_accum_52__46_, prod_accum_52__45_, prod_accum_52__44_, prod_accum_52__43_, prod_accum_52__42_, prod_accum_52__41_, prod_accum_52__40_, prod_accum_52__39_, prod_accum_52__38_, prod_accum_52__37_, prod_accum_52__36_, prod_accum_52__35_, prod_accum_52__34_, prod_accum_52__33_, prod_accum_52__32_, prod_accum_52__31_, prod_accum_52__30_, prod_accum_52__29_, prod_accum_52__28_, prod_accum_52__27_, prod_accum_52__26_, prod_accum_52__25_, prod_accum_52__24_, prod_accum_52__23_, prod_accum_52__22_, prod_accum_52__21_, prod_accum_52__20_, prod_accum_52__19_, prod_accum_52__18_, prod_accum_52__17_, prod_accum_52__16_, prod_accum_52__15_, prod_accum_52__14_, prod_accum_52__13_, prod_accum_52__12_, prod_accum_52__11_, prod_accum_52__10_, prod_accum_52__9_, prod_accum_52__8_, prod_accum_52__7_, prod_accum_52__6_, prod_accum_52__5_, prod_accum_52__4_, prod_accum_52__3_, prod_accum_52__2_, prod_accum_52__1_, prod_accum_52__0_ }),
    .a_o(a_r[6911:6784]),
    .b_o(b_r[6911:6784]),
    .s_o({ s_r_53__127_, s_r_53__126_, s_r_53__125_, s_r_53__124_, s_r_53__123_, s_r_53__122_, s_r_53__121_, s_r_53__120_, s_r_53__119_, s_r_53__118_, s_r_53__117_, s_r_53__116_, s_r_53__115_, s_r_53__114_, s_r_53__113_, s_r_53__112_, s_r_53__111_, s_r_53__110_, s_r_53__109_, s_r_53__108_, s_r_53__107_, s_r_53__106_, s_r_53__105_, s_r_53__104_, s_r_53__103_, s_r_53__102_, s_r_53__101_, s_r_53__100_, s_r_53__99_, s_r_53__98_, s_r_53__97_, s_r_53__96_, s_r_53__95_, s_r_53__94_, s_r_53__93_, s_r_53__92_, s_r_53__91_, s_r_53__90_, s_r_53__89_, s_r_53__88_, s_r_53__87_, s_r_53__86_, s_r_53__85_, s_r_53__84_, s_r_53__83_, s_r_53__82_, s_r_53__81_, s_r_53__80_, s_r_53__79_, s_r_53__78_, s_r_53__77_, s_r_53__76_, s_r_53__75_, s_r_53__74_, s_r_53__73_, s_r_53__72_, s_r_53__71_, s_r_53__70_, s_r_53__69_, s_r_53__68_, s_r_53__67_, s_r_53__66_, s_r_53__65_, s_r_53__64_, s_r_53__63_, s_r_53__62_, s_r_53__61_, s_r_53__60_, s_r_53__59_, s_r_53__58_, s_r_53__57_, s_r_53__56_, s_r_53__55_, s_r_53__54_, s_r_53__53_, s_r_53__52_, s_r_53__51_, s_r_53__50_, s_r_53__49_, s_r_53__48_, s_r_53__47_, s_r_53__46_, s_r_53__45_, s_r_53__44_, s_r_53__43_, s_r_53__42_, s_r_53__41_, s_r_53__40_, s_r_53__39_, s_r_53__38_, s_r_53__37_, s_r_53__36_, s_r_53__35_, s_r_53__34_, s_r_53__33_, s_r_53__32_, s_r_53__31_, s_r_53__30_, s_r_53__29_, s_r_53__28_, s_r_53__27_, s_r_53__26_, s_r_53__25_, s_r_53__24_, s_r_53__23_, s_r_53__22_, s_r_53__21_, s_r_53__20_, s_r_53__19_, s_r_53__18_, s_r_53__17_, s_r_53__16_, s_r_53__15_, s_r_53__14_, s_r_53__13_, s_r_53__12_, s_r_53__11_, s_r_53__10_, s_r_53__9_, s_r_53__8_, s_r_53__7_, s_r_53__6_, s_r_53__5_, s_r_53__4_, s_r_53__3_, s_r_53__2_, s_r_53__1_, s_r_53__0_ }),
    .c_o(c_r[53]),
    .prod_accum_o({ prod_accum_53__54_, prod_accum_53__53_, prod_accum_53__52_, prod_accum_53__51_, prod_accum_53__50_, prod_accum_53__49_, prod_accum_53__48_, prod_accum_53__47_, prod_accum_53__46_, prod_accum_53__45_, prod_accum_53__44_, prod_accum_53__43_, prod_accum_53__42_, prod_accum_53__41_, prod_accum_53__40_, prod_accum_53__39_, prod_accum_53__38_, prod_accum_53__37_, prod_accum_53__36_, prod_accum_53__35_, prod_accum_53__34_, prod_accum_53__33_, prod_accum_53__32_, prod_accum_53__31_, prod_accum_53__30_, prod_accum_53__29_, prod_accum_53__28_, prod_accum_53__27_, prod_accum_53__26_, prod_accum_53__25_, prod_accum_53__24_, prod_accum_53__23_, prod_accum_53__22_, prod_accum_53__21_, prod_accum_53__20_, prod_accum_53__19_, prod_accum_53__18_, prod_accum_53__17_, prod_accum_53__16_, prod_accum_53__15_, prod_accum_53__14_, prod_accum_53__13_, prod_accum_53__12_, prod_accum_53__11_, prod_accum_53__10_, prod_accum_53__9_, prod_accum_53__8_, prod_accum_53__7_, prod_accum_53__6_, prod_accum_53__5_, prod_accum_53__4_, prod_accum_53__3_, prod_accum_53__2_, prod_accum_53__1_, prod_accum_53__0_ })
  );


  bsg_mul_array_row_128_54_x
  genblk1_54__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[6911:6784]),
    .b_i(b_r[6911:6784]),
    .s_i({ s_r_53__127_, s_r_53__126_, s_r_53__125_, s_r_53__124_, s_r_53__123_, s_r_53__122_, s_r_53__121_, s_r_53__120_, s_r_53__119_, s_r_53__118_, s_r_53__117_, s_r_53__116_, s_r_53__115_, s_r_53__114_, s_r_53__113_, s_r_53__112_, s_r_53__111_, s_r_53__110_, s_r_53__109_, s_r_53__108_, s_r_53__107_, s_r_53__106_, s_r_53__105_, s_r_53__104_, s_r_53__103_, s_r_53__102_, s_r_53__101_, s_r_53__100_, s_r_53__99_, s_r_53__98_, s_r_53__97_, s_r_53__96_, s_r_53__95_, s_r_53__94_, s_r_53__93_, s_r_53__92_, s_r_53__91_, s_r_53__90_, s_r_53__89_, s_r_53__88_, s_r_53__87_, s_r_53__86_, s_r_53__85_, s_r_53__84_, s_r_53__83_, s_r_53__82_, s_r_53__81_, s_r_53__80_, s_r_53__79_, s_r_53__78_, s_r_53__77_, s_r_53__76_, s_r_53__75_, s_r_53__74_, s_r_53__73_, s_r_53__72_, s_r_53__71_, s_r_53__70_, s_r_53__69_, s_r_53__68_, s_r_53__67_, s_r_53__66_, s_r_53__65_, s_r_53__64_, s_r_53__63_, s_r_53__62_, s_r_53__61_, s_r_53__60_, s_r_53__59_, s_r_53__58_, s_r_53__57_, s_r_53__56_, s_r_53__55_, s_r_53__54_, s_r_53__53_, s_r_53__52_, s_r_53__51_, s_r_53__50_, s_r_53__49_, s_r_53__48_, s_r_53__47_, s_r_53__46_, s_r_53__45_, s_r_53__44_, s_r_53__43_, s_r_53__42_, s_r_53__41_, s_r_53__40_, s_r_53__39_, s_r_53__38_, s_r_53__37_, s_r_53__36_, s_r_53__35_, s_r_53__34_, s_r_53__33_, s_r_53__32_, s_r_53__31_, s_r_53__30_, s_r_53__29_, s_r_53__28_, s_r_53__27_, s_r_53__26_, s_r_53__25_, s_r_53__24_, s_r_53__23_, s_r_53__22_, s_r_53__21_, s_r_53__20_, s_r_53__19_, s_r_53__18_, s_r_53__17_, s_r_53__16_, s_r_53__15_, s_r_53__14_, s_r_53__13_, s_r_53__12_, s_r_53__11_, s_r_53__10_, s_r_53__9_, s_r_53__8_, s_r_53__7_, s_r_53__6_, s_r_53__5_, s_r_53__4_, s_r_53__3_, s_r_53__2_, s_r_53__1_, s_r_53__0_ }),
    .c_i(c_r[53]),
    .prod_accum_i({ prod_accum_53__54_, prod_accum_53__53_, prod_accum_53__52_, prod_accum_53__51_, prod_accum_53__50_, prod_accum_53__49_, prod_accum_53__48_, prod_accum_53__47_, prod_accum_53__46_, prod_accum_53__45_, prod_accum_53__44_, prod_accum_53__43_, prod_accum_53__42_, prod_accum_53__41_, prod_accum_53__40_, prod_accum_53__39_, prod_accum_53__38_, prod_accum_53__37_, prod_accum_53__36_, prod_accum_53__35_, prod_accum_53__34_, prod_accum_53__33_, prod_accum_53__32_, prod_accum_53__31_, prod_accum_53__30_, prod_accum_53__29_, prod_accum_53__28_, prod_accum_53__27_, prod_accum_53__26_, prod_accum_53__25_, prod_accum_53__24_, prod_accum_53__23_, prod_accum_53__22_, prod_accum_53__21_, prod_accum_53__20_, prod_accum_53__19_, prod_accum_53__18_, prod_accum_53__17_, prod_accum_53__16_, prod_accum_53__15_, prod_accum_53__14_, prod_accum_53__13_, prod_accum_53__12_, prod_accum_53__11_, prod_accum_53__10_, prod_accum_53__9_, prod_accum_53__8_, prod_accum_53__7_, prod_accum_53__6_, prod_accum_53__5_, prod_accum_53__4_, prod_accum_53__3_, prod_accum_53__2_, prod_accum_53__1_, prod_accum_53__0_ }),
    .a_o(a_r[7039:6912]),
    .b_o(b_r[7039:6912]),
    .s_o({ s_r_54__127_, s_r_54__126_, s_r_54__125_, s_r_54__124_, s_r_54__123_, s_r_54__122_, s_r_54__121_, s_r_54__120_, s_r_54__119_, s_r_54__118_, s_r_54__117_, s_r_54__116_, s_r_54__115_, s_r_54__114_, s_r_54__113_, s_r_54__112_, s_r_54__111_, s_r_54__110_, s_r_54__109_, s_r_54__108_, s_r_54__107_, s_r_54__106_, s_r_54__105_, s_r_54__104_, s_r_54__103_, s_r_54__102_, s_r_54__101_, s_r_54__100_, s_r_54__99_, s_r_54__98_, s_r_54__97_, s_r_54__96_, s_r_54__95_, s_r_54__94_, s_r_54__93_, s_r_54__92_, s_r_54__91_, s_r_54__90_, s_r_54__89_, s_r_54__88_, s_r_54__87_, s_r_54__86_, s_r_54__85_, s_r_54__84_, s_r_54__83_, s_r_54__82_, s_r_54__81_, s_r_54__80_, s_r_54__79_, s_r_54__78_, s_r_54__77_, s_r_54__76_, s_r_54__75_, s_r_54__74_, s_r_54__73_, s_r_54__72_, s_r_54__71_, s_r_54__70_, s_r_54__69_, s_r_54__68_, s_r_54__67_, s_r_54__66_, s_r_54__65_, s_r_54__64_, s_r_54__63_, s_r_54__62_, s_r_54__61_, s_r_54__60_, s_r_54__59_, s_r_54__58_, s_r_54__57_, s_r_54__56_, s_r_54__55_, s_r_54__54_, s_r_54__53_, s_r_54__52_, s_r_54__51_, s_r_54__50_, s_r_54__49_, s_r_54__48_, s_r_54__47_, s_r_54__46_, s_r_54__45_, s_r_54__44_, s_r_54__43_, s_r_54__42_, s_r_54__41_, s_r_54__40_, s_r_54__39_, s_r_54__38_, s_r_54__37_, s_r_54__36_, s_r_54__35_, s_r_54__34_, s_r_54__33_, s_r_54__32_, s_r_54__31_, s_r_54__30_, s_r_54__29_, s_r_54__28_, s_r_54__27_, s_r_54__26_, s_r_54__25_, s_r_54__24_, s_r_54__23_, s_r_54__22_, s_r_54__21_, s_r_54__20_, s_r_54__19_, s_r_54__18_, s_r_54__17_, s_r_54__16_, s_r_54__15_, s_r_54__14_, s_r_54__13_, s_r_54__12_, s_r_54__11_, s_r_54__10_, s_r_54__9_, s_r_54__8_, s_r_54__7_, s_r_54__6_, s_r_54__5_, s_r_54__4_, s_r_54__3_, s_r_54__2_, s_r_54__1_, s_r_54__0_ }),
    .c_o(c_r[54]),
    .prod_accum_o({ prod_accum_54__55_, prod_accum_54__54_, prod_accum_54__53_, prod_accum_54__52_, prod_accum_54__51_, prod_accum_54__50_, prod_accum_54__49_, prod_accum_54__48_, prod_accum_54__47_, prod_accum_54__46_, prod_accum_54__45_, prod_accum_54__44_, prod_accum_54__43_, prod_accum_54__42_, prod_accum_54__41_, prod_accum_54__40_, prod_accum_54__39_, prod_accum_54__38_, prod_accum_54__37_, prod_accum_54__36_, prod_accum_54__35_, prod_accum_54__34_, prod_accum_54__33_, prod_accum_54__32_, prod_accum_54__31_, prod_accum_54__30_, prod_accum_54__29_, prod_accum_54__28_, prod_accum_54__27_, prod_accum_54__26_, prod_accum_54__25_, prod_accum_54__24_, prod_accum_54__23_, prod_accum_54__22_, prod_accum_54__21_, prod_accum_54__20_, prod_accum_54__19_, prod_accum_54__18_, prod_accum_54__17_, prod_accum_54__16_, prod_accum_54__15_, prod_accum_54__14_, prod_accum_54__13_, prod_accum_54__12_, prod_accum_54__11_, prod_accum_54__10_, prod_accum_54__9_, prod_accum_54__8_, prod_accum_54__7_, prod_accum_54__6_, prod_accum_54__5_, prod_accum_54__4_, prod_accum_54__3_, prod_accum_54__2_, prod_accum_54__1_, prod_accum_54__0_ })
  );


  bsg_mul_array_row_128_55_x
  genblk1_55__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[7039:6912]),
    .b_i(b_r[7039:6912]),
    .s_i({ s_r_54__127_, s_r_54__126_, s_r_54__125_, s_r_54__124_, s_r_54__123_, s_r_54__122_, s_r_54__121_, s_r_54__120_, s_r_54__119_, s_r_54__118_, s_r_54__117_, s_r_54__116_, s_r_54__115_, s_r_54__114_, s_r_54__113_, s_r_54__112_, s_r_54__111_, s_r_54__110_, s_r_54__109_, s_r_54__108_, s_r_54__107_, s_r_54__106_, s_r_54__105_, s_r_54__104_, s_r_54__103_, s_r_54__102_, s_r_54__101_, s_r_54__100_, s_r_54__99_, s_r_54__98_, s_r_54__97_, s_r_54__96_, s_r_54__95_, s_r_54__94_, s_r_54__93_, s_r_54__92_, s_r_54__91_, s_r_54__90_, s_r_54__89_, s_r_54__88_, s_r_54__87_, s_r_54__86_, s_r_54__85_, s_r_54__84_, s_r_54__83_, s_r_54__82_, s_r_54__81_, s_r_54__80_, s_r_54__79_, s_r_54__78_, s_r_54__77_, s_r_54__76_, s_r_54__75_, s_r_54__74_, s_r_54__73_, s_r_54__72_, s_r_54__71_, s_r_54__70_, s_r_54__69_, s_r_54__68_, s_r_54__67_, s_r_54__66_, s_r_54__65_, s_r_54__64_, s_r_54__63_, s_r_54__62_, s_r_54__61_, s_r_54__60_, s_r_54__59_, s_r_54__58_, s_r_54__57_, s_r_54__56_, s_r_54__55_, s_r_54__54_, s_r_54__53_, s_r_54__52_, s_r_54__51_, s_r_54__50_, s_r_54__49_, s_r_54__48_, s_r_54__47_, s_r_54__46_, s_r_54__45_, s_r_54__44_, s_r_54__43_, s_r_54__42_, s_r_54__41_, s_r_54__40_, s_r_54__39_, s_r_54__38_, s_r_54__37_, s_r_54__36_, s_r_54__35_, s_r_54__34_, s_r_54__33_, s_r_54__32_, s_r_54__31_, s_r_54__30_, s_r_54__29_, s_r_54__28_, s_r_54__27_, s_r_54__26_, s_r_54__25_, s_r_54__24_, s_r_54__23_, s_r_54__22_, s_r_54__21_, s_r_54__20_, s_r_54__19_, s_r_54__18_, s_r_54__17_, s_r_54__16_, s_r_54__15_, s_r_54__14_, s_r_54__13_, s_r_54__12_, s_r_54__11_, s_r_54__10_, s_r_54__9_, s_r_54__8_, s_r_54__7_, s_r_54__6_, s_r_54__5_, s_r_54__4_, s_r_54__3_, s_r_54__2_, s_r_54__1_, s_r_54__0_ }),
    .c_i(c_r[54]),
    .prod_accum_i({ prod_accum_54__55_, prod_accum_54__54_, prod_accum_54__53_, prod_accum_54__52_, prod_accum_54__51_, prod_accum_54__50_, prod_accum_54__49_, prod_accum_54__48_, prod_accum_54__47_, prod_accum_54__46_, prod_accum_54__45_, prod_accum_54__44_, prod_accum_54__43_, prod_accum_54__42_, prod_accum_54__41_, prod_accum_54__40_, prod_accum_54__39_, prod_accum_54__38_, prod_accum_54__37_, prod_accum_54__36_, prod_accum_54__35_, prod_accum_54__34_, prod_accum_54__33_, prod_accum_54__32_, prod_accum_54__31_, prod_accum_54__30_, prod_accum_54__29_, prod_accum_54__28_, prod_accum_54__27_, prod_accum_54__26_, prod_accum_54__25_, prod_accum_54__24_, prod_accum_54__23_, prod_accum_54__22_, prod_accum_54__21_, prod_accum_54__20_, prod_accum_54__19_, prod_accum_54__18_, prod_accum_54__17_, prod_accum_54__16_, prod_accum_54__15_, prod_accum_54__14_, prod_accum_54__13_, prod_accum_54__12_, prod_accum_54__11_, prod_accum_54__10_, prod_accum_54__9_, prod_accum_54__8_, prod_accum_54__7_, prod_accum_54__6_, prod_accum_54__5_, prod_accum_54__4_, prod_accum_54__3_, prod_accum_54__2_, prod_accum_54__1_, prod_accum_54__0_ }),
    .a_o(a_r[7167:7040]),
    .b_o(b_r[7167:7040]),
    .s_o({ s_r_55__127_, s_r_55__126_, s_r_55__125_, s_r_55__124_, s_r_55__123_, s_r_55__122_, s_r_55__121_, s_r_55__120_, s_r_55__119_, s_r_55__118_, s_r_55__117_, s_r_55__116_, s_r_55__115_, s_r_55__114_, s_r_55__113_, s_r_55__112_, s_r_55__111_, s_r_55__110_, s_r_55__109_, s_r_55__108_, s_r_55__107_, s_r_55__106_, s_r_55__105_, s_r_55__104_, s_r_55__103_, s_r_55__102_, s_r_55__101_, s_r_55__100_, s_r_55__99_, s_r_55__98_, s_r_55__97_, s_r_55__96_, s_r_55__95_, s_r_55__94_, s_r_55__93_, s_r_55__92_, s_r_55__91_, s_r_55__90_, s_r_55__89_, s_r_55__88_, s_r_55__87_, s_r_55__86_, s_r_55__85_, s_r_55__84_, s_r_55__83_, s_r_55__82_, s_r_55__81_, s_r_55__80_, s_r_55__79_, s_r_55__78_, s_r_55__77_, s_r_55__76_, s_r_55__75_, s_r_55__74_, s_r_55__73_, s_r_55__72_, s_r_55__71_, s_r_55__70_, s_r_55__69_, s_r_55__68_, s_r_55__67_, s_r_55__66_, s_r_55__65_, s_r_55__64_, s_r_55__63_, s_r_55__62_, s_r_55__61_, s_r_55__60_, s_r_55__59_, s_r_55__58_, s_r_55__57_, s_r_55__56_, s_r_55__55_, s_r_55__54_, s_r_55__53_, s_r_55__52_, s_r_55__51_, s_r_55__50_, s_r_55__49_, s_r_55__48_, s_r_55__47_, s_r_55__46_, s_r_55__45_, s_r_55__44_, s_r_55__43_, s_r_55__42_, s_r_55__41_, s_r_55__40_, s_r_55__39_, s_r_55__38_, s_r_55__37_, s_r_55__36_, s_r_55__35_, s_r_55__34_, s_r_55__33_, s_r_55__32_, s_r_55__31_, s_r_55__30_, s_r_55__29_, s_r_55__28_, s_r_55__27_, s_r_55__26_, s_r_55__25_, s_r_55__24_, s_r_55__23_, s_r_55__22_, s_r_55__21_, s_r_55__20_, s_r_55__19_, s_r_55__18_, s_r_55__17_, s_r_55__16_, s_r_55__15_, s_r_55__14_, s_r_55__13_, s_r_55__12_, s_r_55__11_, s_r_55__10_, s_r_55__9_, s_r_55__8_, s_r_55__7_, s_r_55__6_, s_r_55__5_, s_r_55__4_, s_r_55__3_, s_r_55__2_, s_r_55__1_, s_r_55__0_ }),
    .c_o(c_r[55]),
    .prod_accum_o({ prod_accum_55__56_, prod_accum_55__55_, prod_accum_55__54_, prod_accum_55__53_, prod_accum_55__52_, prod_accum_55__51_, prod_accum_55__50_, prod_accum_55__49_, prod_accum_55__48_, prod_accum_55__47_, prod_accum_55__46_, prod_accum_55__45_, prod_accum_55__44_, prod_accum_55__43_, prod_accum_55__42_, prod_accum_55__41_, prod_accum_55__40_, prod_accum_55__39_, prod_accum_55__38_, prod_accum_55__37_, prod_accum_55__36_, prod_accum_55__35_, prod_accum_55__34_, prod_accum_55__33_, prod_accum_55__32_, prod_accum_55__31_, prod_accum_55__30_, prod_accum_55__29_, prod_accum_55__28_, prod_accum_55__27_, prod_accum_55__26_, prod_accum_55__25_, prod_accum_55__24_, prod_accum_55__23_, prod_accum_55__22_, prod_accum_55__21_, prod_accum_55__20_, prod_accum_55__19_, prod_accum_55__18_, prod_accum_55__17_, prod_accum_55__16_, prod_accum_55__15_, prod_accum_55__14_, prod_accum_55__13_, prod_accum_55__12_, prod_accum_55__11_, prod_accum_55__10_, prod_accum_55__9_, prod_accum_55__8_, prod_accum_55__7_, prod_accum_55__6_, prod_accum_55__5_, prod_accum_55__4_, prod_accum_55__3_, prod_accum_55__2_, prod_accum_55__1_, prod_accum_55__0_ })
  );


  bsg_mul_array_row_128_56_x
  genblk1_56__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[7167:7040]),
    .b_i(b_r[7167:7040]),
    .s_i({ s_r_55__127_, s_r_55__126_, s_r_55__125_, s_r_55__124_, s_r_55__123_, s_r_55__122_, s_r_55__121_, s_r_55__120_, s_r_55__119_, s_r_55__118_, s_r_55__117_, s_r_55__116_, s_r_55__115_, s_r_55__114_, s_r_55__113_, s_r_55__112_, s_r_55__111_, s_r_55__110_, s_r_55__109_, s_r_55__108_, s_r_55__107_, s_r_55__106_, s_r_55__105_, s_r_55__104_, s_r_55__103_, s_r_55__102_, s_r_55__101_, s_r_55__100_, s_r_55__99_, s_r_55__98_, s_r_55__97_, s_r_55__96_, s_r_55__95_, s_r_55__94_, s_r_55__93_, s_r_55__92_, s_r_55__91_, s_r_55__90_, s_r_55__89_, s_r_55__88_, s_r_55__87_, s_r_55__86_, s_r_55__85_, s_r_55__84_, s_r_55__83_, s_r_55__82_, s_r_55__81_, s_r_55__80_, s_r_55__79_, s_r_55__78_, s_r_55__77_, s_r_55__76_, s_r_55__75_, s_r_55__74_, s_r_55__73_, s_r_55__72_, s_r_55__71_, s_r_55__70_, s_r_55__69_, s_r_55__68_, s_r_55__67_, s_r_55__66_, s_r_55__65_, s_r_55__64_, s_r_55__63_, s_r_55__62_, s_r_55__61_, s_r_55__60_, s_r_55__59_, s_r_55__58_, s_r_55__57_, s_r_55__56_, s_r_55__55_, s_r_55__54_, s_r_55__53_, s_r_55__52_, s_r_55__51_, s_r_55__50_, s_r_55__49_, s_r_55__48_, s_r_55__47_, s_r_55__46_, s_r_55__45_, s_r_55__44_, s_r_55__43_, s_r_55__42_, s_r_55__41_, s_r_55__40_, s_r_55__39_, s_r_55__38_, s_r_55__37_, s_r_55__36_, s_r_55__35_, s_r_55__34_, s_r_55__33_, s_r_55__32_, s_r_55__31_, s_r_55__30_, s_r_55__29_, s_r_55__28_, s_r_55__27_, s_r_55__26_, s_r_55__25_, s_r_55__24_, s_r_55__23_, s_r_55__22_, s_r_55__21_, s_r_55__20_, s_r_55__19_, s_r_55__18_, s_r_55__17_, s_r_55__16_, s_r_55__15_, s_r_55__14_, s_r_55__13_, s_r_55__12_, s_r_55__11_, s_r_55__10_, s_r_55__9_, s_r_55__8_, s_r_55__7_, s_r_55__6_, s_r_55__5_, s_r_55__4_, s_r_55__3_, s_r_55__2_, s_r_55__1_, s_r_55__0_ }),
    .c_i(c_r[55]),
    .prod_accum_i({ prod_accum_55__56_, prod_accum_55__55_, prod_accum_55__54_, prod_accum_55__53_, prod_accum_55__52_, prod_accum_55__51_, prod_accum_55__50_, prod_accum_55__49_, prod_accum_55__48_, prod_accum_55__47_, prod_accum_55__46_, prod_accum_55__45_, prod_accum_55__44_, prod_accum_55__43_, prod_accum_55__42_, prod_accum_55__41_, prod_accum_55__40_, prod_accum_55__39_, prod_accum_55__38_, prod_accum_55__37_, prod_accum_55__36_, prod_accum_55__35_, prod_accum_55__34_, prod_accum_55__33_, prod_accum_55__32_, prod_accum_55__31_, prod_accum_55__30_, prod_accum_55__29_, prod_accum_55__28_, prod_accum_55__27_, prod_accum_55__26_, prod_accum_55__25_, prod_accum_55__24_, prod_accum_55__23_, prod_accum_55__22_, prod_accum_55__21_, prod_accum_55__20_, prod_accum_55__19_, prod_accum_55__18_, prod_accum_55__17_, prod_accum_55__16_, prod_accum_55__15_, prod_accum_55__14_, prod_accum_55__13_, prod_accum_55__12_, prod_accum_55__11_, prod_accum_55__10_, prod_accum_55__9_, prod_accum_55__8_, prod_accum_55__7_, prod_accum_55__6_, prod_accum_55__5_, prod_accum_55__4_, prod_accum_55__3_, prod_accum_55__2_, prod_accum_55__1_, prod_accum_55__0_ }),
    .a_o(a_r[7295:7168]),
    .b_o(b_r[7295:7168]),
    .s_o({ s_r_56__127_, s_r_56__126_, s_r_56__125_, s_r_56__124_, s_r_56__123_, s_r_56__122_, s_r_56__121_, s_r_56__120_, s_r_56__119_, s_r_56__118_, s_r_56__117_, s_r_56__116_, s_r_56__115_, s_r_56__114_, s_r_56__113_, s_r_56__112_, s_r_56__111_, s_r_56__110_, s_r_56__109_, s_r_56__108_, s_r_56__107_, s_r_56__106_, s_r_56__105_, s_r_56__104_, s_r_56__103_, s_r_56__102_, s_r_56__101_, s_r_56__100_, s_r_56__99_, s_r_56__98_, s_r_56__97_, s_r_56__96_, s_r_56__95_, s_r_56__94_, s_r_56__93_, s_r_56__92_, s_r_56__91_, s_r_56__90_, s_r_56__89_, s_r_56__88_, s_r_56__87_, s_r_56__86_, s_r_56__85_, s_r_56__84_, s_r_56__83_, s_r_56__82_, s_r_56__81_, s_r_56__80_, s_r_56__79_, s_r_56__78_, s_r_56__77_, s_r_56__76_, s_r_56__75_, s_r_56__74_, s_r_56__73_, s_r_56__72_, s_r_56__71_, s_r_56__70_, s_r_56__69_, s_r_56__68_, s_r_56__67_, s_r_56__66_, s_r_56__65_, s_r_56__64_, s_r_56__63_, s_r_56__62_, s_r_56__61_, s_r_56__60_, s_r_56__59_, s_r_56__58_, s_r_56__57_, s_r_56__56_, s_r_56__55_, s_r_56__54_, s_r_56__53_, s_r_56__52_, s_r_56__51_, s_r_56__50_, s_r_56__49_, s_r_56__48_, s_r_56__47_, s_r_56__46_, s_r_56__45_, s_r_56__44_, s_r_56__43_, s_r_56__42_, s_r_56__41_, s_r_56__40_, s_r_56__39_, s_r_56__38_, s_r_56__37_, s_r_56__36_, s_r_56__35_, s_r_56__34_, s_r_56__33_, s_r_56__32_, s_r_56__31_, s_r_56__30_, s_r_56__29_, s_r_56__28_, s_r_56__27_, s_r_56__26_, s_r_56__25_, s_r_56__24_, s_r_56__23_, s_r_56__22_, s_r_56__21_, s_r_56__20_, s_r_56__19_, s_r_56__18_, s_r_56__17_, s_r_56__16_, s_r_56__15_, s_r_56__14_, s_r_56__13_, s_r_56__12_, s_r_56__11_, s_r_56__10_, s_r_56__9_, s_r_56__8_, s_r_56__7_, s_r_56__6_, s_r_56__5_, s_r_56__4_, s_r_56__3_, s_r_56__2_, s_r_56__1_, s_r_56__0_ }),
    .c_o(c_r[56]),
    .prod_accum_o({ prod_accum_56__57_, prod_accum_56__56_, prod_accum_56__55_, prod_accum_56__54_, prod_accum_56__53_, prod_accum_56__52_, prod_accum_56__51_, prod_accum_56__50_, prod_accum_56__49_, prod_accum_56__48_, prod_accum_56__47_, prod_accum_56__46_, prod_accum_56__45_, prod_accum_56__44_, prod_accum_56__43_, prod_accum_56__42_, prod_accum_56__41_, prod_accum_56__40_, prod_accum_56__39_, prod_accum_56__38_, prod_accum_56__37_, prod_accum_56__36_, prod_accum_56__35_, prod_accum_56__34_, prod_accum_56__33_, prod_accum_56__32_, prod_accum_56__31_, prod_accum_56__30_, prod_accum_56__29_, prod_accum_56__28_, prod_accum_56__27_, prod_accum_56__26_, prod_accum_56__25_, prod_accum_56__24_, prod_accum_56__23_, prod_accum_56__22_, prod_accum_56__21_, prod_accum_56__20_, prod_accum_56__19_, prod_accum_56__18_, prod_accum_56__17_, prod_accum_56__16_, prod_accum_56__15_, prod_accum_56__14_, prod_accum_56__13_, prod_accum_56__12_, prod_accum_56__11_, prod_accum_56__10_, prod_accum_56__9_, prod_accum_56__8_, prod_accum_56__7_, prod_accum_56__6_, prod_accum_56__5_, prod_accum_56__4_, prod_accum_56__3_, prod_accum_56__2_, prod_accum_56__1_, prod_accum_56__0_ })
  );


  bsg_mul_array_row_128_57_x
  genblk1_57__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[7295:7168]),
    .b_i(b_r[7295:7168]),
    .s_i({ s_r_56__127_, s_r_56__126_, s_r_56__125_, s_r_56__124_, s_r_56__123_, s_r_56__122_, s_r_56__121_, s_r_56__120_, s_r_56__119_, s_r_56__118_, s_r_56__117_, s_r_56__116_, s_r_56__115_, s_r_56__114_, s_r_56__113_, s_r_56__112_, s_r_56__111_, s_r_56__110_, s_r_56__109_, s_r_56__108_, s_r_56__107_, s_r_56__106_, s_r_56__105_, s_r_56__104_, s_r_56__103_, s_r_56__102_, s_r_56__101_, s_r_56__100_, s_r_56__99_, s_r_56__98_, s_r_56__97_, s_r_56__96_, s_r_56__95_, s_r_56__94_, s_r_56__93_, s_r_56__92_, s_r_56__91_, s_r_56__90_, s_r_56__89_, s_r_56__88_, s_r_56__87_, s_r_56__86_, s_r_56__85_, s_r_56__84_, s_r_56__83_, s_r_56__82_, s_r_56__81_, s_r_56__80_, s_r_56__79_, s_r_56__78_, s_r_56__77_, s_r_56__76_, s_r_56__75_, s_r_56__74_, s_r_56__73_, s_r_56__72_, s_r_56__71_, s_r_56__70_, s_r_56__69_, s_r_56__68_, s_r_56__67_, s_r_56__66_, s_r_56__65_, s_r_56__64_, s_r_56__63_, s_r_56__62_, s_r_56__61_, s_r_56__60_, s_r_56__59_, s_r_56__58_, s_r_56__57_, s_r_56__56_, s_r_56__55_, s_r_56__54_, s_r_56__53_, s_r_56__52_, s_r_56__51_, s_r_56__50_, s_r_56__49_, s_r_56__48_, s_r_56__47_, s_r_56__46_, s_r_56__45_, s_r_56__44_, s_r_56__43_, s_r_56__42_, s_r_56__41_, s_r_56__40_, s_r_56__39_, s_r_56__38_, s_r_56__37_, s_r_56__36_, s_r_56__35_, s_r_56__34_, s_r_56__33_, s_r_56__32_, s_r_56__31_, s_r_56__30_, s_r_56__29_, s_r_56__28_, s_r_56__27_, s_r_56__26_, s_r_56__25_, s_r_56__24_, s_r_56__23_, s_r_56__22_, s_r_56__21_, s_r_56__20_, s_r_56__19_, s_r_56__18_, s_r_56__17_, s_r_56__16_, s_r_56__15_, s_r_56__14_, s_r_56__13_, s_r_56__12_, s_r_56__11_, s_r_56__10_, s_r_56__9_, s_r_56__8_, s_r_56__7_, s_r_56__6_, s_r_56__5_, s_r_56__4_, s_r_56__3_, s_r_56__2_, s_r_56__1_, s_r_56__0_ }),
    .c_i(c_r[56]),
    .prod_accum_i({ prod_accum_56__57_, prod_accum_56__56_, prod_accum_56__55_, prod_accum_56__54_, prod_accum_56__53_, prod_accum_56__52_, prod_accum_56__51_, prod_accum_56__50_, prod_accum_56__49_, prod_accum_56__48_, prod_accum_56__47_, prod_accum_56__46_, prod_accum_56__45_, prod_accum_56__44_, prod_accum_56__43_, prod_accum_56__42_, prod_accum_56__41_, prod_accum_56__40_, prod_accum_56__39_, prod_accum_56__38_, prod_accum_56__37_, prod_accum_56__36_, prod_accum_56__35_, prod_accum_56__34_, prod_accum_56__33_, prod_accum_56__32_, prod_accum_56__31_, prod_accum_56__30_, prod_accum_56__29_, prod_accum_56__28_, prod_accum_56__27_, prod_accum_56__26_, prod_accum_56__25_, prod_accum_56__24_, prod_accum_56__23_, prod_accum_56__22_, prod_accum_56__21_, prod_accum_56__20_, prod_accum_56__19_, prod_accum_56__18_, prod_accum_56__17_, prod_accum_56__16_, prod_accum_56__15_, prod_accum_56__14_, prod_accum_56__13_, prod_accum_56__12_, prod_accum_56__11_, prod_accum_56__10_, prod_accum_56__9_, prod_accum_56__8_, prod_accum_56__7_, prod_accum_56__6_, prod_accum_56__5_, prod_accum_56__4_, prod_accum_56__3_, prod_accum_56__2_, prod_accum_56__1_, prod_accum_56__0_ }),
    .a_o(a_r[7423:7296]),
    .b_o(b_r[7423:7296]),
    .s_o({ s_r_57__127_, s_r_57__126_, s_r_57__125_, s_r_57__124_, s_r_57__123_, s_r_57__122_, s_r_57__121_, s_r_57__120_, s_r_57__119_, s_r_57__118_, s_r_57__117_, s_r_57__116_, s_r_57__115_, s_r_57__114_, s_r_57__113_, s_r_57__112_, s_r_57__111_, s_r_57__110_, s_r_57__109_, s_r_57__108_, s_r_57__107_, s_r_57__106_, s_r_57__105_, s_r_57__104_, s_r_57__103_, s_r_57__102_, s_r_57__101_, s_r_57__100_, s_r_57__99_, s_r_57__98_, s_r_57__97_, s_r_57__96_, s_r_57__95_, s_r_57__94_, s_r_57__93_, s_r_57__92_, s_r_57__91_, s_r_57__90_, s_r_57__89_, s_r_57__88_, s_r_57__87_, s_r_57__86_, s_r_57__85_, s_r_57__84_, s_r_57__83_, s_r_57__82_, s_r_57__81_, s_r_57__80_, s_r_57__79_, s_r_57__78_, s_r_57__77_, s_r_57__76_, s_r_57__75_, s_r_57__74_, s_r_57__73_, s_r_57__72_, s_r_57__71_, s_r_57__70_, s_r_57__69_, s_r_57__68_, s_r_57__67_, s_r_57__66_, s_r_57__65_, s_r_57__64_, s_r_57__63_, s_r_57__62_, s_r_57__61_, s_r_57__60_, s_r_57__59_, s_r_57__58_, s_r_57__57_, s_r_57__56_, s_r_57__55_, s_r_57__54_, s_r_57__53_, s_r_57__52_, s_r_57__51_, s_r_57__50_, s_r_57__49_, s_r_57__48_, s_r_57__47_, s_r_57__46_, s_r_57__45_, s_r_57__44_, s_r_57__43_, s_r_57__42_, s_r_57__41_, s_r_57__40_, s_r_57__39_, s_r_57__38_, s_r_57__37_, s_r_57__36_, s_r_57__35_, s_r_57__34_, s_r_57__33_, s_r_57__32_, s_r_57__31_, s_r_57__30_, s_r_57__29_, s_r_57__28_, s_r_57__27_, s_r_57__26_, s_r_57__25_, s_r_57__24_, s_r_57__23_, s_r_57__22_, s_r_57__21_, s_r_57__20_, s_r_57__19_, s_r_57__18_, s_r_57__17_, s_r_57__16_, s_r_57__15_, s_r_57__14_, s_r_57__13_, s_r_57__12_, s_r_57__11_, s_r_57__10_, s_r_57__9_, s_r_57__8_, s_r_57__7_, s_r_57__6_, s_r_57__5_, s_r_57__4_, s_r_57__3_, s_r_57__2_, s_r_57__1_, s_r_57__0_ }),
    .c_o(c_r[57]),
    .prod_accum_o({ prod_accum_57__58_, prod_accum_57__57_, prod_accum_57__56_, prod_accum_57__55_, prod_accum_57__54_, prod_accum_57__53_, prod_accum_57__52_, prod_accum_57__51_, prod_accum_57__50_, prod_accum_57__49_, prod_accum_57__48_, prod_accum_57__47_, prod_accum_57__46_, prod_accum_57__45_, prod_accum_57__44_, prod_accum_57__43_, prod_accum_57__42_, prod_accum_57__41_, prod_accum_57__40_, prod_accum_57__39_, prod_accum_57__38_, prod_accum_57__37_, prod_accum_57__36_, prod_accum_57__35_, prod_accum_57__34_, prod_accum_57__33_, prod_accum_57__32_, prod_accum_57__31_, prod_accum_57__30_, prod_accum_57__29_, prod_accum_57__28_, prod_accum_57__27_, prod_accum_57__26_, prod_accum_57__25_, prod_accum_57__24_, prod_accum_57__23_, prod_accum_57__22_, prod_accum_57__21_, prod_accum_57__20_, prod_accum_57__19_, prod_accum_57__18_, prod_accum_57__17_, prod_accum_57__16_, prod_accum_57__15_, prod_accum_57__14_, prod_accum_57__13_, prod_accum_57__12_, prod_accum_57__11_, prod_accum_57__10_, prod_accum_57__9_, prod_accum_57__8_, prod_accum_57__7_, prod_accum_57__6_, prod_accum_57__5_, prod_accum_57__4_, prod_accum_57__3_, prod_accum_57__2_, prod_accum_57__1_, prod_accum_57__0_ })
  );


  bsg_mul_array_row_128_58_x
  genblk1_58__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[7423:7296]),
    .b_i(b_r[7423:7296]),
    .s_i({ s_r_57__127_, s_r_57__126_, s_r_57__125_, s_r_57__124_, s_r_57__123_, s_r_57__122_, s_r_57__121_, s_r_57__120_, s_r_57__119_, s_r_57__118_, s_r_57__117_, s_r_57__116_, s_r_57__115_, s_r_57__114_, s_r_57__113_, s_r_57__112_, s_r_57__111_, s_r_57__110_, s_r_57__109_, s_r_57__108_, s_r_57__107_, s_r_57__106_, s_r_57__105_, s_r_57__104_, s_r_57__103_, s_r_57__102_, s_r_57__101_, s_r_57__100_, s_r_57__99_, s_r_57__98_, s_r_57__97_, s_r_57__96_, s_r_57__95_, s_r_57__94_, s_r_57__93_, s_r_57__92_, s_r_57__91_, s_r_57__90_, s_r_57__89_, s_r_57__88_, s_r_57__87_, s_r_57__86_, s_r_57__85_, s_r_57__84_, s_r_57__83_, s_r_57__82_, s_r_57__81_, s_r_57__80_, s_r_57__79_, s_r_57__78_, s_r_57__77_, s_r_57__76_, s_r_57__75_, s_r_57__74_, s_r_57__73_, s_r_57__72_, s_r_57__71_, s_r_57__70_, s_r_57__69_, s_r_57__68_, s_r_57__67_, s_r_57__66_, s_r_57__65_, s_r_57__64_, s_r_57__63_, s_r_57__62_, s_r_57__61_, s_r_57__60_, s_r_57__59_, s_r_57__58_, s_r_57__57_, s_r_57__56_, s_r_57__55_, s_r_57__54_, s_r_57__53_, s_r_57__52_, s_r_57__51_, s_r_57__50_, s_r_57__49_, s_r_57__48_, s_r_57__47_, s_r_57__46_, s_r_57__45_, s_r_57__44_, s_r_57__43_, s_r_57__42_, s_r_57__41_, s_r_57__40_, s_r_57__39_, s_r_57__38_, s_r_57__37_, s_r_57__36_, s_r_57__35_, s_r_57__34_, s_r_57__33_, s_r_57__32_, s_r_57__31_, s_r_57__30_, s_r_57__29_, s_r_57__28_, s_r_57__27_, s_r_57__26_, s_r_57__25_, s_r_57__24_, s_r_57__23_, s_r_57__22_, s_r_57__21_, s_r_57__20_, s_r_57__19_, s_r_57__18_, s_r_57__17_, s_r_57__16_, s_r_57__15_, s_r_57__14_, s_r_57__13_, s_r_57__12_, s_r_57__11_, s_r_57__10_, s_r_57__9_, s_r_57__8_, s_r_57__7_, s_r_57__6_, s_r_57__5_, s_r_57__4_, s_r_57__3_, s_r_57__2_, s_r_57__1_, s_r_57__0_ }),
    .c_i(c_r[57]),
    .prod_accum_i({ prod_accum_57__58_, prod_accum_57__57_, prod_accum_57__56_, prod_accum_57__55_, prod_accum_57__54_, prod_accum_57__53_, prod_accum_57__52_, prod_accum_57__51_, prod_accum_57__50_, prod_accum_57__49_, prod_accum_57__48_, prod_accum_57__47_, prod_accum_57__46_, prod_accum_57__45_, prod_accum_57__44_, prod_accum_57__43_, prod_accum_57__42_, prod_accum_57__41_, prod_accum_57__40_, prod_accum_57__39_, prod_accum_57__38_, prod_accum_57__37_, prod_accum_57__36_, prod_accum_57__35_, prod_accum_57__34_, prod_accum_57__33_, prod_accum_57__32_, prod_accum_57__31_, prod_accum_57__30_, prod_accum_57__29_, prod_accum_57__28_, prod_accum_57__27_, prod_accum_57__26_, prod_accum_57__25_, prod_accum_57__24_, prod_accum_57__23_, prod_accum_57__22_, prod_accum_57__21_, prod_accum_57__20_, prod_accum_57__19_, prod_accum_57__18_, prod_accum_57__17_, prod_accum_57__16_, prod_accum_57__15_, prod_accum_57__14_, prod_accum_57__13_, prod_accum_57__12_, prod_accum_57__11_, prod_accum_57__10_, prod_accum_57__9_, prod_accum_57__8_, prod_accum_57__7_, prod_accum_57__6_, prod_accum_57__5_, prod_accum_57__4_, prod_accum_57__3_, prod_accum_57__2_, prod_accum_57__1_, prod_accum_57__0_ }),
    .a_o(a_r[7551:7424]),
    .b_o(b_r[7551:7424]),
    .s_o({ s_r_58__127_, s_r_58__126_, s_r_58__125_, s_r_58__124_, s_r_58__123_, s_r_58__122_, s_r_58__121_, s_r_58__120_, s_r_58__119_, s_r_58__118_, s_r_58__117_, s_r_58__116_, s_r_58__115_, s_r_58__114_, s_r_58__113_, s_r_58__112_, s_r_58__111_, s_r_58__110_, s_r_58__109_, s_r_58__108_, s_r_58__107_, s_r_58__106_, s_r_58__105_, s_r_58__104_, s_r_58__103_, s_r_58__102_, s_r_58__101_, s_r_58__100_, s_r_58__99_, s_r_58__98_, s_r_58__97_, s_r_58__96_, s_r_58__95_, s_r_58__94_, s_r_58__93_, s_r_58__92_, s_r_58__91_, s_r_58__90_, s_r_58__89_, s_r_58__88_, s_r_58__87_, s_r_58__86_, s_r_58__85_, s_r_58__84_, s_r_58__83_, s_r_58__82_, s_r_58__81_, s_r_58__80_, s_r_58__79_, s_r_58__78_, s_r_58__77_, s_r_58__76_, s_r_58__75_, s_r_58__74_, s_r_58__73_, s_r_58__72_, s_r_58__71_, s_r_58__70_, s_r_58__69_, s_r_58__68_, s_r_58__67_, s_r_58__66_, s_r_58__65_, s_r_58__64_, s_r_58__63_, s_r_58__62_, s_r_58__61_, s_r_58__60_, s_r_58__59_, s_r_58__58_, s_r_58__57_, s_r_58__56_, s_r_58__55_, s_r_58__54_, s_r_58__53_, s_r_58__52_, s_r_58__51_, s_r_58__50_, s_r_58__49_, s_r_58__48_, s_r_58__47_, s_r_58__46_, s_r_58__45_, s_r_58__44_, s_r_58__43_, s_r_58__42_, s_r_58__41_, s_r_58__40_, s_r_58__39_, s_r_58__38_, s_r_58__37_, s_r_58__36_, s_r_58__35_, s_r_58__34_, s_r_58__33_, s_r_58__32_, s_r_58__31_, s_r_58__30_, s_r_58__29_, s_r_58__28_, s_r_58__27_, s_r_58__26_, s_r_58__25_, s_r_58__24_, s_r_58__23_, s_r_58__22_, s_r_58__21_, s_r_58__20_, s_r_58__19_, s_r_58__18_, s_r_58__17_, s_r_58__16_, s_r_58__15_, s_r_58__14_, s_r_58__13_, s_r_58__12_, s_r_58__11_, s_r_58__10_, s_r_58__9_, s_r_58__8_, s_r_58__7_, s_r_58__6_, s_r_58__5_, s_r_58__4_, s_r_58__3_, s_r_58__2_, s_r_58__1_, s_r_58__0_ }),
    .c_o(c_r[58]),
    .prod_accum_o({ prod_accum_58__59_, prod_accum_58__58_, prod_accum_58__57_, prod_accum_58__56_, prod_accum_58__55_, prod_accum_58__54_, prod_accum_58__53_, prod_accum_58__52_, prod_accum_58__51_, prod_accum_58__50_, prod_accum_58__49_, prod_accum_58__48_, prod_accum_58__47_, prod_accum_58__46_, prod_accum_58__45_, prod_accum_58__44_, prod_accum_58__43_, prod_accum_58__42_, prod_accum_58__41_, prod_accum_58__40_, prod_accum_58__39_, prod_accum_58__38_, prod_accum_58__37_, prod_accum_58__36_, prod_accum_58__35_, prod_accum_58__34_, prod_accum_58__33_, prod_accum_58__32_, prod_accum_58__31_, prod_accum_58__30_, prod_accum_58__29_, prod_accum_58__28_, prod_accum_58__27_, prod_accum_58__26_, prod_accum_58__25_, prod_accum_58__24_, prod_accum_58__23_, prod_accum_58__22_, prod_accum_58__21_, prod_accum_58__20_, prod_accum_58__19_, prod_accum_58__18_, prod_accum_58__17_, prod_accum_58__16_, prod_accum_58__15_, prod_accum_58__14_, prod_accum_58__13_, prod_accum_58__12_, prod_accum_58__11_, prod_accum_58__10_, prod_accum_58__9_, prod_accum_58__8_, prod_accum_58__7_, prod_accum_58__6_, prod_accum_58__5_, prod_accum_58__4_, prod_accum_58__3_, prod_accum_58__2_, prod_accum_58__1_, prod_accum_58__0_ })
  );


  bsg_mul_array_row_128_59_x
  genblk1_59__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[7551:7424]),
    .b_i(b_r[7551:7424]),
    .s_i({ s_r_58__127_, s_r_58__126_, s_r_58__125_, s_r_58__124_, s_r_58__123_, s_r_58__122_, s_r_58__121_, s_r_58__120_, s_r_58__119_, s_r_58__118_, s_r_58__117_, s_r_58__116_, s_r_58__115_, s_r_58__114_, s_r_58__113_, s_r_58__112_, s_r_58__111_, s_r_58__110_, s_r_58__109_, s_r_58__108_, s_r_58__107_, s_r_58__106_, s_r_58__105_, s_r_58__104_, s_r_58__103_, s_r_58__102_, s_r_58__101_, s_r_58__100_, s_r_58__99_, s_r_58__98_, s_r_58__97_, s_r_58__96_, s_r_58__95_, s_r_58__94_, s_r_58__93_, s_r_58__92_, s_r_58__91_, s_r_58__90_, s_r_58__89_, s_r_58__88_, s_r_58__87_, s_r_58__86_, s_r_58__85_, s_r_58__84_, s_r_58__83_, s_r_58__82_, s_r_58__81_, s_r_58__80_, s_r_58__79_, s_r_58__78_, s_r_58__77_, s_r_58__76_, s_r_58__75_, s_r_58__74_, s_r_58__73_, s_r_58__72_, s_r_58__71_, s_r_58__70_, s_r_58__69_, s_r_58__68_, s_r_58__67_, s_r_58__66_, s_r_58__65_, s_r_58__64_, s_r_58__63_, s_r_58__62_, s_r_58__61_, s_r_58__60_, s_r_58__59_, s_r_58__58_, s_r_58__57_, s_r_58__56_, s_r_58__55_, s_r_58__54_, s_r_58__53_, s_r_58__52_, s_r_58__51_, s_r_58__50_, s_r_58__49_, s_r_58__48_, s_r_58__47_, s_r_58__46_, s_r_58__45_, s_r_58__44_, s_r_58__43_, s_r_58__42_, s_r_58__41_, s_r_58__40_, s_r_58__39_, s_r_58__38_, s_r_58__37_, s_r_58__36_, s_r_58__35_, s_r_58__34_, s_r_58__33_, s_r_58__32_, s_r_58__31_, s_r_58__30_, s_r_58__29_, s_r_58__28_, s_r_58__27_, s_r_58__26_, s_r_58__25_, s_r_58__24_, s_r_58__23_, s_r_58__22_, s_r_58__21_, s_r_58__20_, s_r_58__19_, s_r_58__18_, s_r_58__17_, s_r_58__16_, s_r_58__15_, s_r_58__14_, s_r_58__13_, s_r_58__12_, s_r_58__11_, s_r_58__10_, s_r_58__9_, s_r_58__8_, s_r_58__7_, s_r_58__6_, s_r_58__5_, s_r_58__4_, s_r_58__3_, s_r_58__2_, s_r_58__1_, s_r_58__0_ }),
    .c_i(c_r[58]),
    .prod_accum_i({ prod_accum_58__59_, prod_accum_58__58_, prod_accum_58__57_, prod_accum_58__56_, prod_accum_58__55_, prod_accum_58__54_, prod_accum_58__53_, prod_accum_58__52_, prod_accum_58__51_, prod_accum_58__50_, prod_accum_58__49_, prod_accum_58__48_, prod_accum_58__47_, prod_accum_58__46_, prod_accum_58__45_, prod_accum_58__44_, prod_accum_58__43_, prod_accum_58__42_, prod_accum_58__41_, prod_accum_58__40_, prod_accum_58__39_, prod_accum_58__38_, prod_accum_58__37_, prod_accum_58__36_, prod_accum_58__35_, prod_accum_58__34_, prod_accum_58__33_, prod_accum_58__32_, prod_accum_58__31_, prod_accum_58__30_, prod_accum_58__29_, prod_accum_58__28_, prod_accum_58__27_, prod_accum_58__26_, prod_accum_58__25_, prod_accum_58__24_, prod_accum_58__23_, prod_accum_58__22_, prod_accum_58__21_, prod_accum_58__20_, prod_accum_58__19_, prod_accum_58__18_, prod_accum_58__17_, prod_accum_58__16_, prod_accum_58__15_, prod_accum_58__14_, prod_accum_58__13_, prod_accum_58__12_, prod_accum_58__11_, prod_accum_58__10_, prod_accum_58__9_, prod_accum_58__8_, prod_accum_58__7_, prod_accum_58__6_, prod_accum_58__5_, prod_accum_58__4_, prod_accum_58__3_, prod_accum_58__2_, prod_accum_58__1_, prod_accum_58__0_ }),
    .a_o(a_r[7679:7552]),
    .b_o(b_r[7679:7552]),
    .s_o({ s_r_59__127_, s_r_59__126_, s_r_59__125_, s_r_59__124_, s_r_59__123_, s_r_59__122_, s_r_59__121_, s_r_59__120_, s_r_59__119_, s_r_59__118_, s_r_59__117_, s_r_59__116_, s_r_59__115_, s_r_59__114_, s_r_59__113_, s_r_59__112_, s_r_59__111_, s_r_59__110_, s_r_59__109_, s_r_59__108_, s_r_59__107_, s_r_59__106_, s_r_59__105_, s_r_59__104_, s_r_59__103_, s_r_59__102_, s_r_59__101_, s_r_59__100_, s_r_59__99_, s_r_59__98_, s_r_59__97_, s_r_59__96_, s_r_59__95_, s_r_59__94_, s_r_59__93_, s_r_59__92_, s_r_59__91_, s_r_59__90_, s_r_59__89_, s_r_59__88_, s_r_59__87_, s_r_59__86_, s_r_59__85_, s_r_59__84_, s_r_59__83_, s_r_59__82_, s_r_59__81_, s_r_59__80_, s_r_59__79_, s_r_59__78_, s_r_59__77_, s_r_59__76_, s_r_59__75_, s_r_59__74_, s_r_59__73_, s_r_59__72_, s_r_59__71_, s_r_59__70_, s_r_59__69_, s_r_59__68_, s_r_59__67_, s_r_59__66_, s_r_59__65_, s_r_59__64_, s_r_59__63_, s_r_59__62_, s_r_59__61_, s_r_59__60_, s_r_59__59_, s_r_59__58_, s_r_59__57_, s_r_59__56_, s_r_59__55_, s_r_59__54_, s_r_59__53_, s_r_59__52_, s_r_59__51_, s_r_59__50_, s_r_59__49_, s_r_59__48_, s_r_59__47_, s_r_59__46_, s_r_59__45_, s_r_59__44_, s_r_59__43_, s_r_59__42_, s_r_59__41_, s_r_59__40_, s_r_59__39_, s_r_59__38_, s_r_59__37_, s_r_59__36_, s_r_59__35_, s_r_59__34_, s_r_59__33_, s_r_59__32_, s_r_59__31_, s_r_59__30_, s_r_59__29_, s_r_59__28_, s_r_59__27_, s_r_59__26_, s_r_59__25_, s_r_59__24_, s_r_59__23_, s_r_59__22_, s_r_59__21_, s_r_59__20_, s_r_59__19_, s_r_59__18_, s_r_59__17_, s_r_59__16_, s_r_59__15_, s_r_59__14_, s_r_59__13_, s_r_59__12_, s_r_59__11_, s_r_59__10_, s_r_59__9_, s_r_59__8_, s_r_59__7_, s_r_59__6_, s_r_59__5_, s_r_59__4_, s_r_59__3_, s_r_59__2_, s_r_59__1_, s_r_59__0_ }),
    .c_o(c_r[59]),
    .prod_accum_o({ prod_accum_59__60_, prod_accum_59__59_, prod_accum_59__58_, prod_accum_59__57_, prod_accum_59__56_, prod_accum_59__55_, prod_accum_59__54_, prod_accum_59__53_, prod_accum_59__52_, prod_accum_59__51_, prod_accum_59__50_, prod_accum_59__49_, prod_accum_59__48_, prod_accum_59__47_, prod_accum_59__46_, prod_accum_59__45_, prod_accum_59__44_, prod_accum_59__43_, prod_accum_59__42_, prod_accum_59__41_, prod_accum_59__40_, prod_accum_59__39_, prod_accum_59__38_, prod_accum_59__37_, prod_accum_59__36_, prod_accum_59__35_, prod_accum_59__34_, prod_accum_59__33_, prod_accum_59__32_, prod_accum_59__31_, prod_accum_59__30_, prod_accum_59__29_, prod_accum_59__28_, prod_accum_59__27_, prod_accum_59__26_, prod_accum_59__25_, prod_accum_59__24_, prod_accum_59__23_, prod_accum_59__22_, prod_accum_59__21_, prod_accum_59__20_, prod_accum_59__19_, prod_accum_59__18_, prod_accum_59__17_, prod_accum_59__16_, prod_accum_59__15_, prod_accum_59__14_, prod_accum_59__13_, prod_accum_59__12_, prod_accum_59__11_, prod_accum_59__10_, prod_accum_59__9_, prod_accum_59__8_, prod_accum_59__7_, prod_accum_59__6_, prod_accum_59__5_, prod_accum_59__4_, prod_accum_59__3_, prod_accum_59__2_, prod_accum_59__1_, prod_accum_59__0_ })
  );


  bsg_mul_array_row_128_60_x
  genblk1_60__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[7679:7552]),
    .b_i(b_r[7679:7552]),
    .s_i({ s_r_59__127_, s_r_59__126_, s_r_59__125_, s_r_59__124_, s_r_59__123_, s_r_59__122_, s_r_59__121_, s_r_59__120_, s_r_59__119_, s_r_59__118_, s_r_59__117_, s_r_59__116_, s_r_59__115_, s_r_59__114_, s_r_59__113_, s_r_59__112_, s_r_59__111_, s_r_59__110_, s_r_59__109_, s_r_59__108_, s_r_59__107_, s_r_59__106_, s_r_59__105_, s_r_59__104_, s_r_59__103_, s_r_59__102_, s_r_59__101_, s_r_59__100_, s_r_59__99_, s_r_59__98_, s_r_59__97_, s_r_59__96_, s_r_59__95_, s_r_59__94_, s_r_59__93_, s_r_59__92_, s_r_59__91_, s_r_59__90_, s_r_59__89_, s_r_59__88_, s_r_59__87_, s_r_59__86_, s_r_59__85_, s_r_59__84_, s_r_59__83_, s_r_59__82_, s_r_59__81_, s_r_59__80_, s_r_59__79_, s_r_59__78_, s_r_59__77_, s_r_59__76_, s_r_59__75_, s_r_59__74_, s_r_59__73_, s_r_59__72_, s_r_59__71_, s_r_59__70_, s_r_59__69_, s_r_59__68_, s_r_59__67_, s_r_59__66_, s_r_59__65_, s_r_59__64_, s_r_59__63_, s_r_59__62_, s_r_59__61_, s_r_59__60_, s_r_59__59_, s_r_59__58_, s_r_59__57_, s_r_59__56_, s_r_59__55_, s_r_59__54_, s_r_59__53_, s_r_59__52_, s_r_59__51_, s_r_59__50_, s_r_59__49_, s_r_59__48_, s_r_59__47_, s_r_59__46_, s_r_59__45_, s_r_59__44_, s_r_59__43_, s_r_59__42_, s_r_59__41_, s_r_59__40_, s_r_59__39_, s_r_59__38_, s_r_59__37_, s_r_59__36_, s_r_59__35_, s_r_59__34_, s_r_59__33_, s_r_59__32_, s_r_59__31_, s_r_59__30_, s_r_59__29_, s_r_59__28_, s_r_59__27_, s_r_59__26_, s_r_59__25_, s_r_59__24_, s_r_59__23_, s_r_59__22_, s_r_59__21_, s_r_59__20_, s_r_59__19_, s_r_59__18_, s_r_59__17_, s_r_59__16_, s_r_59__15_, s_r_59__14_, s_r_59__13_, s_r_59__12_, s_r_59__11_, s_r_59__10_, s_r_59__9_, s_r_59__8_, s_r_59__7_, s_r_59__6_, s_r_59__5_, s_r_59__4_, s_r_59__3_, s_r_59__2_, s_r_59__1_, s_r_59__0_ }),
    .c_i(c_r[59]),
    .prod_accum_i({ prod_accum_59__60_, prod_accum_59__59_, prod_accum_59__58_, prod_accum_59__57_, prod_accum_59__56_, prod_accum_59__55_, prod_accum_59__54_, prod_accum_59__53_, prod_accum_59__52_, prod_accum_59__51_, prod_accum_59__50_, prod_accum_59__49_, prod_accum_59__48_, prod_accum_59__47_, prod_accum_59__46_, prod_accum_59__45_, prod_accum_59__44_, prod_accum_59__43_, prod_accum_59__42_, prod_accum_59__41_, prod_accum_59__40_, prod_accum_59__39_, prod_accum_59__38_, prod_accum_59__37_, prod_accum_59__36_, prod_accum_59__35_, prod_accum_59__34_, prod_accum_59__33_, prod_accum_59__32_, prod_accum_59__31_, prod_accum_59__30_, prod_accum_59__29_, prod_accum_59__28_, prod_accum_59__27_, prod_accum_59__26_, prod_accum_59__25_, prod_accum_59__24_, prod_accum_59__23_, prod_accum_59__22_, prod_accum_59__21_, prod_accum_59__20_, prod_accum_59__19_, prod_accum_59__18_, prod_accum_59__17_, prod_accum_59__16_, prod_accum_59__15_, prod_accum_59__14_, prod_accum_59__13_, prod_accum_59__12_, prod_accum_59__11_, prod_accum_59__10_, prod_accum_59__9_, prod_accum_59__8_, prod_accum_59__7_, prod_accum_59__6_, prod_accum_59__5_, prod_accum_59__4_, prod_accum_59__3_, prod_accum_59__2_, prod_accum_59__1_, prod_accum_59__0_ }),
    .a_o(a_r[7807:7680]),
    .b_o(b_r[7807:7680]),
    .s_o({ s_r_60__127_, s_r_60__126_, s_r_60__125_, s_r_60__124_, s_r_60__123_, s_r_60__122_, s_r_60__121_, s_r_60__120_, s_r_60__119_, s_r_60__118_, s_r_60__117_, s_r_60__116_, s_r_60__115_, s_r_60__114_, s_r_60__113_, s_r_60__112_, s_r_60__111_, s_r_60__110_, s_r_60__109_, s_r_60__108_, s_r_60__107_, s_r_60__106_, s_r_60__105_, s_r_60__104_, s_r_60__103_, s_r_60__102_, s_r_60__101_, s_r_60__100_, s_r_60__99_, s_r_60__98_, s_r_60__97_, s_r_60__96_, s_r_60__95_, s_r_60__94_, s_r_60__93_, s_r_60__92_, s_r_60__91_, s_r_60__90_, s_r_60__89_, s_r_60__88_, s_r_60__87_, s_r_60__86_, s_r_60__85_, s_r_60__84_, s_r_60__83_, s_r_60__82_, s_r_60__81_, s_r_60__80_, s_r_60__79_, s_r_60__78_, s_r_60__77_, s_r_60__76_, s_r_60__75_, s_r_60__74_, s_r_60__73_, s_r_60__72_, s_r_60__71_, s_r_60__70_, s_r_60__69_, s_r_60__68_, s_r_60__67_, s_r_60__66_, s_r_60__65_, s_r_60__64_, s_r_60__63_, s_r_60__62_, s_r_60__61_, s_r_60__60_, s_r_60__59_, s_r_60__58_, s_r_60__57_, s_r_60__56_, s_r_60__55_, s_r_60__54_, s_r_60__53_, s_r_60__52_, s_r_60__51_, s_r_60__50_, s_r_60__49_, s_r_60__48_, s_r_60__47_, s_r_60__46_, s_r_60__45_, s_r_60__44_, s_r_60__43_, s_r_60__42_, s_r_60__41_, s_r_60__40_, s_r_60__39_, s_r_60__38_, s_r_60__37_, s_r_60__36_, s_r_60__35_, s_r_60__34_, s_r_60__33_, s_r_60__32_, s_r_60__31_, s_r_60__30_, s_r_60__29_, s_r_60__28_, s_r_60__27_, s_r_60__26_, s_r_60__25_, s_r_60__24_, s_r_60__23_, s_r_60__22_, s_r_60__21_, s_r_60__20_, s_r_60__19_, s_r_60__18_, s_r_60__17_, s_r_60__16_, s_r_60__15_, s_r_60__14_, s_r_60__13_, s_r_60__12_, s_r_60__11_, s_r_60__10_, s_r_60__9_, s_r_60__8_, s_r_60__7_, s_r_60__6_, s_r_60__5_, s_r_60__4_, s_r_60__3_, s_r_60__2_, s_r_60__1_, s_r_60__0_ }),
    .c_o(c_r[60]),
    .prod_accum_o({ prod_accum_60__61_, prod_accum_60__60_, prod_accum_60__59_, prod_accum_60__58_, prod_accum_60__57_, prod_accum_60__56_, prod_accum_60__55_, prod_accum_60__54_, prod_accum_60__53_, prod_accum_60__52_, prod_accum_60__51_, prod_accum_60__50_, prod_accum_60__49_, prod_accum_60__48_, prod_accum_60__47_, prod_accum_60__46_, prod_accum_60__45_, prod_accum_60__44_, prod_accum_60__43_, prod_accum_60__42_, prod_accum_60__41_, prod_accum_60__40_, prod_accum_60__39_, prod_accum_60__38_, prod_accum_60__37_, prod_accum_60__36_, prod_accum_60__35_, prod_accum_60__34_, prod_accum_60__33_, prod_accum_60__32_, prod_accum_60__31_, prod_accum_60__30_, prod_accum_60__29_, prod_accum_60__28_, prod_accum_60__27_, prod_accum_60__26_, prod_accum_60__25_, prod_accum_60__24_, prod_accum_60__23_, prod_accum_60__22_, prod_accum_60__21_, prod_accum_60__20_, prod_accum_60__19_, prod_accum_60__18_, prod_accum_60__17_, prod_accum_60__16_, prod_accum_60__15_, prod_accum_60__14_, prod_accum_60__13_, prod_accum_60__12_, prod_accum_60__11_, prod_accum_60__10_, prod_accum_60__9_, prod_accum_60__8_, prod_accum_60__7_, prod_accum_60__6_, prod_accum_60__5_, prod_accum_60__4_, prod_accum_60__3_, prod_accum_60__2_, prod_accum_60__1_, prod_accum_60__0_ })
  );


  bsg_mul_array_row_128_61_x
  genblk1_61__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[7807:7680]),
    .b_i(b_r[7807:7680]),
    .s_i({ s_r_60__127_, s_r_60__126_, s_r_60__125_, s_r_60__124_, s_r_60__123_, s_r_60__122_, s_r_60__121_, s_r_60__120_, s_r_60__119_, s_r_60__118_, s_r_60__117_, s_r_60__116_, s_r_60__115_, s_r_60__114_, s_r_60__113_, s_r_60__112_, s_r_60__111_, s_r_60__110_, s_r_60__109_, s_r_60__108_, s_r_60__107_, s_r_60__106_, s_r_60__105_, s_r_60__104_, s_r_60__103_, s_r_60__102_, s_r_60__101_, s_r_60__100_, s_r_60__99_, s_r_60__98_, s_r_60__97_, s_r_60__96_, s_r_60__95_, s_r_60__94_, s_r_60__93_, s_r_60__92_, s_r_60__91_, s_r_60__90_, s_r_60__89_, s_r_60__88_, s_r_60__87_, s_r_60__86_, s_r_60__85_, s_r_60__84_, s_r_60__83_, s_r_60__82_, s_r_60__81_, s_r_60__80_, s_r_60__79_, s_r_60__78_, s_r_60__77_, s_r_60__76_, s_r_60__75_, s_r_60__74_, s_r_60__73_, s_r_60__72_, s_r_60__71_, s_r_60__70_, s_r_60__69_, s_r_60__68_, s_r_60__67_, s_r_60__66_, s_r_60__65_, s_r_60__64_, s_r_60__63_, s_r_60__62_, s_r_60__61_, s_r_60__60_, s_r_60__59_, s_r_60__58_, s_r_60__57_, s_r_60__56_, s_r_60__55_, s_r_60__54_, s_r_60__53_, s_r_60__52_, s_r_60__51_, s_r_60__50_, s_r_60__49_, s_r_60__48_, s_r_60__47_, s_r_60__46_, s_r_60__45_, s_r_60__44_, s_r_60__43_, s_r_60__42_, s_r_60__41_, s_r_60__40_, s_r_60__39_, s_r_60__38_, s_r_60__37_, s_r_60__36_, s_r_60__35_, s_r_60__34_, s_r_60__33_, s_r_60__32_, s_r_60__31_, s_r_60__30_, s_r_60__29_, s_r_60__28_, s_r_60__27_, s_r_60__26_, s_r_60__25_, s_r_60__24_, s_r_60__23_, s_r_60__22_, s_r_60__21_, s_r_60__20_, s_r_60__19_, s_r_60__18_, s_r_60__17_, s_r_60__16_, s_r_60__15_, s_r_60__14_, s_r_60__13_, s_r_60__12_, s_r_60__11_, s_r_60__10_, s_r_60__9_, s_r_60__8_, s_r_60__7_, s_r_60__6_, s_r_60__5_, s_r_60__4_, s_r_60__3_, s_r_60__2_, s_r_60__1_, s_r_60__0_ }),
    .c_i(c_r[60]),
    .prod_accum_i({ prod_accum_60__61_, prod_accum_60__60_, prod_accum_60__59_, prod_accum_60__58_, prod_accum_60__57_, prod_accum_60__56_, prod_accum_60__55_, prod_accum_60__54_, prod_accum_60__53_, prod_accum_60__52_, prod_accum_60__51_, prod_accum_60__50_, prod_accum_60__49_, prod_accum_60__48_, prod_accum_60__47_, prod_accum_60__46_, prod_accum_60__45_, prod_accum_60__44_, prod_accum_60__43_, prod_accum_60__42_, prod_accum_60__41_, prod_accum_60__40_, prod_accum_60__39_, prod_accum_60__38_, prod_accum_60__37_, prod_accum_60__36_, prod_accum_60__35_, prod_accum_60__34_, prod_accum_60__33_, prod_accum_60__32_, prod_accum_60__31_, prod_accum_60__30_, prod_accum_60__29_, prod_accum_60__28_, prod_accum_60__27_, prod_accum_60__26_, prod_accum_60__25_, prod_accum_60__24_, prod_accum_60__23_, prod_accum_60__22_, prod_accum_60__21_, prod_accum_60__20_, prod_accum_60__19_, prod_accum_60__18_, prod_accum_60__17_, prod_accum_60__16_, prod_accum_60__15_, prod_accum_60__14_, prod_accum_60__13_, prod_accum_60__12_, prod_accum_60__11_, prod_accum_60__10_, prod_accum_60__9_, prod_accum_60__8_, prod_accum_60__7_, prod_accum_60__6_, prod_accum_60__5_, prod_accum_60__4_, prod_accum_60__3_, prod_accum_60__2_, prod_accum_60__1_, prod_accum_60__0_ }),
    .a_o(a_r[7935:7808]),
    .b_o(b_r[7935:7808]),
    .s_o({ s_r_61__127_, s_r_61__126_, s_r_61__125_, s_r_61__124_, s_r_61__123_, s_r_61__122_, s_r_61__121_, s_r_61__120_, s_r_61__119_, s_r_61__118_, s_r_61__117_, s_r_61__116_, s_r_61__115_, s_r_61__114_, s_r_61__113_, s_r_61__112_, s_r_61__111_, s_r_61__110_, s_r_61__109_, s_r_61__108_, s_r_61__107_, s_r_61__106_, s_r_61__105_, s_r_61__104_, s_r_61__103_, s_r_61__102_, s_r_61__101_, s_r_61__100_, s_r_61__99_, s_r_61__98_, s_r_61__97_, s_r_61__96_, s_r_61__95_, s_r_61__94_, s_r_61__93_, s_r_61__92_, s_r_61__91_, s_r_61__90_, s_r_61__89_, s_r_61__88_, s_r_61__87_, s_r_61__86_, s_r_61__85_, s_r_61__84_, s_r_61__83_, s_r_61__82_, s_r_61__81_, s_r_61__80_, s_r_61__79_, s_r_61__78_, s_r_61__77_, s_r_61__76_, s_r_61__75_, s_r_61__74_, s_r_61__73_, s_r_61__72_, s_r_61__71_, s_r_61__70_, s_r_61__69_, s_r_61__68_, s_r_61__67_, s_r_61__66_, s_r_61__65_, s_r_61__64_, s_r_61__63_, s_r_61__62_, s_r_61__61_, s_r_61__60_, s_r_61__59_, s_r_61__58_, s_r_61__57_, s_r_61__56_, s_r_61__55_, s_r_61__54_, s_r_61__53_, s_r_61__52_, s_r_61__51_, s_r_61__50_, s_r_61__49_, s_r_61__48_, s_r_61__47_, s_r_61__46_, s_r_61__45_, s_r_61__44_, s_r_61__43_, s_r_61__42_, s_r_61__41_, s_r_61__40_, s_r_61__39_, s_r_61__38_, s_r_61__37_, s_r_61__36_, s_r_61__35_, s_r_61__34_, s_r_61__33_, s_r_61__32_, s_r_61__31_, s_r_61__30_, s_r_61__29_, s_r_61__28_, s_r_61__27_, s_r_61__26_, s_r_61__25_, s_r_61__24_, s_r_61__23_, s_r_61__22_, s_r_61__21_, s_r_61__20_, s_r_61__19_, s_r_61__18_, s_r_61__17_, s_r_61__16_, s_r_61__15_, s_r_61__14_, s_r_61__13_, s_r_61__12_, s_r_61__11_, s_r_61__10_, s_r_61__9_, s_r_61__8_, s_r_61__7_, s_r_61__6_, s_r_61__5_, s_r_61__4_, s_r_61__3_, s_r_61__2_, s_r_61__1_, s_r_61__0_ }),
    .c_o(c_r[61]),
    .prod_accum_o({ prod_accum_61__62_, prod_accum_61__61_, prod_accum_61__60_, prod_accum_61__59_, prod_accum_61__58_, prod_accum_61__57_, prod_accum_61__56_, prod_accum_61__55_, prod_accum_61__54_, prod_accum_61__53_, prod_accum_61__52_, prod_accum_61__51_, prod_accum_61__50_, prod_accum_61__49_, prod_accum_61__48_, prod_accum_61__47_, prod_accum_61__46_, prod_accum_61__45_, prod_accum_61__44_, prod_accum_61__43_, prod_accum_61__42_, prod_accum_61__41_, prod_accum_61__40_, prod_accum_61__39_, prod_accum_61__38_, prod_accum_61__37_, prod_accum_61__36_, prod_accum_61__35_, prod_accum_61__34_, prod_accum_61__33_, prod_accum_61__32_, prod_accum_61__31_, prod_accum_61__30_, prod_accum_61__29_, prod_accum_61__28_, prod_accum_61__27_, prod_accum_61__26_, prod_accum_61__25_, prod_accum_61__24_, prod_accum_61__23_, prod_accum_61__22_, prod_accum_61__21_, prod_accum_61__20_, prod_accum_61__19_, prod_accum_61__18_, prod_accum_61__17_, prod_accum_61__16_, prod_accum_61__15_, prod_accum_61__14_, prod_accum_61__13_, prod_accum_61__12_, prod_accum_61__11_, prod_accum_61__10_, prod_accum_61__9_, prod_accum_61__8_, prod_accum_61__7_, prod_accum_61__6_, prod_accum_61__5_, prod_accum_61__4_, prod_accum_61__3_, prod_accum_61__2_, prod_accum_61__1_, prod_accum_61__0_ })
  );


  bsg_mul_array_row_128_62_x
  genblk1_62__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[7935:7808]),
    .b_i(b_r[7935:7808]),
    .s_i({ s_r_61__127_, s_r_61__126_, s_r_61__125_, s_r_61__124_, s_r_61__123_, s_r_61__122_, s_r_61__121_, s_r_61__120_, s_r_61__119_, s_r_61__118_, s_r_61__117_, s_r_61__116_, s_r_61__115_, s_r_61__114_, s_r_61__113_, s_r_61__112_, s_r_61__111_, s_r_61__110_, s_r_61__109_, s_r_61__108_, s_r_61__107_, s_r_61__106_, s_r_61__105_, s_r_61__104_, s_r_61__103_, s_r_61__102_, s_r_61__101_, s_r_61__100_, s_r_61__99_, s_r_61__98_, s_r_61__97_, s_r_61__96_, s_r_61__95_, s_r_61__94_, s_r_61__93_, s_r_61__92_, s_r_61__91_, s_r_61__90_, s_r_61__89_, s_r_61__88_, s_r_61__87_, s_r_61__86_, s_r_61__85_, s_r_61__84_, s_r_61__83_, s_r_61__82_, s_r_61__81_, s_r_61__80_, s_r_61__79_, s_r_61__78_, s_r_61__77_, s_r_61__76_, s_r_61__75_, s_r_61__74_, s_r_61__73_, s_r_61__72_, s_r_61__71_, s_r_61__70_, s_r_61__69_, s_r_61__68_, s_r_61__67_, s_r_61__66_, s_r_61__65_, s_r_61__64_, s_r_61__63_, s_r_61__62_, s_r_61__61_, s_r_61__60_, s_r_61__59_, s_r_61__58_, s_r_61__57_, s_r_61__56_, s_r_61__55_, s_r_61__54_, s_r_61__53_, s_r_61__52_, s_r_61__51_, s_r_61__50_, s_r_61__49_, s_r_61__48_, s_r_61__47_, s_r_61__46_, s_r_61__45_, s_r_61__44_, s_r_61__43_, s_r_61__42_, s_r_61__41_, s_r_61__40_, s_r_61__39_, s_r_61__38_, s_r_61__37_, s_r_61__36_, s_r_61__35_, s_r_61__34_, s_r_61__33_, s_r_61__32_, s_r_61__31_, s_r_61__30_, s_r_61__29_, s_r_61__28_, s_r_61__27_, s_r_61__26_, s_r_61__25_, s_r_61__24_, s_r_61__23_, s_r_61__22_, s_r_61__21_, s_r_61__20_, s_r_61__19_, s_r_61__18_, s_r_61__17_, s_r_61__16_, s_r_61__15_, s_r_61__14_, s_r_61__13_, s_r_61__12_, s_r_61__11_, s_r_61__10_, s_r_61__9_, s_r_61__8_, s_r_61__7_, s_r_61__6_, s_r_61__5_, s_r_61__4_, s_r_61__3_, s_r_61__2_, s_r_61__1_, s_r_61__0_ }),
    .c_i(c_r[61]),
    .prod_accum_i({ prod_accum_61__62_, prod_accum_61__61_, prod_accum_61__60_, prod_accum_61__59_, prod_accum_61__58_, prod_accum_61__57_, prod_accum_61__56_, prod_accum_61__55_, prod_accum_61__54_, prod_accum_61__53_, prod_accum_61__52_, prod_accum_61__51_, prod_accum_61__50_, prod_accum_61__49_, prod_accum_61__48_, prod_accum_61__47_, prod_accum_61__46_, prod_accum_61__45_, prod_accum_61__44_, prod_accum_61__43_, prod_accum_61__42_, prod_accum_61__41_, prod_accum_61__40_, prod_accum_61__39_, prod_accum_61__38_, prod_accum_61__37_, prod_accum_61__36_, prod_accum_61__35_, prod_accum_61__34_, prod_accum_61__33_, prod_accum_61__32_, prod_accum_61__31_, prod_accum_61__30_, prod_accum_61__29_, prod_accum_61__28_, prod_accum_61__27_, prod_accum_61__26_, prod_accum_61__25_, prod_accum_61__24_, prod_accum_61__23_, prod_accum_61__22_, prod_accum_61__21_, prod_accum_61__20_, prod_accum_61__19_, prod_accum_61__18_, prod_accum_61__17_, prod_accum_61__16_, prod_accum_61__15_, prod_accum_61__14_, prod_accum_61__13_, prod_accum_61__12_, prod_accum_61__11_, prod_accum_61__10_, prod_accum_61__9_, prod_accum_61__8_, prod_accum_61__7_, prod_accum_61__6_, prod_accum_61__5_, prod_accum_61__4_, prod_accum_61__3_, prod_accum_61__2_, prod_accum_61__1_, prod_accum_61__0_ }),
    .a_o(a_r[8063:7936]),
    .b_o(b_r[8063:7936]),
    .s_o({ s_r_62__127_, s_r_62__126_, s_r_62__125_, s_r_62__124_, s_r_62__123_, s_r_62__122_, s_r_62__121_, s_r_62__120_, s_r_62__119_, s_r_62__118_, s_r_62__117_, s_r_62__116_, s_r_62__115_, s_r_62__114_, s_r_62__113_, s_r_62__112_, s_r_62__111_, s_r_62__110_, s_r_62__109_, s_r_62__108_, s_r_62__107_, s_r_62__106_, s_r_62__105_, s_r_62__104_, s_r_62__103_, s_r_62__102_, s_r_62__101_, s_r_62__100_, s_r_62__99_, s_r_62__98_, s_r_62__97_, s_r_62__96_, s_r_62__95_, s_r_62__94_, s_r_62__93_, s_r_62__92_, s_r_62__91_, s_r_62__90_, s_r_62__89_, s_r_62__88_, s_r_62__87_, s_r_62__86_, s_r_62__85_, s_r_62__84_, s_r_62__83_, s_r_62__82_, s_r_62__81_, s_r_62__80_, s_r_62__79_, s_r_62__78_, s_r_62__77_, s_r_62__76_, s_r_62__75_, s_r_62__74_, s_r_62__73_, s_r_62__72_, s_r_62__71_, s_r_62__70_, s_r_62__69_, s_r_62__68_, s_r_62__67_, s_r_62__66_, s_r_62__65_, s_r_62__64_, s_r_62__63_, s_r_62__62_, s_r_62__61_, s_r_62__60_, s_r_62__59_, s_r_62__58_, s_r_62__57_, s_r_62__56_, s_r_62__55_, s_r_62__54_, s_r_62__53_, s_r_62__52_, s_r_62__51_, s_r_62__50_, s_r_62__49_, s_r_62__48_, s_r_62__47_, s_r_62__46_, s_r_62__45_, s_r_62__44_, s_r_62__43_, s_r_62__42_, s_r_62__41_, s_r_62__40_, s_r_62__39_, s_r_62__38_, s_r_62__37_, s_r_62__36_, s_r_62__35_, s_r_62__34_, s_r_62__33_, s_r_62__32_, s_r_62__31_, s_r_62__30_, s_r_62__29_, s_r_62__28_, s_r_62__27_, s_r_62__26_, s_r_62__25_, s_r_62__24_, s_r_62__23_, s_r_62__22_, s_r_62__21_, s_r_62__20_, s_r_62__19_, s_r_62__18_, s_r_62__17_, s_r_62__16_, s_r_62__15_, s_r_62__14_, s_r_62__13_, s_r_62__12_, s_r_62__11_, s_r_62__10_, s_r_62__9_, s_r_62__8_, s_r_62__7_, s_r_62__6_, s_r_62__5_, s_r_62__4_, s_r_62__3_, s_r_62__2_, s_r_62__1_, s_r_62__0_ }),
    .c_o(c_r[62]),
    .prod_accum_o({ prod_accum_62__63_, prod_accum_62__62_, prod_accum_62__61_, prod_accum_62__60_, prod_accum_62__59_, prod_accum_62__58_, prod_accum_62__57_, prod_accum_62__56_, prod_accum_62__55_, prod_accum_62__54_, prod_accum_62__53_, prod_accum_62__52_, prod_accum_62__51_, prod_accum_62__50_, prod_accum_62__49_, prod_accum_62__48_, prod_accum_62__47_, prod_accum_62__46_, prod_accum_62__45_, prod_accum_62__44_, prod_accum_62__43_, prod_accum_62__42_, prod_accum_62__41_, prod_accum_62__40_, prod_accum_62__39_, prod_accum_62__38_, prod_accum_62__37_, prod_accum_62__36_, prod_accum_62__35_, prod_accum_62__34_, prod_accum_62__33_, prod_accum_62__32_, prod_accum_62__31_, prod_accum_62__30_, prod_accum_62__29_, prod_accum_62__28_, prod_accum_62__27_, prod_accum_62__26_, prod_accum_62__25_, prod_accum_62__24_, prod_accum_62__23_, prod_accum_62__22_, prod_accum_62__21_, prod_accum_62__20_, prod_accum_62__19_, prod_accum_62__18_, prod_accum_62__17_, prod_accum_62__16_, prod_accum_62__15_, prod_accum_62__14_, prod_accum_62__13_, prod_accum_62__12_, prod_accum_62__11_, prod_accum_62__10_, prod_accum_62__9_, prod_accum_62__8_, prod_accum_62__7_, prod_accum_62__6_, prod_accum_62__5_, prod_accum_62__4_, prod_accum_62__3_, prod_accum_62__2_, prod_accum_62__1_, prod_accum_62__0_ })
  );


  bsg_mul_array_row_128_63_x
  genblk1_63__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[8063:7936]),
    .b_i(b_r[8063:7936]),
    .s_i({ s_r_62__127_, s_r_62__126_, s_r_62__125_, s_r_62__124_, s_r_62__123_, s_r_62__122_, s_r_62__121_, s_r_62__120_, s_r_62__119_, s_r_62__118_, s_r_62__117_, s_r_62__116_, s_r_62__115_, s_r_62__114_, s_r_62__113_, s_r_62__112_, s_r_62__111_, s_r_62__110_, s_r_62__109_, s_r_62__108_, s_r_62__107_, s_r_62__106_, s_r_62__105_, s_r_62__104_, s_r_62__103_, s_r_62__102_, s_r_62__101_, s_r_62__100_, s_r_62__99_, s_r_62__98_, s_r_62__97_, s_r_62__96_, s_r_62__95_, s_r_62__94_, s_r_62__93_, s_r_62__92_, s_r_62__91_, s_r_62__90_, s_r_62__89_, s_r_62__88_, s_r_62__87_, s_r_62__86_, s_r_62__85_, s_r_62__84_, s_r_62__83_, s_r_62__82_, s_r_62__81_, s_r_62__80_, s_r_62__79_, s_r_62__78_, s_r_62__77_, s_r_62__76_, s_r_62__75_, s_r_62__74_, s_r_62__73_, s_r_62__72_, s_r_62__71_, s_r_62__70_, s_r_62__69_, s_r_62__68_, s_r_62__67_, s_r_62__66_, s_r_62__65_, s_r_62__64_, s_r_62__63_, s_r_62__62_, s_r_62__61_, s_r_62__60_, s_r_62__59_, s_r_62__58_, s_r_62__57_, s_r_62__56_, s_r_62__55_, s_r_62__54_, s_r_62__53_, s_r_62__52_, s_r_62__51_, s_r_62__50_, s_r_62__49_, s_r_62__48_, s_r_62__47_, s_r_62__46_, s_r_62__45_, s_r_62__44_, s_r_62__43_, s_r_62__42_, s_r_62__41_, s_r_62__40_, s_r_62__39_, s_r_62__38_, s_r_62__37_, s_r_62__36_, s_r_62__35_, s_r_62__34_, s_r_62__33_, s_r_62__32_, s_r_62__31_, s_r_62__30_, s_r_62__29_, s_r_62__28_, s_r_62__27_, s_r_62__26_, s_r_62__25_, s_r_62__24_, s_r_62__23_, s_r_62__22_, s_r_62__21_, s_r_62__20_, s_r_62__19_, s_r_62__18_, s_r_62__17_, s_r_62__16_, s_r_62__15_, s_r_62__14_, s_r_62__13_, s_r_62__12_, s_r_62__11_, s_r_62__10_, s_r_62__9_, s_r_62__8_, s_r_62__7_, s_r_62__6_, s_r_62__5_, s_r_62__4_, s_r_62__3_, s_r_62__2_, s_r_62__1_, s_r_62__0_ }),
    .c_i(c_r[62]),
    .prod_accum_i({ prod_accum_62__63_, prod_accum_62__62_, prod_accum_62__61_, prod_accum_62__60_, prod_accum_62__59_, prod_accum_62__58_, prod_accum_62__57_, prod_accum_62__56_, prod_accum_62__55_, prod_accum_62__54_, prod_accum_62__53_, prod_accum_62__52_, prod_accum_62__51_, prod_accum_62__50_, prod_accum_62__49_, prod_accum_62__48_, prod_accum_62__47_, prod_accum_62__46_, prod_accum_62__45_, prod_accum_62__44_, prod_accum_62__43_, prod_accum_62__42_, prod_accum_62__41_, prod_accum_62__40_, prod_accum_62__39_, prod_accum_62__38_, prod_accum_62__37_, prod_accum_62__36_, prod_accum_62__35_, prod_accum_62__34_, prod_accum_62__33_, prod_accum_62__32_, prod_accum_62__31_, prod_accum_62__30_, prod_accum_62__29_, prod_accum_62__28_, prod_accum_62__27_, prod_accum_62__26_, prod_accum_62__25_, prod_accum_62__24_, prod_accum_62__23_, prod_accum_62__22_, prod_accum_62__21_, prod_accum_62__20_, prod_accum_62__19_, prod_accum_62__18_, prod_accum_62__17_, prod_accum_62__16_, prod_accum_62__15_, prod_accum_62__14_, prod_accum_62__13_, prod_accum_62__12_, prod_accum_62__11_, prod_accum_62__10_, prod_accum_62__9_, prod_accum_62__8_, prod_accum_62__7_, prod_accum_62__6_, prod_accum_62__5_, prod_accum_62__4_, prod_accum_62__3_, prod_accum_62__2_, prod_accum_62__1_, prod_accum_62__0_ }),
    .a_o(a_r[8191:8064]),
    .b_o(b_r[8191:8064]),
    .s_o({ s_r_63__127_, s_r_63__126_, s_r_63__125_, s_r_63__124_, s_r_63__123_, s_r_63__122_, s_r_63__121_, s_r_63__120_, s_r_63__119_, s_r_63__118_, s_r_63__117_, s_r_63__116_, s_r_63__115_, s_r_63__114_, s_r_63__113_, s_r_63__112_, s_r_63__111_, s_r_63__110_, s_r_63__109_, s_r_63__108_, s_r_63__107_, s_r_63__106_, s_r_63__105_, s_r_63__104_, s_r_63__103_, s_r_63__102_, s_r_63__101_, s_r_63__100_, s_r_63__99_, s_r_63__98_, s_r_63__97_, s_r_63__96_, s_r_63__95_, s_r_63__94_, s_r_63__93_, s_r_63__92_, s_r_63__91_, s_r_63__90_, s_r_63__89_, s_r_63__88_, s_r_63__87_, s_r_63__86_, s_r_63__85_, s_r_63__84_, s_r_63__83_, s_r_63__82_, s_r_63__81_, s_r_63__80_, s_r_63__79_, s_r_63__78_, s_r_63__77_, s_r_63__76_, s_r_63__75_, s_r_63__74_, s_r_63__73_, s_r_63__72_, s_r_63__71_, s_r_63__70_, s_r_63__69_, s_r_63__68_, s_r_63__67_, s_r_63__66_, s_r_63__65_, s_r_63__64_, s_r_63__63_, s_r_63__62_, s_r_63__61_, s_r_63__60_, s_r_63__59_, s_r_63__58_, s_r_63__57_, s_r_63__56_, s_r_63__55_, s_r_63__54_, s_r_63__53_, s_r_63__52_, s_r_63__51_, s_r_63__50_, s_r_63__49_, s_r_63__48_, s_r_63__47_, s_r_63__46_, s_r_63__45_, s_r_63__44_, s_r_63__43_, s_r_63__42_, s_r_63__41_, s_r_63__40_, s_r_63__39_, s_r_63__38_, s_r_63__37_, s_r_63__36_, s_r_63__35_, s_r_63__34_, s_r_63__33_, s_r_63__32_, s_r_63__31_, s_r_63__30_, s_r_63__29_, s_r_63__28_, s_r_63__27_, s_r_63__26_, s_r_63__25_, s_r_63__24_, s_r_63__23_, s_r_63__22_, s_r_63__21_, s_r_63__20_, s_r_63__19_, s_r_63__18_, s_r_63__17_, s_r_63__16_, s_r_63__15_, s_r_63__14_, s_r_63__13_, s_r_63__12_, s_r_63__11_, s_r_63__10_, s_r_63__9_, s_r_63__8_, s_r_63__7_, s_r_63__6_, s_r_63__5_, s_r_63__4_, s_r_63__3_, s_r_63__2_, s_r_63__1_, s_r_63__0_ }),
    .c_o(c_r[63]),
    .prod_accum_o({ prod_accum_63__64_, prod_accum_63__63_, prod_accum_63__62_, prod_accum_63__61_, prod_accum_63__60_, prod_accum_63__59_, prod_accum_63__58_, prod_accum_63__57_, prod_accum_63__56_, prod_accum_63__55_, prod_accum_63__54_, prod_accum_63__53_, prod_accum_63__52_, prod_accum_63__51_, prod_accum_63__50_, prod_accum_63__49_, prod_accum_63__48_, prod_accum_63__47_, prod_accum_63__46_, prod_accum_63__45_, prod_accum_63__44_, prod_accum_63__43_, prod_accum_63__42_, prod_accum_63__41_, prod_accum_63__40_, prod_accum_63__39_, prod_accum_63__38_, prod_accum_63__37_, prod_accum_63__36_, prod_accum_63__35_, prod_accum_63__34_, prod_accum_63__33_, prod_accum_63__32_, prod_accum_63__31_, prod_accum_63__30_, prod_accum_63__29_, prod_accum_63__28_, prod_accum_63__27_, prod_accum_63__26_, prod_accum_63__25_, prod_accum_63__24_, prod_accum_63__23_, prod_accum_63__22_, prod_accum_63__21_, prod_accum_63__20_, prod_accum_63__19_, prod_accum_63__18_, prod_accum_63__17_, prod_accum_63__16_, prod_accum_63__15_, prod_accum_63__14_, prod_accum_63__13_, prod_accum_63__12_, prod_accum_63__11_, prod_accum_63__10_, prod_accum_63__9_, prod_accum_63__8_, prod_accum_63__7_, prod_accum_63__6_, prod_accum_63__5_, prod_accum_63__4_, prod_accum_63__3_, prod_accum_63__2_, prod_accum_63__1_, prod_accum_63__0_ })
  );


  bsg_mul_array_row_128_64_x
  genblk1_64__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[8191:8064]),
    .b_i(b_r[8191:8064]),
    .s_i({ s_r_63__127_, s_r_63__126_, s_r_63__125_, s_r_63__124_, s_r_63__123_, s_r_63__122_, s_r_63__121_, s_r_63__120_, s_r_63__119_, s_r_63__118_, s_r_63__117_, s_r_63__116_, s_r_63__115_, s_r_63__114_, s_r_63__113_, s_r_63__112_, s_r_63__111_, s_r_63__110_, s_r_63__109_, s_r_63__108_, s_r_63__107_, s_r_63__106_, s_r_63__105_, s_r_63__104_, s_r_63__103_, s_r_63__102_, s_r_63__101_, s_r_63__100_, s_r_63__99_, s_r_63__98_, s_r_63__97_, s_r_63__96_, s_r_63__95_, s_r_63__94_, s_r_63__93_, s_r_63__92_, s_r_63__91_, s_r_63__90_, s_r_63__89_, s_r_63__88_, s_r_63__87_, s_r_63__86_, s_r_63__85_, s_r_63__84_, s_r_63__83_, s_r_63__82_, s_r_63__81_, s_r_63__80_, s_r_63__79_, s_r_63__78_, s_r_63__77_, s_r_63__76_, s_r_63__75_, s_r_63__74_, s_r_63__73_, s_r_63__72_, s_r_63__71_, s_r_63__70_, s_r_63__69_, s_r_63__68_, s_r_63__67_, s_r_63__66_, s_r_63__65_, s_r_63__64_, s_r_63__63_, s_r_63__62_, s_r_63__61_, s_r_63__60_, s_r_63__59_, s_r_63__58_, s_r_63__57_, s_r_63__56_, s_r_63__55_, s_r_63__54_, s_r_63__53_, s_r_63__52_, s_r_63__51_, s_r_63__50_, s_r_63__49_, s_r_63__48_, s_r_63__47_, s_r_63__46_, s_r_63__45_, s_r_63__44_, s_r_63__43_, s_r_63__42_, s_r_63__41_, s_r_63__40_, s_r_63__39_, s_r_63__38_, s_r_63__37_, s_r_63__36_, s_r_63__35_, s_r_63__34_, s_r_63__33_, s_r_63__32_, s_r_63__31_, s_r_63__30_, s_r_63__29_, s_r_63__28_, s_r_63__27_, s_r_63__26_, s_r_63__25_, s_r_63__24_, s_r_63__23_, s_r_63__22_, s_r_63__21_, s_r_63__20_, s_r_63__19_, s_r_63__18_, s_r_63__17_, s_r_63__16_, s_r_63__15_, s_r_63__14_, s_r_63__13_, s_r_63__12_, s_r_63__11_, s_r_63__10_, s_r_63__9_, s_r_63__8_, s_r_63__7_, s_r_63__6_, s_r_63__5_, s_r_63__4_, s_r_63__3_, s_r_63__2_, s_r_63__1_, s_r_63__0_ }),
    .c_i(c_r[63]),
    .prod_accum_i({ prod_accum_63__64_, prod_accum_63__63_, prod_accum_63__62_, prod_accum_63__61_, prod_accum_63__60_, prod_accum_63__59_, prod_accum_63__58_, prod_accum_63__57_, prod_accum_63__56_, prod_accum_63__55_, prod_accum_63__54_, prod_accum_63__53_, prod_accum_63__52_, prod_accum_63__51_, prod_accum_63__50_, prod_accum_63__49_, prod_accum_63__48_, prod_accum_63__47_, prod_accum_63__46_, prod_accum_63__45_, prod_accum_63__44_, prod_accum_63__43_, prod_accum_63__42_, prod_accum_63__41_, prod_accum_63__40_, prod_accum_63__39_, prod_accum_63__38_, prod_accum_63__37_, prod_accum_63__36_, prod_accum_63__35_, prod_accum_63__34_, prod_accum_63__33_, prod_accum_63__32_, prod_accum_63__31_, prod_accum_63__30_, prod_accum_63__29_, prod_accum_63__28_, prod_accum_63__27_, prod_accum_63__26_, prod_accum_63__25_, prod_accum_63__24_, prod_accum_63__23_, prod_accum_63__22_, prod_accum_63__21_, prod_accum_63__20_, prod_accum_63__19_, prod_accum_63__18_, prod_accum_63__17_, prod_accum_63__16_, prod_accum_63__15_, prod_accum_63__14_, prod_accum_63__13_, prod_accum_63__12_, prod_accum_63__11_, prod_accum_63__10_, prod_accum_63__9_, prod_accum_63__8_, prod_accum_63__7_, prod_accum_63__6_, prod_accum_63__5_, prod_accum_63__4_, prod_accum_63__3_, prod_accum_63__2_, prod_accum_63__1_, prod_accum_63__0_ }),
    .a_o(a_r[8319:8192]),
    .b_o(b_r[8319:8192]),
    .s_o({ s_r_64__127_, s_r_64__126_, s_r_64__125_, s_r_64__124_, s_r_64__123_, s_r_64__122_, s_r_64__121_, s_r_64__120_, s_r_64__119_, s_r_64__118_, s_r_64__117_, s_r_64__116_, s_r_64__115_, s_r_64__114_, s_r_64__113_, s_r_64__112_, s_r_64__111_, s_r_64__110_, s_r_64__109_, s_r_64__108_, s_r_64__107_, s_r_64__106_, s_r_64__105_, s_r_64__104_, s_r_64__103_, s_r_64__102_, s_r_64__101_, s_r_64__100_, s_r_64__99_, s_r_64__98_, s_r_64__97_, s_r_64__96_, s_r_64__95_, s_r_64__94_, s_r_64__93_, s_r_64__92_, s_r_64__91_, s_r_64__90_, s_r_64__89_, s_r_64__88_, s_r_64__87_, s_r_64__86_, s_r_64__85_, s_r_64__84_, s_r_64__83_, s_r_64__82_, s_r_64__81_, s_r_64__80_, s_r_64__79_, s_r_64__78_, s_r_64__77_, s_r_64__76_, s_r_64__75_, s_r_64__74_, s_r_64__73_, s_r_64__72_, s_r_64__71_, s_r_64__70_, s_r_64__69_, s_r_64__68_, s_r_64__67_, s_r_64__66_, s_r_64__65_, s_r_64__64_, s_r_64__63_, s_r_64__62_, s_r_64__61_, s_r_64__60_, s_r_64__59_, s_r_64__58_, s_r_64__57_, s_r_64__56_, s_r_64__55_, s_r_64__54_, s_r_64__53_, s_r_64__52_, s_r_64__51_, s_r_64__50_, s_r_64__49_, s_r_64__48_, s_r_64__47_, s_r_64__46_, s_r_64__45_, s_r_64__44_, s_r_64__43_, s_r_64__42_, s_r_64__41_, s_r_64__40_, s_r_64__39_, s_r_64__38_, s_r_64__37_, s_r_64__36_, s_r_64__35_, s_r_64__34_, s_r_64__33_, s_r_64__32_, s_r_64__31_, s_r_64__30_, s_r_64__29_, s_r_64__28_, s_r_64__27_, s_r_64__26_, s_r_64__25_, s_r_64__24_, s_r_64__23_, s_r_64__22_, s_r_64__21_, s_r_64__20_, s_r_64__19_, s_r_64__18_, s_r_64__17_, s_r_64__16_, s_r_64__15_, s_r_64__14_, s_r_64__13_, s_r_64__12_, s_r_64__11_, s_r_64__10_, s_r_64__9_, s_r_64__8_, s_r_64__7_, s_r_64__6_, s_r_64__5_, s_r_64__4_, s_r_64__3_, s_r_64__2_, s_r_64__1_, s_r_64__0_ }),
    .c_o(c_r[64]),
    .prod_accum_o({ prod_accum_64__65_, prod_accum_64__64_, prod_accum_64__63_, prod_accum_64__62_, prod_accum_64__61_, prod_accum_64__60_, prod_accum_64__59_, prod_accum_64__58_, prod_accum_64__57_, prod_accum_64__56_, prod_accum_64__55_, prod_accum_64__54_, prod_accum_64__53_, prod_accum_64__52_, prod_accum_64__51_, prod_accum_64__50_, prod_accum_64__49_, prod_accum_64__48_, prod_accum_64__47_, prod_accum_64__46_, prod_accum_64__45_, prod_accum_64__44_, prod_accum_64__43_, prod_accum_64__42_, prod_accum_64__41_, prod_accum_64__40_, prod_accum_64__39_, prod_accum_64__38_, prod_accum_64__37_, prod_accum_64__36_, prod_accum_64__35_, prod_accum_64__34_, prod_accum_64__33_, prod_accum_64__32_, prod_accum_64__31_, prod_accum_64__30_, prod_accum_64__29_, prod_accum_64__28_, prod_accum_64__27_, prod_accum_64__26_, prod_accum_64__25_, prod_accum_64__24_, prod_accum_64__23_, prod_accum_64__22_, prod_accum_64__21_, prod_accum_64__20_, prod_accum_64__19_, prod_accum_64__18_, prod_accum_64__17_, prod_accum_64__16_, prod_accum_64__15_, prod_accum_64__14_, prod_accum_64__13_, prod_accum_64__12_, prod_accum_64__11_, prod_accum_64__10_, prod_accum_64__9_, prod_accum_64__8_, prod_accum_64__7_, prod_accum_64__6_, prod_accum_64__5_, prod_accum_64__4_, prod_accum_64__3_, prod_accum_64__2_, prod_accum_64__1_, prod_accum_64__0_ })
  );


  bsg_mul_array_row_128_65_x
  genblk1_65__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[8319:8192]),
    .b_i(b_r[8319:8192]),
    .s_i({ s_r_64__127_, s_r_64__126_, s_r_64__125_, s_r_64__124_, s_r_64__123_, s_r_64__122_, s_r_64__121_, s_r_64__120_, s_r_64__119_, s_r_64__118_, s_r_64__117_, s_r_64__116_, s_r_64__115_, s_r_64__114_, s_r_64__113_, s_r_64__112_, s_r_64__111_, s_r_64__110_, s_r_64__109_, s_r_64__108_, s_r_64__107_, s_r_64__106_, s_r_64__105_, s_r_64__104_, s_r_64__103_, s_r_64__102_, s_r_64__101_, s_r_64__100_, s_r_64__99_, s_r_64__98_, s_r_64__97_, s_r_64__96_, s_r_64__95_, s_r_64__94_, s_r_64__93_, s_r_64__92_, s_r_64__91_, s_r_64__90_, s_r_64__89_, s_r_64__88_, s_r_64__87_, s_r_64__86_, s_r_64__85_, s_r_64__84_, s_r_64__83_, s_r_64__82_, s_r_64__81_, s_r_64__80_, s_r_64__79_, s_r_64__78_, s_r_64__77_, s_r_64__76_, s_r_64__75_, s_r_64__74_, s_r_64__73_, s_r_64__72_, s_r_64__71_, s_r_64__70_, s_r_64__69_, s_r_64__68_, s_r_64__67_, s_r_64__66_, s_r_64__65_, s_r_64__64_, s_r_64__63_, s_r_64__62_, s_r_64__61_, s_r_64__60_, s_r_64__59_, s_r_64__58_, s_r_64__57_, s_r_64__56_, s_r_64__55_, s_r_64__54_, s_r_64__53_, s_r_64__52_, s_r_64__51_, s_r_64__50_, s_r_64__49_, s_r_64__48_, s_r_64__47_, s_r_64__46_, s_r_64__45_, s_r_64__44_, s_r_64__43_, s_r_64__42_, s_r_64__41_, s_r_64__40_, s_r_64__39_, s_r_64__38_, s_r_64__37_, s_r_64__36_, s_r_64__35_, s_r_64__34_, s_r_64__33_, s_r_64__32_, s_r_64__31_, s_r_64__30_, s_r_64__29_, s_r_64__28_, s_r_64__27_, s_r_64__26_, s_r_64__25_, s_r_64__24_, s_r_64__23_, s_r_64__22_, s_r_64__21_, s_r_64__20_, s_r_64__19_, s_r_64__18_, s_r_64__17_, s_r_64__16_, s_r_64__15_, s_r_64__14_, s_r_64__13_, s_r_64__12_, s_r_64__11_, s_r_64__10_, s_r_64__9_, s_r_64__8_, s_r_64__7_, s_r_64__6_, s_r_64__5_, s_r_64__4_, s_r_64__3_, s_r_64__2_, s_r_64__1_, s_r_64__0_ }),
    .c_i(c_r[64]),
    .prod_accum_i({ prod_accum_64__65_, prod_accum_64__64_, prod_accum_64__63_, prod_accum_64__62_, prod_accum_64__61_, prod_accum_64__60_, prod_accum_64__59_, prod_accum_64__58_, prod_accum_64__57_, prod_accum_64__56_, prod_accum_64__55_, prod_accum_64__54_, prod_accum_64__53_, prod_accum_64__52_, prod_accum_64__51_, prod_accum_64__50_, prod_accum_64__49_, prod_accum_64__48_, prod_accum_64__47_, prod_accum_64__46_, prod_accum_64__45_, prod_accum_64__44_, prod_accum_64__43_, prod_accum_64__42_, prod_accum_64__41_, prod_accum_64__40_, prod_accum_64__39_, prod_accum_64__38_, prod_accum_64__37_, prod_accum_64__36_, prod_accum_64__35_, prod_accum_64__34_, prod_accum_64__33_, prod_accum_64__32_, prod_accum_64__31_, prod_accum_64__30_, prod_accum_64__29_, prod_accum_64__28_, prod_accum_64__27_, prod_accum_64__26_, prod_accum_64__25_, prod_accum_64__24_, prod_accum_64__23_, prod_accum_64__22_, prod_accum_64__21_, prod_accum_64__20_, prod_accum_64__19_, prod_accum_64__18_, prod_accum_64__17_, prod_accum_64__16_, prod_accum_64__15_, prod_accum_64__14_, prod_accum_64__13_, prod_accum_64__12_, prod_accum_64__11_, prod_accum_64__10_, prod_accum_64__9_, prod_accum_64__8_, prod_accum_64__7_, prod_accum_64__6_, prod_accum_64__5_, prod_accum_64__4_, prod_accum_64__3_, prod_accum_64__2_, prod_accum_64__1_, prod_accum_64__0_ }),
    .a_o(a_r[8447:8320]),
    .b_o(b_r[8447:8320]),
    .s_o({ s_r_65__127_, s_r_65__126_, s_r_65__125_, s_r_65__124_, s_r_65__123_, s_r_65__122_, s_r_65__121_, s_r_65__120_, s_r_65__119_, s_r_65__118_, s_r_65__117_, s_r_65__116_, s_r_65__115_, s_r_65__114_, s_r_65__113_, s_r_65__112_, s_r_65__111_, s_r_65__110_, s_r_65__109_, s_r_65__108_, s_r_65__107_, s_r_65__106_, s_r_65__105_, s_r_65__104_, s_r_65__103_, s_r_65__102_, s_r_65__101_, s_r_65__100_, s_r_65__99_, s_r_65__98_, s_r_65__97_, s_r_65__96_, s_r_65__95_, s_r_65__94_, s_r_65__93_, s_r_65__92_, s_r_65__91_, s_r_65__90_, s_r_65__89_, s_r_65__88_, s_r_65__87_, s_r_65__86_, s_r_65__85_, s_r_65__84_, s_r_65__83_, s_r_65__82_, s_r_65__81_, s_r_65__80_, s_r_65__79_, s_r_65__78_, s_r_65__77_, s_r_65__76_, s_r_65__75_, s_r_65__74_, s_r_65__73_, s_r_65__72_, s_r_65__71_, s_r_65__70_, s_r_65__69_, s_r_65__68_, s_r_65__67_, s_r_65__66_, s_r_65__65_, s_r_65__64_, s_r_65__63_, s_r_65__62_, s_r_65__61_, s_r_65__60_, s_r_65__59_, s_r_65__58_, s_r_65__57_, s_r_65__56_, s_r_65__55_, s_r_65__54_, s_r_65__53_, s_r_65__52_, s_r_65__51_, s_r_65__50_, s_r_65__49_, s_r_65__48_, s_r_65__47_, s_r_65__46_, s_r_65__45_, s_r_65__44_, s_r_65__43_, s_r_65__42_, s_r_65__41_, s_r_65__40_, s_r_65__39_, s_r_65__38_, s_r_65__37_, s_r_65__36_, s_r_65__35_, s_r_65__34_, s_r_65__33_, s_r_65__32_, s_r_65__31_, s_r_65__30_, s_r_65__29_, s_r_65__28_, s_r_65__27_, s_r_65__26_, s_r_65__25_, s_r_65__24_, s_r_65__23_, s_r_65__22_, s_r_65__21_, s_r_65__20_, s_r_65__19_, s_r_65__18_, s_r_65__17_, s_r_65__16_, s_r_65__15_, s_r_65__14_, s_r_65__13_, s_r_65__12_, s_r_65__11_, s_r_65__10_, s_r_65__9_, s_r_65__8_, s_r_65__7_, s_r_65__6_, s_r_65__5_, s_r_65__4_, s_r_65__3_, s_r_65__2_, s_r_65__1_, s_r_65__0_ }),
    .c_o(c_r[65]),
    .prod_accum_o({ prod_accum_65__66_, prod_accum_65__65_, prod_accum_65__64_, prod_accum_65__63_, prod_accum_65__62_, prod_accum_65__61_, prod_accum_65__60_, prod_accum_65__59_, prod_accum_65__58_, prod_accum_65__57_, prod_accum_65__56_, prod_accum_65__55_, prod_accum_65__54_, prod_accum_65__53_, prod_accum_65__52_, prod_accum_65__51_, prod_accum_65__50_, prod_accum_65__49_, prod_accum_65__48_, prod_accum_65__47_, prod_accum_65__46_, prod_accum_65__45_, prod_accum_65__44_, prod_accum_65__43_, prod_accum_65__42_, prod_accum_65__41_, prod_accum_65__40_, prod_accum_65__39_, prod_accum_65__38_, prod_accum_65__37_, prod_accum_65__36_, prod_accum_65__35_, prod_accum_65__34_, prod_accum_65__33_, prod_accum_65__32_, prod_accum_65__31_, prod_accum_65__30_, prod_accum_65__29_, prod_accum_65__28_, prod_accum_65__27_, prod_accum_65__26_, prod_accum_65__25_, prod_accum_65__24_, prod_accum_65__23_, prod_accum_65__22_, prod_accum_65__21_, prod_accum_65__20_, prod_accum_65__19_, prod_accum_65__18_, prod_accum_65__17_, prod_accum_65__16_, prod_accum_65__15_, prod_accum_65__14_, prod_accum_65__13_, prod_accum_65__12_, prod_accum_65__11_, prod_accum_65__10_, prod_accum_65__9_, prod_accum_65__8_, prod_accum_65__7_, prod_accum_65__6_, prod_accum_65__5_, prod_accum_65__4_, prod_accum_65__3_, prod_accum_65__2_, prod_accum_65__1_, prod_accum_65__0_ })
  );


  bsg_mul_array_row_128_66_x
  genblk1_66__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[8447:8320]),
    .b_i(b_r[8447:8320]),
    .s_i({ s_r_65__127_, s_r_65__126_, s_r_65__125_, s_r_65__124_, s_r_65__123_, s_r_65__122_, s_r_65__121_, s_r_65__120_, s_r_65__119_, s_r_65__118_, s_r_65__117_, s_r_65__116_, s_r_65__115_, s_r_65__114_, s_r_65__113_, s_r_65__112_, s_r_65__111_, s_r_65__110_, s_r_65__109_, s_r_65__108_, s_r_65__107_, s_r_65__106_, s_r_65__105_, s_r_65__104_, s_r_65__103_, s_r_65__102_, s_r_65__101_, s_r_65__100_, s_r_65__99_, s_r_65__98_, s_r_65__97_, s_r_65__96_, s_r_65__95_, s_r_65__94_, s_r_65__93_, s_r_65__92_, s_r_65__91_, s_r_65__90_, s_r_65__89_, s_r_65__88_, s_r_65__87_, s_r_65__86_, s_r_65__85_, s_r_65__84_, s_r_65__83_, s_r_65__82_, s_r_65__81_, s_r_65__80_, s_r_65__79_, s_r_65__78_, s_r_65__77_, s_r_65__76_, s_r_65__75_, s_r_65__74_, s_r_65__73_, s_r_65__72_, s_r_65__71_, s_r_65__70_, s_r_65__69_, s_r_65__68_, s_r_65__67_, s_r_65__66_, s_r_65__65_, s_r_65__64_, s_r_65__63_, s_r_65__62_, s_r_65__61_, s_r_65__60_, s_r_65__59_, s_r_65__58_, s_r_65__57_, s_r_65__56_, s_r_65__55_, s_r_65__54_, s_r_65__53_, s_r_65__52_, s_r_65__51_, s_r_65__50_, s_r_65__49_, s_r_65__48_, s_r_65__47_, s_r_65__46_, s_r_65__45_, s_r_65__44_, s_r_65__43_, s_r_65__42_, s_r_65__41_, s_r_65__40_, s_r_65__39_, s_r_65__38_, s_r_65__37_, s_r_65__36_, s_r_65__35_, s_r_65__34_, s_r_65__33_, s_r_65__32_, s_r_65__31_, s_r_65__30_, s_r_65__29_, s_r_65__28_, s_r_65__27_, s_r_65__26_, s_r_65__25_, s_r_65__24_, s_r_65__23_, s_r_65__22_, s_r_65__21_, s_r_65__20_, s_r_65__19_, s_r_65__18_, s_r_65__17_, s_r_65__16_, s_r_65__15_, s_r_65__14_, s_r_65__13_, s_r_65__12_, s_r_65__11_, s_r_65__10_, s_r_65__9_, s_r_65__8_, s_r_65__7_, s_r_65__6_, s_r_65__5_, s_r_65__4_, s_r_65__3_, s_r_65__2_, s_r_65__1_, s_r_65__0_ }),
    .c_i(c_r[65]),
    .prod_accum_i({ prod_accum_65__66_, prod_accum_65__65_, prod_accum_65__64_, prod_accum_65__63_, prod_accum_65__62_, prod_accum_65__61_, prod_accum_65__60_, prod_accum_65__59_, prod_accum_65__58_, prod_accum_65__57_, prod_accum_65__56_, prod_accum_65__55_, prod_accum_65__54_, prod_accum_65__53_, prod_accum_65__52_, prod_accum_65__51_, prod_accum_65__50_, prod_accum_65__49_, prod_accum_65__48_, prod_accum_65__47_, prod_accum_65__46_, prod_accum_65__45_, prod_accum_65__44_, prod_accum_65__43_, prod_accum_65__42_, prod_accum_65__41_, prod_accum_65__40_, prod_accum_65__39_, prod_accum_65__38_, prod_accum_65__37_, prod_accum_65__36_, prod_accum_65__35_, prod_accum_65__34_, prod_accum_65__33_, prod_accum_65__32_, prod_accum_65__31_, prod_accum_65__30_, prod_accum_65__29_, prod_accum_65__28_, prod_accum_65__27_, prod_accum_65__26_, prod_accum_65__25_, prod_accum_65__24_, prod_accum_65__23_, prod_accum_65__22_, prod_accum_65__21_, prod_accum_65__20_, prod_accum_65__19_, prod_accum_65__18_, prod_accum_65__17_, prod_accum_65__16_, prod_accum_65__15_, prod_accum_65__14_, prod_accum_65__13_, prod_accum_65__12_, prod_accum_65__11_, prod_accum_65__10_, prod_accum_65__9_, prod_accum_65__8_, prod_accum_65__7_, prod_accum_65__6_, prod_accum_65__5_, prod_accum_65__4_, prod_accum_65__3_, prod_accum_65__2_, prod_accum_65__1_, prod_accum_65__0_ }),
    .a_o(a_r[8575:8448]),
    .b_o(b_r[8575:8448]),
    .s_o({ s_r_66__127_, s_r_66__126_, s_r_66__125_, s_r_66__124_, s_r_66__123_, s_r_66__122_, s_r_66__121_, s_r_66__120_, s_r_66__119_, s_r_66__118_, s_r_66__117_, s_r_66__116_, s_r_66__115_, s_r_66__114_, s_r_66__113_, s_r_66__112_, s_r_66__111_, s_r_66__110_, s_r_66__109_, s_r_66__108_, s_r_66__107_, s_r_66__106_, s_r_66__105_, s_r_66__104_, s_r_66__103_, s_r_66__102_, s_r_66__101_, s_r_66__100_, s_r_66__99_, s_r_66__98_, s_r_66__97_, s_r_66__96_, s_r_66__95_, s_r_66__94_, s_r_66__93_, s_r_66__92_, s_r_66__91_, s_r_66__90_, s_r_66__89_, s_r_66__88_, s_r_66__87_, s_r_66__86_, s_r_66__85_, s_r_66__84_, s_r_66__83_, s_r_66__82_, s_r_66__81_, s_r_66__80_, s_r_66__79_, s_r_66__78_, s_r_66__77_, s_r_66__76_, s_r_66__75_, s_r_66__74_, s_r_66__73_, s_r_66__72_, s_r_66__71_, s_r_66__70_, s_r_66__69_, s_r_66__68_, s_r_66__67_, s_r_66__66_, s_r_66__65_, s_r_66__64_, s_r_66__63_, s_r_66__62_, s_r_66__61_, s_r_66__60_, s_r_66__59_, s_r_66__58_, s_r_66__57_, s_r_66__56_, s_r_66__55_, s_r_66__54_, s_r_66__53_, s_r_66__52_, s_r_66__51_, s_r_66__50_, s_r_66__49_, s_r_66__48_, s_r_66__47_, s_r_66__46_, s_r_66__45_, s_r_66__44_, s_r_66__43_, s_r_66__42_, s_r_66__41_, s_r_66__40_, s_r_66__39_, s_r_66__38_, s_r_66__37_, s_r_66__36_, s_r_66__35_, s_r_66__34_, s_r_66__33_, s_r_66__32_, s_r_66__31_, s_r_66__30_, s_r_66__29_, s_r_66__28_, s_r_66__27_, s_r_66__26_, s_r_66__25_, s_r_66__24_, s_r_66__23_, s_r_66__22_, s_r_66__21_, s_r_66__20_, s_r_66__19_, s_r_66__18_, s_r_66__17_, s_r_66__16_, s_r_66__15_, s_r_66__14_, s_r_66__13_, s_r_66__12_, s_r_66__11_, s_r_66__10_, s_r_66__9_, s_r_66__8_, s_r_66__7_, s_r_66__6_, s_r_66__5_, s_r_66__4_, s_r_66__3_, s_r_66__2_, s_r_66__1_, s_r_66__0_ }),
    .c_o(c_r[66]),
    .prod_accum_o({ prod_accum_66__67_, prod_accum_66__66_, prod_accum_66__65_, prod_accum_66__64_, prod_accum_66__63_, prod_accum_66__62_, prod_accum_66__61_, prod_accum_66__60_, prod_accum_66__59_, prod_accum_66__58_, prod_accum_66__57_, prod_accum_66__56_, prod_accum_66__55_, prod_accum_66__54_, prod_accum_66__53_, prod_accum_66__52_, prod_accum_66__51_, prod_accum_66__50_, prod_accum_66__49_, prod_accum_66__48_, prod_accum_66__47_, prod_accum_66__46_, prod_accum_66__45_, prod_accum_66__44_, prod_accum_66__43_, prod_accum_66__42_, prod_accum_66__41_, prod_accum_66__40_, prod_accum_66__39_, prod_accum_66__38_, prod_accum_66__37_, prod_accum_66__36_, prod_accum_66__35_, prod_accum_66__34_, prod_accum_66__33_, prod_accum_66__32_, prod_accum_66__31_, prod_accum_66__30_, prod_accum_66__29_, prod_accum_66__28_, prod_accum_66__27_, prod_accum_66__26_, prod_accum_66__25_, prod_accum_66__24_, prod_accum_66__23_, prod_accum_66__22_, prod_accum_66__21_, prod_accum_66__20_, prod_accum_66__19_, prod_accum_66__18_, prod_accum_66__17_, prod_accum_66__16_, prod_accum_66__15_, prod_accum_66__14_, prod_accum_66__13_, prod_accum_66__12_, prod_accum_66__11_, prod_accum_66__10_, prod_accum_66__9_, prod_accum_66__8_, prod_accum_66__7_, prod_accum_66__6_, prod_accum_66__5_, prod_accum_66__4_, prod_accum_66__3_, prod_accum_66__2_, prod_accum_66__1_, prod_accum_66__0_ })
  );


  bsg_mul_array_row_128_67_x
  genblk1_67__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[8575:8448]),
    .b_i(b_r[8575:8448]),
    .s_i({ s_r_66__127_, s_r_66__126_, s_r_66__125_, s_r_66__124_, s_r_66__123_, s_r_66__122_, s_r_66__121_, s_r_66__120_, s_r_66__119_, s_r_66__118_, s_r_66__117_, s_r_66__116_, s_r_66__115_, s_r_66__114_, s_r_66__113_, s_r_66__112_, s_r_66__111_, s_r_66__110_, s_r_66__109_, s_r_66__108_, s_r_66__107_, s_r_66__106_, s_r_66__105_, s_r_66__104_, s_r_66__103_, s_r_66__102_, s_r_66__101_, s_r_66__100_, s_r_66__99_, s_r_66__98_, s_r_66__97_, s_r_66__96_, s_r_66__95_, s_r_66__94_, s_r_66__93_, s_r_66__92_, s_r_66__91_, s_r_66__90_, s_r_66__89_, s_r_66__88_, s_r_66__87_, s_r_66__86_, s_r_66__85_, s_r_66__84_, s_r_66__83_, s_r_66__82_, s_r_66__81_, s_r_66__80_, s_r_66__79_, s_r_66__78_, s_r_66__77_, s_r_66__76_, s_r_66__75_, s_r_66__74_, s_r_66__73_, s_r_66__72_, s_r_66__71_, s_r_66__70_, s_r_66__69_, s_r_66__68_, s_r_66__67_, s_r_66__66_, s_r_66__65_, s_r_66__64_, s_r_66__63_, s_r_66__62_, s_r_66__61_, s_r_66__60_, s_r_66__59_, s_r_66__58_, s_r_66__57_, s_r_66__56_, s_r_66__55_, s_r_66__54_, s_r_66__53_, s_r_66__52_, s_r_66__51_, s_r_66__50_, s_r_66__49_, s_r_66__48_, s_r_66__47_, s_r_66__46_, s_r_66__45_, s_r_66__44_, s_r_66__43_, s_r_66__42_, s_r_66__41_, s_r_66__40_, s_r_66__39_, s_r_66__38_, s_r_66__37_, s_r_66__36_, s_r_66__35_, s_r_66__34_, s_r_66__33_, s_r_66__32_, s_r_66__31_, s_r_66__30_, s_r_66__29_, s_r_66__28_, s_r_66__27_, s_r_66__26_, s_r_66__25_, s_r_66__24_, s_r_66__23_, s_r_66__22_, s_r_66__21_, s_r_66__20_, s_r_66__19_, s_r_66__18_, s_r_66__17_, s_r_66__16_, s_r_66__15_, s_r_66__14_, s_r_66__13_, s_r_66__12_, s_r_66__11_, s_r_66__10_, s_r_66__9_, s_r_66__8_, s_r_66__7_, s_r_66__6_, s_r_66__5_, s_r_66__4_, s_r_66__3_, s_r_66__2_, s_r_66__1_, s_r_66__0_ }),
    .c_i(c_r[66]),
    .prod_accum_i({ prod_accum_66__67_, prod_accum_66__66_, prod_accum_66__65_, prod_accum_66__64_, prod_accum_66__63_, prod_accum_66__62_, prod_accum_66__61_, prod_accum_66__60_, prod_accum_66__59_, prod_accum_66__58_, prod_accum_66__57_, prod_accum_66__56_, prod_accum_66__55_, prod_accum_66__54_, prod_accum_66__53_, prod_accum_66__52_, prod_accum_66__51_, prod_accum_66__50_, prod_accum_66__49_, prod_accum_66__48_, prod_accum_66__47_, prod_accum_66__46_, prod_accum_66__45_, prod_accum_66__44_, prod_accum_66__43_, prod_accum_66__42_, prod_accum_66__41_, prod_accum_66__40_, prod_accum_66__39_, prod_accum_66__38_, prod_accum_66__37_, prod_accum_66__36_, prod_accum_66__35_, prod_accum_66__34_, prod_accum_66__33_, prod_accum_66__32_, prod_accum_66__31_, prod_accum_66__30_, prod_accum_66__29_, prod_accum_66__28_, prod_accum_66__27_, prod_accum_66__26_, prod_accum_66__25_, prod_accum_66__24_, prod_accum_66__23_, prod_accum_66__22_, prod_accum_66__21_, prod_accum_66__20_, prod_accum_66__19_, prod_accum_66__18_, prod_accum_66__17_, prod_accum_66__16_, prod_accum_66__15_, prod_accum_66__14_, prod_accum_66__13_, prod_accum_66__12_, prod_accum_66__11_, prod_accum_66__10_, prod_accum_66__9_, prod_accum_66__8_, prod_accum_66__7_, prod_accum_66__6_, prod_accum_66__5_, prod_accum_66__4_, prod_accum_66__3_, prod_accum_66__2_, prod_accum_66__1_, prod_accum_66__0_ }),
    .a_o(a_r[8703:8576]),
    .b_o(b_r[8703:8576]),
    .s_o({ s_r_67__127_, s_r_67__126_, s_r_67__125_, s_r_67__124_, s_r_67__123_, s_r_67__122_, s_r_67__121_, s_r_67__120_, s_r_67__119_, s_r_67__118_, s_r_67__117_, s_r_67__116_, s_r_67__115_, s_r_67__114_, s_r_67__113_, s_r_67__112_, s_r_67__111_, s_r_67__110_, s_r_67__109_, s_r_67__108_, s_r_67__107_, s_r_67__106_, s_r_67__105_, s_r_67__104_, s_r_67__103_, s_r_67__102_, s_r_67__101_, s_r_67__100_, s_r_67__99_, s_r_67__98_, s_r_67__97_, s_r_67__96_, s_r_67__95_, s_r_67__94_, s_r_67__93_, s_r_67__92_, s_r_67__91_, s_r_67__90_, s_r_67__89_, s_r_67__88_, s_r_67__87_, s_r_67__86_, s_r_67__85_, s_r_67__84_, s_r_67__83_, s_r_67__82_, s_r_67__81_, s_r_67__80_, s_r_67__79_, s_r_67__78_, s_r_67__77_, s_r_67__76_, s_r_67__75_, s_r_67__74_, s_r_67__73_, s_r_67__72_, s_r_67__71_, s_r_67__70_, s_r_67__69_, s_r_67__68_, s_r_67__67_, s_r_67__66_, s_r_67__65_, s_r_67__64_, s_r_67__63_, s_r_67__62_, s_r_67__61_, s_r_67__60_, s_r_67__59_, s_r_67__58_, s_r_67__57_, s_r_67__56_, s_r_67__55_, s_r_67__54_, s_r_67__53_, s_r_67__52_, s_r_67__51_, s_r_67__50_, s_r_67__49_, s_r_67__48_, s_r_67__47_, s_r_67__46_, s_r_67__45_, s_r_67__44_, s_r_67__43_, s_r_67__42_, s_r_67__41_, s_r_67__40_, s_r_67__39_, s_r_67__38_, s_r_67__37_, s_r_67__36_, s_r_67__35_, s_r_67__34_, s_r_67__33_, s_r_67__32_, s_r_67__31_, s_r_67__30_, s_r_67__29_, s_r_67__28_, s_r_67__27_, s_r_67__26_, s_r_67__25_, s_r_67__24_, s_r_67__23_, s_r_67__22_, s_r_67__21_, s_r_67__20_, s_r_67__19_, s_r_67__18_, s_r_67__17_, s_r_67__16_, s_r_67__15_, s_r_67__14_, s_r_67__13_, s_r_67__12_, s_r_67__11_, s_r_67__10_, s_r_67__9_, s_r_67__8_, s_r_67__7_, s_r_67__6_, s_r_67__5_, s_r_67__4_, s_r_67__3_, s_r_67__2_, s_r_67__1_, s_r_67__0_ }),
    .c_o(c_r[67]),
    .prod_accum_o({ prod_accum_67__68_, prod_accum_67__67_, prod_accum_67__66_, prod_accum_67__65_, prod_accum_67__64_, prod_accum_67__63_, prod_accum_67__62_, prod_accum_67__61_, prod_accum_67__60_, prod_accum_67__59_, prod_accum_67__58_, prod_accum_67__57_, prod_accum_67__56_, prod_accum_67__55_, prod_accum_67__54_, prod_accum_67__53_, prod_accum_67__52_, prod_accum_67__51_, prod_accum_67__50_, prod_accum_67__49_, prod_accum_67__48_, prod_accum_67__47_, prod_accum_67__46_, prod_accum_67__45_, prod_accum_67__44_, prod_accum_67__43_, prod_accum_67__42_, prod_accum_67__41_, prod_accum_67__40_, prod_accum_67__39_, prod_accum_67__38_, prod_accum_67__37_, prod_accum_67__36_, prod_accum_67__35_, prod_accum_67__34_, prod_accum_67__33_, prod_accum_67__32_, prod_accum_67__31_, prod_accum_67__30_, prod_accum_67__29_, prod_accum_67__28_, prod_accum_67__27_, prod_accum_67__26_, prod_accum_67__25_, prod_accum_67__24_, prod_accum_67__23_, prod_accum_67__22_, prod_accum_67__21_, prod_accum_67__20_, prod_accum_67__19_, prod_accum_67__18_, prod_accum_67__17_, prod_accum_67__16_, prod_accum_67__15_, prod_accum_67__14_, prod_accum_67__13_, prod_accum_67__12_, prod_accum_67__11_, prod_accum_67__10_, prod_accum_67__9_, prod_accum_67__8_, prod_accum_67__7_, prod_accum_67__6_, prod_accum_67__5_, prod_accum_67__4_, prod_accum_67__3_, prod_accum_67__2_, prod_accum_67__1_, prod_accum_67__0_ })
  );


  bsg_mul_array_row_128_68_x
  genblk1_68__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[8703:8576]),
    .b_i(b_r[8703:8576]),
    .s_i({ s_r_67__127_, s_r_67__126_, s_r_67__125_, s_r_67__124_, s_r_67__123_, s_r_67__122_, s_r_67__121_, s_r_67__120_, s_r_67__119_, s_r_67__118_, s_r_67__117_, s_r_67__116_, s_r_67__115_, s_r_67__114_, s_r_67__113_, s_r_67__112_, s_r_67__111_, s_r_67__110_, s_r_67__109_, s_r_67__108_, s_r_67__107_, s_r_67__106_, s_r_67__105_, s_r_67__104_, s_r_67__103_, s_r_67__102_, s_r_67__101_, s_r_67__100_, s_r_67__99_, s_r_67__98_, s_r_67__97_, s_r_67__96_, s_r_67__95_, s_r_67__94_, s_r_67__93_, s_r_67__92_, s_r_67__91_, s_r_67__90_, s_r_67__89_, s_r_67__88_, s_r_67__87_, s_r_67__86_, s_r_67__85_, s_r_67__84_, s_r_67__83_, s_r_67__82_, s_r_67__81_, s_r_67__80_, s_r_67__79_, s_r_67__78_, s_r_67__77_, s_r_67__76_, s_r_67__75_, s_r_67__74_, s_r_67__73_, s_r_67__72_, s_r_67__71_, s_r_67__70_, s_r_67__69_, s_r_67__68_, s_r_67__67_, s_r_67__66_, s_r_67__65_, s_r_67__64_, s_r_67__63_, s_r_67__62_, s_r_67__61_, s_r_67__60_, s_r_67__59_, s_r_67__58_, s_r_67__57_, s_r_67__56_, s_r_67__55_, s_r_67__54_, s_r_67__53_, s_r_67__52_, s_r_67__51_, s_r_67__50_, s_r_67__49_, s_r_67__48_, s_r_67__47_, s_r_67__46_, s_r_67__45_, s_r_67__44_, s_r_67__43_, s_r_67__42_, s_r_67__41_, s_r_67__40_, s_r_67__39_, s_r_67__38_, s_r_67__37_, s_r_67__36_, s_r_67__35_, s_r_67__34_, s_r_67__33_, s_r_67__32_, s_r_67__31_, s_r_67__30_, s_r_67__29_, s_r_67__28_, s_r_67__27_, s_r_67__26_, s_r_67__25_, s_r_67__24_, s_r_67__23_, s_r_67__22_, s_r_67__21_, s_r_67__20_, s_r_67__19_, s_r_67__18_, s_r_67__17_, s_r_67__16_, s_r_67__15_, s_r_67__14_, s_r_67__13_, s_r_67__12_, s_r_67__11_, s_r_67__10_, s_r_67__9_, s_r_67__8_, s_r_67__7_, s_r_67__6_, s_r_67__5_, s_r_67__4_, s_r_67__3_, s_r_67__2_, s_r_67__1_, s_r_67__0_ }),
    .c_i(c_r[67]),
    .prod_accum_i({ prod_accum_67__68_, prod_accum_67__67_, prod_accum_67__66_, prod_accum_67__65_, prod_accum_67__64_, prod_accum_67__63_, prod_accum_67__62_, prod_accum_67__61_, prod_accum_67__60_, prod_accum_67__59_, prod_accum_67__58_, prod_accum_67__57_, prod_accum_67__56_, prod_accum_67__55_, prod_accum_67__54_, prod_accum_67__53_, prod_accum_67__52_, prod_accum_67__51_, prod_accum_67__50_, prod_accum_67__49_, prod_accum_67__48_, prod_accum_67__47_, prod_accum_67__46_, prod_accum_67__45_, prod_accum_67__44_, prod_accum_67__43_, prod_accum_67__42_, prod_accum_67__41_, prod_accum_67__40_, prod_accum_67__39_, prod_accum_67__38_, prod_accum_67__37_, prod_accum_67__36_, prod_accum_67__35_, prod_accum_67__34_, prod_accum_67__33_, prod_accum_67__32_, prod_accum_67__31_, prod_accum_67__30_, prod_accum_67__29_, prod_accum_67__28_, prod_accum_67__27_, prod_accum_67__26_, prod_accum_67__25_, prod_accum_67__24_, prod_accum_67__23_, prod_accum_67__22_, prod_accum_67__21_, prod_accum_67__20_, prod_accum_67__19_, prod_accum_67__18_, prod_accum_67__17_, prod_accum_67__16_, prod_accum_67__15_, prod_accum_67__14_, prod_accum_67__13_, prod_accum_67__12_, prod_accum_67__11_, prod_accum_67__10_, prod_accum_67__9_, prod_accum_67__8_, prod_accum_67__7_, prod_accum_67__6_, prod_accum_67__5_, prod_accum_67__4_, prod_accum_67__3_, prod_accum_67__2_, prod_accum_67__1_, prod_accum_67__0_ }),
    .a_o(a_r[8831:8704]),
    .b_o(b_r[8831:8704]),
    .s_o({ s_r_68__127_, s_r_68__126_, s_r_68__125_, s_r_68__124_, s_r_68__123_, s_r_68__122_, s_r_68__121_, s_r_68__120_, s_r_68__119_, s_r_68__118_, s_r_68__117_, s_r_68__116_, s_r_68__115_, s_r_68__114_, s_r_68__113_, s_r_68__112_, s_r_68__111_, s_r_68__110_, s_r_68__109_, s_r_68__108_, s_r_68__107_, s_r_68__106_, s_r_68__105_, s_r_68__104_, s_r_68__103_, s_r_68__102_, s_r_68__101_, s_r_68__100_, s_r_68__99_, s_r_68__98_, s_r_68__97_, s_r_68__96_, s_r_68__95_, s_r_68__94_, s_r_68__93_, s_r_68__92_, s_r_68__91_, s_r_68__90_, s_r_68__89_, s_r_68__88_, s_r_68__87_, s_r_68__86_, s_r_68__85_, s_r_68__84_, s_r_68__83_, s_r_68__82_, s_r_68__81_, s_r_68__80_, s_r_68__79_, s_r_68__78_, s_r_68__77_, s_r_68__76_, s_r_68__75_, s_r_68__74_, s_r_68__73_, s_r_68__72_, s_r_68__71_, s_r_68__70_, s_r_68__69_, s_r_68__68_, s_r_68__67_, s_r_68__66_, s_r_68__65_, s_r_68__64_, s_r_68__63_, s_r_68__62_, s_r_68__61_, s_r_68__60_, s_r_68__59_, s_r_68__58_, s_r_68__57_, s_r_68__56_, s_r_68__55_, s_r_68__54_, s_r_68__53_, s_r_68__52_, s_r_68__51_, s_r_68__50_, s_r_68__49_, s_r_68__48_, s_r_68__47_, s_r_68__46_, s_r_68__45_, s_r_68__44_, s_r_68__43_, s_r_68__42_, s_r_68__41_, s_r_68__40_, s_r_68__39_, s_r_68__38_, s_r_68__37_, s_r_68__36_, s_r_68__35_, s_r_68__34_, s_r_68__33_, s_r_68__32_, s_r_68__31_, s_r_68__30_, s_r_68__29_, s_r_68__28_, s_r_68__27_, s_r_68__26_, s_r_68__25_, s_r_68__24_, s_r_68__23_, s_r_68__22_, s_r_68__21_, s_r_68__20_, s_r_68__19_, s_r_68__18_, s_r_68__17_, s_r_68__16_, s_r_68__15_, s_r_68__14_, s_r_68__13_, s_r_68__12_, s_r_68__11_, s_r_68__10_, s_r_68__9_, s_r_68__8_, s_r_68__7_, s_r_68__6_, s_r_68__5_, s_r_68__4_, s_r_68__3_, s_r_68__2_, s_r_68__1_, s_r_68__0_ }),
    .c_o(c_r[68]),
    .prod_accum_o({ prod_accum_68__69_, prod_accum_68__68_, prod_accum_68__67_, prod_accum_68__66_, prod_accum_68__65_, prod_accum_68__64_, prod_accum_68__63_, prod_accum_68__62_, prod_accum_68__61_, prod_accum_68__60_, prod_accum_68__59_, prod_accum_68__58_, prod_accum_68__57_, prod_accum_68__56_, prod_accum_68__55_, prod_accum_68__54_, prod_accum_68__53_, prod_accum_68__52_, prod_accum_68__51_, prod_accum_68__50_, prod_accum_68__49_, prod_accum_68__48_, prod_accum_68__47_, prod_accum_68__46_, prod_accum_68__45_, prod_accum_68__44_, prod_accum_68__43_, prod_accum_68__42_, prod_accum_68__41_, prod_accum_68__40_, prod_accum_68__39_, prod_accum_68__38_, prod_accum_68__37_, prod_accum_68__36_, prod_accum_68__35_, prod_accum_68__34_, prod_accum_68__33_, prod_accum_68__32_, prod_accum_68__31_, prod_accum_68__30_, prod_accum_68__29_, prod_accum_68__28_, prod_accum_68__27_, prod_accum_68__26_, prod_accum_68__25_, prod_accum_68__24_, prod_accum_68__23_, prod_accum_68__22_, prod_accum_68__21_, prod_accum_68__20_, prod_accum_68__19_, prod_accum_68__18_, prod_accum_68__17_, prod_accum_68__16_, prod_accum_68__15_, prod_accum_68__14_, prod_accum_68__13_, prod_accum_68__12_, prod_accum_68__11_, prod_accum_68__10_, prod_accum_68__9_, prod_accum_68__8_, prod_accum_68__7_, prod_accum_68__6_, prod_accum_68__5_, prod_accum_68__4_, prod_accum_68__3_, prod_accum_68__2_, prod_accum_68__1_, prod_accum_68__0_ })
  );


  bsg_mul_array_row_128_69_x
  genblk1_69__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[8831:8704]),
    .b_i(b_r[8831:8704]),
    .s_i({ s_r_68__127_, s_r_68__126_, s_r_68__125_, s_r_68__124_, s_r_68__123_, s_r_68__122_, s_r_68__121_, s_r_68__120_, s_r_68__119_, s_r_68__118_, s_r_68__117_, s_r_68__116_, s_r_68__115_, s_r_68__114_, s_r_68__113_, s_r_68__112_, s_r_68__111_, s_r_68__110_, s_r_68__109_, s_r_68__108_, s_r_68__107_, s_r_68__106_, s_r_68__105_, s_r_68__104_, s_r_68__103_, s_r_68__102_, s_r_68__101_, s_r_68__100_, s_r_68__99_, s_r_68__98_, s_r_68__97_, s_r_68__96_, s_r_68__95_, s_r_68__94_, s_r_68__93_, s_r_68__92_, s_r_68__91_, s_r_68__90_, s_r_68__89_, s_r_68__88_, s_r_68__87_, s_r_68__86_, s_r_68__85_, s_r_68__84_, s_r_68__83_, s_r_68__82_, s_r_68__81_, s_r_68__80_, s_r_68__79_, s_r_68__78_, s_r_68__77_, s_r_68__76_, s_r_68__75_, s_r_68__74_, s_r_68__73_, s_r_68__72_, s_r_68__71_, s_r_68__70_, s_r_68__69_, s_r_68__68_, s_r_68__67_, s_r_68__66_, s_r_68__65_, s_r_68__64_, s_r_68__63_, s_r_68__62_, s_r_68__61_, s_r_68__60_, s_r_68__59_, s_r_68__58_, s_r_68__57_, s_r_68__56_, s_r_68__55_, s_r_68__54_, s_r_68__53_, s_r_68__52_, s_r_68__51_, s_r_68__50_, s_r_68__49_, s_r_68__48_, s_r_68__47_, s_r_68__46_, s_r_68__45_, s_r_68__44_, s_r_68__43_, s_r_68__42_, s_r_68__41_, s_r_68__40_, s_r_68__39_, s_r_68__38_, s_r_68__37_, s_r_68__36_, s_r_68__35_, s_r_68__34_, s_r_68__33_, s_r_68__32_, s_r_68__31_, s_r_68__30_, s_r_68__29_, s_r_68__28_, s_r_68__27_, s_r_68__26_, s_r_68__25_, s_r_68__24_, s_r_68__23_, s_r_68__22_, s_r_68__21_, s_r_68__20_, s_r_68__19_, s_r_68__18_, s_r_68__17_, s_r_68__16_, s_r_68__15_, s_r_68__14_, s_r_68__13_, s_r_68__12_, s_r_68__11_, s_r_68__10_, s_r_68__9_, s_r_68__8_, s_r_68__7_, s_r_68__6_, s_r_68__5_, s_r_68__4_, s_r_68__3_, s_r_68__2_, s_r_68__1_, s_r_68__0_ }),
    .c_i(c_r[68]),
    .prod_accum_i({ prod_accum_68__69_, prod_accum_68__68_, prod_accum_68__67_, prod_accum_68__66_, prod_accum_68__65_, prod_accum_68__64_, prod_accum_68__63_, prod_accum_68__62_, prod_accum_68__61_, prod_accum_68__60_, prod_accum_68__59_, prod_accum_68__58_, prod_accum_68__57_, prod_accum_68__56_, prod_accum_68__55_, prod_accum_68__54_, prod_accum_68__53_, prod_accum_68__52_, prod_accum_68__51_, prod_accum_68__50_, prod_accum_68__49_, prod_accum_68__48_, prod_accum_68__47_, prod_accum_68__46_, prod_accum_68__45_, prod_accum_68__44_, prod_accum_68__43_, prod_accum_68__42_, prod_accum_68__41_, prod_accum_68__40_, prod_accum_68__39_, prod_accum_68__38_, prod_accum_68__37_, prod_accum_68__36_, prod_accum_68__35_, prod_accum_68__34_, prod_accum_68__33_, prod_accum_68__32_, prod_accum_68__31_, prod_accum_68__30_, prod_accum_68__29_, prod_accum_68__28_, prod_accum_68__27_, prod_accum_68__26_, prod_accum_68__25_, prod_accum_68__24_, prod_accum_68__23_, prod_accum_68__22_, prod_accum_68__21_, prod_accum_68__20_, prod_accum_68__19_, prod_accum_68__18_, prod_accum_68__17_, prod_accum_68__16_, prod_accum_68__15_, prod_accum_68__14_, prod_accum_68__13_, prod_accum_68__12_, prod_accum_68__11_, prod_accum_68__10_, prod_accum_68__9_, prod_accum_68__8_, prod_accum_68__7_, prod_accum_68__6_, prod_accum_68__5_, prod_accum_68__4_, prod_accum_68__3_, prod_accum_68__2_, prod_accum_68__1_, prod_accum_68__0_ }),
    .a_o(a_r[8959:8832]),
    .b_o(b_r[8959:8832]),
    .s_o({ s_r_69__127_, s_r_69__126_, s_r_69__125_, s_r_69__124_, s_r_69__123_, s_r_69__122_, s_r_69__121_, s_r_69__120_, s_r_69__119_, s_r_69__118_, s_r_69__117_, s_r_69__116_, s_r_69__115_, s_r_69__114_, s_r_69__113_, s_r_69__112_, s_r_69__111_, s_r_69__110_, s_r_69__109_, s_r_69__108_, s_r_69__107_, s_r_69__106_, s_r_69__105_, s_r_69__104_, s_r_69__103_, s_r_69__102_, s_r_69__101_, s_r_69__100_, s_r_69__99_, s_r_69__98_, s_r_69__97_, s_r_69__96_, s_r_69__95_, s_r_69__94_, s_r_69__93_, s_r_69__92_, s_r_69__91_, s_r_69__90_, s_r_69__89_, s_r_69__88_, s_r_69__87_, s_r_69__86_, s_r_69__85_, s_r_69__84_, s_r_69__83_, s_r_69__82_, s_r_69__81_, s_r_69__80_, s_r_69__79_, s_r_69__78_, s_r_69__77_, s_r_69__76_, s_r_69__75_, s_r_69__74_, s_r_69__73_, s_r_69__72_, s_r_69__71_, s_r_69__70_, s_r_69__69_, s_r_69__68_, s_r_69__67_, s_r_69__66_, s_r_69__65_, s_r_69__64_, s_r_69__63_, s_r_69__62_, s_r_69__61_, s_r_69__60_, s_r_69__59_, s_r_69__58_, s_r_69__57_, s_r_69__56_, s_r_69__55_, s_r_69__54_, s_r_69__53_, s_r_69__52_, s_r_69__51_, s_r_69__50_, s_r_69__49_, s_r_69__48_, s_r_69__47_, s_r_69__46_, s_r_69__45_, s_r_69__44_, s_r_69__43_, s_r_69__42_, s_r_69__41_, s_r_69__40_, s_r_69__39_, s_r_69__38_, s_r_69__37_, s_r_69__36_, s_r_69__35_, s_r_69__34_, s_r_69__33_, s_r_69__32_, s_r_69__31_, s_r_69__30_, s_r_69__29_, s_r_69__28_, s_r_69__27_, s_r_69__26_, s_r_69__25_, s_r_69__24_, s_r_69__23_, s_r_69__22_, s_r_69__21_, s_r_69__20_, s_r_69__19_, s_r_69__18_, s_r_69__17_, s_r_69__16_, s_r_69__15_, s_r_69__14_, s_r_69__13_, s_r_69__12_, s_r_69__11_, s_r_69__10_, s_r_69__9_, s_r_69__8_, s_r_69__7_, s_r_69__6_, s_r_69__5_, s_r_69__4_, s_r_69__3_, s_r_69__2_, s_r_69__1_, s_r_69__0_ }),
    .c_o(c_r[69]),
    .prod_accum_o({ prod_accum_69__70_, prod_accum_69__69_, prod_accum_69__68_, prod_accum_69__67_, prod_accum_69__66_, prod_accum_69__65_, prod_accum_69__64_, prod_accum_69__63_, prod_accum_69__62_, prod_accum_69__61_, prod_accum_69__60_, prod_accum_69__59_, prod_accum_69__58_, prod_accum_69__57_, prod_accum_69__56_, prod_accum_69__55_, prod_accum_69__54_, prod_accum_69__53_, prod_accum_69__52_, prod_accum_69__51_, prod_accum_69__50_, prod_accum_69__49_, prod_accum_69__48_, prod_accum_69__47_, prod_accum_69__46_, prod_accum_69__45_, prod_accum_69__44_, prod_accum_69__43_, prod_accum_69__42_, prod_accum_69__41_, prod_accum_69__40_, prod_accum_69__39_, prod_accum_69__38_, prod_accum_69__37_, prod_accum_69__36_, prod_accum_69__35_, prod_accum_69__34_, prod_accum_69__33_, prod_accum_69__32_, prod_accum_69__31_, prod_accum_69__30_, prod_accum_69__29_, prod_accum_69__28_, prod_accum_69__27_, prod_accum_69__26_, prod_accum_69__25_, prod_accum_69__24_, prod_accum_69__23_, prod_accum_69__22_, prod_accum_69__21_, prod_accum_69__20_, prod_accum_69__19_, prod_accum_69__18_, prod_accum_69__17_, prod_accum_69__16_, prod_accum_69__15_, prod_accum_69__14_, prod_accum_69__13_, prod_accum_69__12_, prod_accum_69__11_, prod_accum_69__10_, prod_accum_69__9_, prod_accum_69__8_, prod_accum_69__7_, prod_accum_69__6_, prod_accum_69__5_, prod_accum_69__4_, prod_accum_69__3_, prod_accum_69__2_, prod_accum_69__1_, prod_accum_69__0_ })
  );


  bsg_mul_array_row_128_70_x
  genblk1_70__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[8959:8832]),
    .b_i(b_r[8959:8832]),
    .s_i({ s_r_69__127_, s_r_69__126_, s_r_69__125_, s_r_69__124_, s_r_69__123_, s_r_69__122_, s_r_69__121_, s_r_69__120_, s_r_69__119_, s_r_69__118_, s_r_69__117_, s_r_69__116_, s_r_69__115_, s_r_69__114_, s_r_69__113_, s_r_69__112_, s_r_69__111_, s_r_69__110_, s_r_69__109_, s_r_69__108_, s_r_69__107_, s_r_69__106_, s_r_69__105_, s_r_69__104_, s_r_69__103_, s_r_69__102_, s_r_69__101_, s_r_69__100_, s_r_69__99_, s_r_69__98_, s_r_69__97_, s_r_69__96_, s_r_69__95_, s_r_69__94_, s_r_69__93_, s_r_69__92_, s_r_69__91_, s_r_69__90_, s_r_69__89_, s_r_69__88_, s_r_69__87_, s_r_69__86_, s_r_69__85_, s_r_69__84_, s_r_69__83_, s_r_69__82_, s_r_69__81_, s_r_69__80_, s_r_69__79_, s_r_69__78_, s_r_69__77_, s_r_69__76_, s_r_69__75_, s_r_69__74_, s_r_69__73_, s_r_69__72_, s_r_69__71_, s_r_69__70_, s_r_69__69_, s_r_69__68_, s_r_69__67_, s_r_69__66_, s_r_69__65_, s_r_69__64_, s_r_69__63_, s_r_69__62_, s_r_69__61_, s_r_69__60_, s_r_69__59_, s_r_69__58_, s_r_69__57_, s_r_69__56_, s_r_69__55_, s_r_69__54_, s_r_69__53_, s_r_69__52_, s_r_69__51_, s_r_69__50_, s_r_69__49_, s_r_69__48_, s_r_69__47_, s_r_69__46_, s_r_69__45_, s_r_69__44_, s_r_69__43_, s_r_69__42_, s_r_69__41_, s_r_69__40_, s_r_69__39_, s_r_69__38_, s_r_69__37_, s_r_69__36_, s_r_69__35_, s_r_69__34_, s_r_69__33_, s_r_69__32_, s_r_69__31_, s_r_69__30_, s_r_69__29_, s_r_69__28_, s_r_69__27_, s_r_69__26_, s_r_69__25_, s_r_69__24_, s_r_69__23_, s_r_69__22_, s_r_69__21_, s_r_69__20_, s_r_69__19_, s_r_69__18_, s_r_69__17_, s_r_69__16_, s_r_69__15_, s_r_69__14_, s_r_69__13_, s_r_69__12_, s_r_69__11_, s_r_69__10_, s_r_69__9_, s_r_69__8_, s_r_69__7_, s_r_69__6_, s_r_69__5_, s_r_69__4_, s_r_69__3_, s_r_69__2_, s_r_69__1_, s_r_69__0_ }),
    .c_i(c_r[69]),
    .prod_accum_i({ prod_accum_69__70_, prod_accum_69__69_, prod_accum_69__68_, prod_accum_69__67_, prod_accum_69__66_, prod_accum_69__65_, prod_accum_69__64_, prod_accum_69__63_, prod_accum_69__62_, prod_accum_69__61_, prod_accum_69__60_, prod_accum_69__59_, prod_accum_69__58_, prod_accum_69__57_, prod_accum_69__56_, prod_accum_69__55_, prod_accum_69__54_, prod_accum_69__53_, prod_accum_69__52_, prod_accum_69__51_, prod_accum_69__50_, prod_accum_69__49_, prod_accum_69__48_, prod_accum_69__47_, prod_accum_69__46_, prod_accum_69__45_, prod_accum_69__44_, prod_accum_69__43_, prod_accum_69__42_, prod_accum_69__41_, prod_accum_69__40_, prod_accum_69__39_, prod_accum_69__38_, prod_accum_69__37_, prod_accum_69__36_, prod_accum_69__35_, prod_accum_69__34_, prod_accum_69__33_, prod_accum_69__32_, prod_accum_69__31_, prod_accum_69__30_, prod_accum_69__29_, prod_accum_69__28_, prod_accum_69__27_, prod_accum_69__26_, prod_accum_69__25_, prod_accum_69__24_, prod_accum_69__23_, prod_accum_69__22_, prod_accum_69__21_, prod_accum_69__20_, prod_accum_69__19_, prod_accum_69__18_, prod_accum_69__17_, prod_accum_69__16_, prod_accum_69__15_, prod_accum_69__14_, prod_accum_69__13_, prod_accum_69__12_, prod_accum_69__11_, prod_accum_69__10_, prod_accum_69__9_, prod_accum_69__8_, prod_accum_69__7_, prod_accum_69__6_, prod_accum_69__5_, prod_accum_69__4_, prod_accum_69__3_, prod_accum_69__2_, prod_accum_69__1_, prod_accum_69__0_ }),
    .a_o(a_r[9087:8960]),
    .b_o(b_r[9087:8960]),
    .s_o({ s_r_70__127_, s_r_70__126_, s_r_70__125_, s_r_70__124_, s_r_70__123_, s_r_70__122_, s_r_70__121_, s_r_70__120_, s_r_70__119_, s_r_70__118_, s_r_70__117_, s_r_70__116_, s_r_70__115_, s_r_70__114_, s_r_70__113_, s_r_70__112_, s_r_70__111_, s_r_70__110_, s_r_70__109_, s_r_70__108_, s_r_70__107_, s_r_70__106_, s_r_70__105_, s_r_70__104_, s_r_70__103_, s_r_70__102_, s_r_70__101_, s_r_70__100_, s_r_70__99_, s_r_70__98_, s_r_70__97_, s_r_70__96_, s_r_70__95_, s_r_70__94_, s_r_70__93_, s_r_70__92_, s_r_70__91_, s_r_70__90_, s_r_70__89_, s_r_70__88_, s_r_70__87_, s_r_70__86_, s_r_70__85_, s_r_70__84_, s_r_70__83_, s_r_70__82_, s_r_70__81_, s_r_70__80_, s_r_70__79_, s_r_70__78_, s_r_70__77_, s_r_70__76_, s_r_70__75_, s_r_70__74_, s_r_70__73_, s_r_70__72_, s_r_70__71_, s_r_70__70_, s_r_70__69_, s_r_70__68_, s_r_70__67_, s_r_70__66_, s_r_70__65_, s_r_70__64_, s_r_70__63_, s_r_70__62_, s_r_70__61_, s_r_70__60_, s_r_70__59_, s_r_70__58_, s_r_70__57_, s_r_70__56_, s_r_70__55_, s_r_70__54_, s_r_70__53_, s_r_70__52_, s_r_70__51_, s_r_70__50_, s_r_70__49_, s_r_70__48_, s_r_70__47_, s_r_70__46_, s_r_70__45_, s_r_70__44_, s_r_70__43_, s_r_70__42_, s_r_70__41_, s_r_70__40_, s_r_70__39_, s_r_70__38_, s_r_70__37_, s_r_70__36_, s_r_70__35_, s_r_70__34_, s_r_70__33_, s_r_70__32_, s_r_70__31_, s_r_70__30_, s_r_70__29_, s_r_70__28_, s_r_70__27_, s_r_70__26_, s_r_70__25_, s_r_70__24_, s_r_70__23_, s_r_70__22_, s_r_70__21_, s_r_70__20_, s_r_70__19_, s_r_70__18_, s_r_70__17_, s_r_70__16_, s_r_70__15_, s_r_70__14_, s_r_70__13_, s_r_70__12_, s_r_70__11_, s_r_70__10_, s_r_70__9_, s_r_70__8_, s_r_70__7_, s_r_70__6_, s_r_70__5_, s_r_70__4_, s_r_70__3_, s_r_70__2_, s_r_70__1_, s_r_70__0_ }),
    .c_o(c_r[70]),
    .prod_accum_o({ prod_accum_70__71_, prod_accum_70__70_, prod_accum_70__69_, prod_accum_70__68_, prod_accum_70__67_, prod_accum_70__66_, prod_accum_70__65_, prod_accum_70__64_, prod_accum_70__63_, prod_accum_70__62_, prod_accum_70__61_, prod_accum_70__60_, prod_accum_70__59_, prod_accum_70__58_, prod_accum_70__57_, prod_accum_70__56_, prod_accum_70__55_, prod_accum_70__54_, prod_accum_70__53_, prod_accum_70__52_, prod_accum_70__51_, prod_accum_70__50_, prod_accum_70__49_, prod_accum_70__48_, prod_accum_70__47_, prod_accum_70__46_, prod_accum_70__45_, prod_accum_70__44_, prod_accum_70__43_, prod_accum_70__42_, prod_accum_70__41_, prod_accum_70__40_, prod_accum_70__39_, prod_accum_70__38_, prod_accum_70__37_, prod_accum_70__36_, prod_accum_70__35_, prod_accum_70__34_, prod_accum_70__33_, prod_accum_70__32_, prod_accum_70__31_, prod_accum_70__30_, prod_accum_70__29_, prod_accum_70__28_, prod_accum_70__27_, prod_accum_70__26_, prod_accum_70__25_, prod_accum_70__24_, prod_accum_70__23_, prod_accum_70__22_, prod_accum_70__21_, prod_accum_70__20_, prod_accum_70__19_, prod_accum_70__18_, prod_accum_70__17_, prod_accum_70__16_, prod_accum_70__15_, prod_accum_70__14_, prod_accum_70__13_, prod_accum_70__12_, prod_accum_70__11_, prod_accum_70__10_, prod_accum_70__9_, prod_accum_70__8_, prod_accum_70__7_, prod_accum_70__6_, prod_accum_70__5_, prod_accum_70__4_, prod_accum_70__3_, prod_accum_70__2_, prod_accum_70__1_, prod_accum_70__0_ })
  );


  bsg_mul_array_row_128_71_x
  genblk1_71__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[9087:8960]),
    .b_i(b_r[9087:8960]),
    .s_i({ s_r_70__127_, s_r_70__126_, s_r_70__125_, s_r_70__124_, s_r_70__123_, s_r_70__122_, s_r_70__121_, s_r_70__120_, s_r_70__119_, s_r_70__118_, s_r_70__117_, s_r_70__116_, s_r_70__115_, s_r_70__114_, s_r_70__113_, s_r_70__112_, s_r_70__111_, s_r_70__110_, s_r_70__109_, s_r_70__108_, s_r_70__107_, s_r_70__106_, s_r_70__105_, s_r_70__104_, s_r_70__103_, s_r_70__102_, s_r_70__101_, s_r_70__100_, s_r_70__99_, s_r_70__98_, s_r_70__97_, s_r_70__96_, s_r_70__95_, s_r_70__94_, s_r_70__93_, s_r_70__92_, s_r_70__91_, s_r_70__90_, s_r_70__89_, s_r_70__88_, s_r_70__87_, s_r_70__86_, s_r_70__85_, s_r_70__84_, s_r_70__83_, s_r_70__82_, s_r_70__81_, s_r_70__80_, s_r_70__79_, s_r_70__78_, s_r_70__77_, s_r_70__76_, s_r_70__75_, s_r_70__74_, s_r_70__73_, s_r_70__72_, s_r_70__71_, s_r_70__70_, s_r_70__69_, s_r_70__68_, s_r_70__67_, s_r_70__66_, s_r_70__65_, s_r_70__64_, s_r_70__63_, s_r_70__62_, s_r_70__61_, s_r_70__60_, s_r_70__59_, s_r_70__58_, s_r_70__57_, s_r_70__56_, s_r_70__55_, s_r_70__54_, s_r_70__53_, s_r_70__52_, s_r_70__51_, s_r_70__50_, s_r_70__49_, s_r_70__48_, s_r_70__47_, s_r_70__46_, s_r_70__45_, s_r_70__44_, s_r_70__43_, s_r_70__42_, s_r_70__41_, s_r_70__40_, s_r_70__39_, s_r_70__38_, s_r_70__37_, s_r_70__36_, s_r_70__35_, s_r_70__34_, s_r_70__33_, s_r_70__32_, s_r_70__31_, s_r_70__30_, s_r_70__29_, s_r_70__28_, s_r_70__27_, s_r_70__26_, s_r_70__25_, s_r_70__24_, s_r_70__23_, s_r_70__22_, s_r_70__21_, s_r_70__20_, s_r_70__19_, s_r_70__18_, s_r_70__17_, s_r_70__16_, s_r_70__15_, s_r_70__14_, s_r_70__13_, s_r_70__12_, s_r_70__11_, s_r_70__10_, s_r_70__9_, s_r_70__8_, s_r_70__7_, s_r_70__6_, s_r_70__5_, s_r_70__4_, s_r_70__3_, s_r_70__2_, s_r_70__1_, s_r_70__0_ }),
    .c_i(c_r[70]),
    .prod_accum_i({ prod_accum_70__71_, prod_accum_70__70_, prod_accum_70__69_, prod_accum_70__68_, prod_accum_70__67_, prod_accum_70__66_, prod_accum_70__65_, prod_accum_70__64_, prod_accum_70__63_, prod_accum_70__62_, prod_accum_70__61_, prod_accum_70__60_, prod_accum_70__59_, prod_accum_70__58_, prod_accum_70__57_, prod_accum_70__56_, prod_accum_70__55_, prod_accum_70__54_, prod_accum_70__53_, prod_accum_70__52_, prod_accum_70__51_, prod_accum_70__50_, prod_accum_70__49_, prod_accum_70__48_, prod_accum_70__47_, prod_accum_70__46_, prod_accum_70__45_, prod_accum_70__44_, prod_accum_70__43_, prod_accum_70__42_, prod_accum_70__41_, prod_accum_70__40_, prod_accum_70__39_, prod_accum_70__38_, prod_accum_70__37_, prod_accum_70__36_, prod_accum_70__35_, prod_accum_70__34_, prod_accum_70__33_, prod_accum_70__32_, prod_accum_70__31_, prod_accum_70__30_, prod_accum_70__29_, prod_accum_70__28_, prod_accum_70__27_, prod_accum_70__26_, prod_accum_70__25_, prod_accum_70__24_, prod_accum_70__23_, prod_accum_70__22_, prod_accum_70__21_, prod_accum_70__20_, prod_accum_70__19_, prod_accum_70__18_, prod_accum_70__17_, prod_accum_70__16_, prod_accum_70__15_, prod_accum_70__14_, prod_accum_70__13_, prod_accum_70__12_, prod_accum_70__11_, prod_accum_70__10_, prod_accum_70__9_, prod_accum_70__8_, prod_accum_70__7_, prod_accum_70__6_, prod_accum_70__5_, prod_accum_70__4_, prod_accum_70__3_, prod_accum_70__2_, prod_accum_70__1_, prod_accum_70__0_ }),
    .a_o(a_r[9215:9088]),
    .b_o(b_r[9215:9088]),
    .s_o({ s_r_71__127_, s_r_71__126_, s_r_71__125_, s_r_71__124_, s_r_71__123_, s_r_71__122_, s_r_71__121_, s_r_71__120_, s_r_71__119_, s_r_71__118_, s_r_71__117_, s_r_71__116_, s_r_71__115_, s_r_71__114_, s_r_71__113_, s_r_71__112_, s_r_71__111_, s_r_71__110_, s_r_71__109_, s_r_71__108_, s_r_71__107_, s_r_71__106_, s_r_71__105_, s_r_71__104_, s_r_71__103_, s_r_71__102_, s_r_71__101_, s_r_71__100_, s_r_71__99_, s_r_71__98_, s_r_71__97_, s_r_71__96_, s_r_71__95_, s_r_71__94_, s_r_71__93_, s_r_71__92_, s_r_71__91_, s_r_71__90_, s_r_71__89_, s_r_71__88_, s_r_71__87_, s_r_71__86_, s_r_71__85_, s_r_71__84_, s_r_71__83_, s_r_71__82_, s_r_71__81_, s_r_71__80_, s_r_71__79_, s_r_71__78_, s_r_71__77_, s_r_71__76_, s_r_71__75_, s_r_71__74_, s_r_71__73_, s_r_71__72_, s_r_71__71_, s_r_71__70_, s_r_71__69_, s_r_71__68_, s_r_71__67_, s_r_71__66_, s_r_71__65_, s_r_71__64_, s_r_71__63_, s_r_71__62_, s_r_71__61_, s_r_71__60_, s_r_71__59_, s_r_71__58_, s_r_71__57_, s_r_71__56_, s_r_71__55_, s_r_71__54_, s_r_71__53_, s_r_71__52_, s_r_71__51_, s_r_71__50_, s_r_71__49_, s_r_71__48_, s_r_71__47_, s_r_71__46_, s_r_71__45_, s_r_71__44_, s_r_71__43_, s_r_71__42_, s_r_71__41_, s_r_71__40_, s_r_71__39_, s_r_71__38_, s_r_71__37_, s_r_71__36_, s_r_71__35_, s_r_71__34_, s_r_71__33_, s_r_71__32_, s_r_71__31_, s_r_71__30_, s_r_71__29_, s_r_71__28_, s_r_71__27_, s_r_71__26_, s_r_71__25_, s_r_71__24_, s_r_71__23_, s_r_71__22_, s_r_71__21_, s_r_71__20_, s_r_71__19_, s_r_71__18_, s_r_71__17_, s_r_71__16_, s_r_71__15_, s_r_71__14_, s_r_71__13_, s_r_71__12_, s_r_71__11_, s_r_71__10_, s_r_71__9_, s_r_71__8_, s_r_71__7_, s_r_71__6_, s_r_71__5_, s_r_71__4_, s_r_71__3_, s_r_71__2_, s_r_71__1_, s_r_71__0_ }),
    .c_o(c_r[71]),
    .prod_accum_o({ prod_accum_71__72_, prod_accum_71__71_, prod_accum_71__70_, prod_accum_71__69_, prod_accum_71__68_, prod_accum_71__67_, prod_accum_71__66_, prod_accum_71__65_, prod_accum_71__64_, prod_accum_71__63_, prod_accum_71__62_, prod_accum_71__61_, prod_accum_71__60_, prod_accum_71__59_, prod_accum_71__58_, prod_accum_71__57_, prod_accum_71__56_, prod_accum_71__55_, prod_accum_71__54_, prod_accum_71__53_, prod_accum_71__52_, prod_accum_71__51_, prod_accum_71__50_, prod_accum_71__49_, prod_accum_71__48_, prod_accum_71__47_, prod_accum_71__46_, prod_accum_71__45_, prod_accum_71__44_, prod_accum_71__43_, prod_accum_71__42_, prod_accum_71__41_, prod_accum_71__40_, prod_accum_71__39_, prod_accum_71__38_, prod_accum_71__37_, prod_accum_71__36_, prod_accum_71__35_, prod_accum_71__34_, prod_accum_71__33_, prod_accum_71__32_, prod_accum_71__31_, prod_accum_71__30_, prod_accum_71__29_, prod_accum_71__28_, prod_accum_71__27_, prod_accum_71__26_, prod_accum_71__25_, prod_accum_71__24_, prod_accum_71__23_, prod_accum_71__22_, prod_accum_71__21_, prod_accum_71__20_, prod_accum_71__19_, prod_accum_71__18_, prod_accum_71__17_, prod_accum_71__16_, prod_accum_71__15_, prod_accum_71__14_, prod_accum_71__13_, prod_accum_71__12_, prod_accum_71__11_, prod_accum_71__10_, prod_accum_71__9_, prod_accum_71__8_, prod_accum_71__7_, prod_accum_71__6_, prod_accum_71__5_, prod_accum_71__4_, prod_accum_71__3_, prod_accum_71__2_, prod_accum_71__1_, prod_accum_71__0_ })
  );


  bsg_mul_array_row_128_72_x
  genblk1_72__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[9215:9088]),
    .b_i(b_r[9215:9088]),
    .s_i({ s_r_71__127_, s_r_71__126_, s_r_71__125_, s_r_71__124_, s_r_71__123_, s_r_71__122_, s_r_71__121_, s_r_71__120_, s_r_71__119_, s_r_71__118_, s_r_71__117_, s_r_71__116_, s_r_71__115_, s_r_71__114_, s_r_71__113_, s_r_71__112_, s_r_71__111_, s_r_71__110_, s_r_71__109_, s_r_71__108_, s_r_71__107_, s_r_71__106_, s_r_71__105_, s_r_71__104_, s_r_71__103_, s_r_71__102_, s_r_71__101_, s_r_71__100_, s_r_71__99_, s_r_71__98_, s_r_71__97_, s_r_71__96_, s_r_71__95_, s_r_71__94_, s_r_71__93_, s_r_71__92_, s_r_71__91_, s_r_71__90_, s_r_71__89_, s_r_71__88_, s_r_71__87_, s_r_71__86_, s_r_71__85_, s_r_71__84_, s_r_71__83_, s_r_71__82_, s_r_71__81_, s_r_71__80_, s_r_71__79_, s_r_71__78_, s_r_71__77_, s_r_71__76_, s_r_71__75_, s_r_71__74_, s_r_71__73_, s_r_71__72_, s_r_71__71_, s_r_71__70_, s_r_71__69_, s_r_71__68_, s_r_71__67_, s_r_71__66_, s_r_71__65_, s_r_71__64_, s_r_71__63_, s_r_71__62_, s_r_71__61_, s_r_71__60_, s_r_71__59_, s_r_71__58_, s_r_71__57_, s_r_71__56_, s_r_71__55_, s_r_71__54_, s_r_71__53_, s_r_71__52_, s_r_71__51_, s_r_71__50_, s_r_71__49_, s_r_71__48_, s_r_71__47_, s_r_71__46_, s_r_71__45_, s_r_71__44_, s_r_71__43_, s_r_71__42_, s_r_71__41_, s_r_71__40_, s_r_71__39_, s_r_71__38_, s_r_71__37_, s_r_71__36_, s_r_71__35_, s_r_71__34_, s_r_71__33_, s_r_71__32_, s_r_71__31_, s_r_71__30_, s_r_71__29_, s_r_71__28_, s_r_71__27_, s_r_71__26_, s_r_71__25_, s_r_71__24_, s_r_71__23_, s_r_71__22_, s_r_71__21_, s_r_71__20_, s_r_71__19_, s_r_71__18_, s_r_71__17_, s_r_71__16_, s_r_71__15_, s_r_71__14_, s_r_71__13_, s_r_71__12_, s_r_71__11_, s_r_71__10_, s_r_71__9_, s_r_71__8_, s_r_71__7_, s_r_71__6_, s_r_71__5_, s_r_71__4_, s_r_71__3_, s_r_71__2_, s_r_71__1_, s_r_71__0_ }),
    .c_i(c_r[71]),
    .prod_accum_i({ prod_accum_71__72_, prod_accum_71__71_, prod_accum_71__70_, prod_accum_71__69_, prod_accum_71__68_, prod_accum_71__67_, prod_accum_71__66_, prod_accum_71__65_, prod_accum_71__64_, prod_accum_71__63_, prod_accum_71__62_, prod_accum_71__61_, prod_accum_71__60_, prod_accum_71__59_, prod_accum_71__58_, prod_accum_71__57_, prod_accum_71__56_, prod_accum_71__55_, prod_accum_71__54_, prod_accum_71__53_, prod_accum_71__52_, prod_accum_71__51_, prod_accum_71__50_, prod_accum_71__49_, prod_accum_71__48_, prod_accum_71__47_, prod_accum_71__46_, prod_accum_71__45_, prod_accum_71__44_, prod_accum_71__43_, prod_accum_71__42_, prod_accum_71__41_, prod_accum_71__40_, prod_accum_71__39_, prod_accum_71__38_, prod_accum_71__37_, prod_accum_71__36_, prod_accum_71__35_, prod_accum_71__34_, prod_accum_71__33_, prod_accum_71__32_, prod_accum_71__31_, prod_accum_71__30_, prod_accum_71__29_, prod_accum_71__28_, prod_accum_71__27_, prod_accum_71__26_, prod_accum_71__25_, prod_accum_71__24_, prod_accum_71__23_, prod_accum_71__22_, prod_accum_71__21_, prod_accum_71__20_, prod_accum_71__19_, prod_accum_71__18_, prod_accum_71__17_, prod_accum_71__16_, prod_accum_71__15_, prod_accum_71__14_, prod_accum_71__13_, prod_accum_71__12_, prod_accum_71__11_, prod_accum_71__10_, prod_accum_71__9_, prod_accum_71__8_, prod_accum_71__7_, prod_accum_71__6_, prod_accum_71__5_, prod_accum_71__4_, prod_accum_71__3_, prod_accum_71__2_, prod_accum_71__1_, prod_accum_71__0_ }),
    .a_o(a_r[9343:9216]),
    .b_o(b_r[9343:9216]),
    .s_o({ s_r_72__127_, s_r_72__126_, s_r_72__125_, s_r_72__124_, s_r_72__123_, s_r_72__122_, s_r_72__121_, s_r_72__120_, s_r_72__119_, s_r_72__118_, s_r_72__117_, s_r_72__116_, s_r_72__115_, s_r_72__114_, s_r_72__113_, s_r_72__112_, s_r_72__111_, s_r_72__110_, s_r_72__109_, s_r_72__108_, s_r_72__107_, s_r_72__106_, s_r_72__105_, s_r_72__104_, s_r_72__103_, s_r_72__102_, s_r_72__101_, s_r_72__100_, s_r_72__99_, s_r_72__98_, s_r_72__97_, s_r_72__96_, s_r_72__95_, s_r_72__94_, s_r_72__93_, s_r_72__92_, s_r_72__91_, s_r_72__90_, s_r_72__89_, s_r_72__88_, s_r_72__87_, s_r_72__86_, s_r_72__85_, s_r_72__84_, s_r_72__83_, s_r_72__82_, s_r_72__81_, s_r_72__80_, s_r_72__79_, s_r_72__78_, s_r_72__77_, s_r_72__76_, s_r_72__75_, s_r_72__74_, s_r_72__73_, s_r_72__72_, s_r_72__71_, s_r_72__70_, s_r_72__69_, s_r_72__68_, s_r_72__67_, s_r_72__66_, s_r_72__65_, s_r_72__64_, s_r_72__63_, s_r_72__62_, s_r_72__61_, s_r_72__60_, s_r_72__59_, s_r_72__58_, s_r_72__57_, s_r_72__56_, s_r_72__55_, s_r_72__54_, s_r_72__53_, s_r_72__52_, s_r_72__51_, s_r_72__50_, s_r_72__49_, s_r_72__48_, s_r_72__47_, s_r_72__46_, s_r_72__45_, s_r_72__44_, s_r_72__43_, s_r_72__42_, s_r_72__41_, s_r_72__40_, s_r_72__39_, s_r_72__38_, s_r_72__37_, s_r_72__36_, s_r_72__35_, s_r_72__34_, s_r_72__33_, s_r_72__32_, s_r_72__31_, s_r_72__30_, s_r_72__29_, s_r_72__28_, s_r_72__27_, s_r_72__26_, s_r_72__25_, s_r_72__24_, s_r_72__23_, s_r_72__22_, s_r_72__21_, s_r_72__20_, s_r_72__19_, s_r_72__18_, s_r_72__17_, s_r_72__16_, s_r_72__15_, s_r_72__14_, s_r_72__13_, s_r_72__12_, s_r_72__11_, s_r_72__10_, s_r_72__9_, s_r_72__8_, s_r_72__7_, s_r_72__6_, s_r_72__5_, s_r_72__4_, s_r_72__3_, s_r_72__2_, s_r_72__1_, s_r_72__0_ }),
    .c_o(c_r[72]),
    .prod_accum_o({ prod_accum_72__73_, prod_accum_72__72_, prod_accum_72__71_, prod_accum_72__70_, prod_accum_72__69_, prod_accum_72__68_, prod_accum_72__67_, prod_accum_72__66_, prod_accum_72__65_, prod_accum_72__64_, prod_accum_72__63_, prod_accum_72__62_, prod_accum_72__61_, prod_accum_72__60_, prod_accum_72__59_, prod_accum_72__58_, prod_accum_72__57_, prod_accum_72__56_, prod_accum_72__55_, prod_accum_72__54_, prod_accum_72__53_, prod_accum_72__52_, prod_accum_72__51_, prod_accum_72__50_, prod_accum_72__49_, prod_accum_72__48_, prod_accum_72__47_, prod_accum_72__46_, prod_accum_72__45_, prod_accum_72__44_, prod_accum_72__43_, prod_accum_72__42_, prod_accum_72__41_, prod_accum_72__40_, prod_accum_72__39_, prod_accum_72__38_, prod_accum_72__37_, prod_accum_72__36_, prod_accum_72__35_, prod_accum_72__34_, prod_accum_72__33_, prod_accum_72__32_, prod_accum_72__31_, prod_accum_72__30_, prod_accum_72__29_, prod_accum_72__28_, prod_accum_72__27_, prod_accum_72__26_, prod_accum_72__25_, prod_accum_72__24_, prod_accum_72__23_, prod_accum_72__22_, prod_accum_72__21_, prod_accum_72__20_, prod_accum_72__19_, prod_accum_72__18_, prod_accum_72__17_, prod_accum_72__16_, prod_accum_72__15_, prod_accum_72__14_, prod_accum_72__13_, prod_accum_72__12_, prod_accum_72__11_, prod_accum_72__10_, prod_accum_72__9_, prod_accum_72__8_, prod_accum_72__7_, prod_accum_72__6_, prod_accum_72__5_, prod_accum_72__4_, prod_accum_72__3_, prod_accum_72__2_, prod_accum_72__1_, prod_accum_72__0_ })
  );


  bsg_mul_array_row_128_73_x
  genblk1_73__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[9343:9216]),
    .b_i(b_r[9343:9216]),
    .s_i({ s_r_72__127_, s_r_72__126_, s_r_72__125_, s_r_72__124_, s_r_72__123_, s_r_72__122_, s_r_72__121_, s_r_72__120_, s_r_72__119_, s_r_72__118_, s_r_72__117_, s_r_72__116_, s_r_72__115_, s_r_72__114_, s_r_72__113_, s_r_72__112_, s_r_72__111_, s_r_72__110_, s_r_72__109_, s_r_72__108_, s_r_72__107_, s_r_72__106_, s_r_72__105_, s_r_72__104_, s_r_72__103_, s_r_72__102_, s_r_72__101_, s_r_72__100_, s_r_72__99_, s_r_72__98_, s_r_72__97_, s_r_72__96_, s_r_72__95_, s_r_72__94_, s_r_72__93_, s_r_72__92_, s_r_72__91_, s_r_72__90_, s_r_72__89_, s_r_72__88_, s_r_72__87_, s_r_72__86_, s_r_72__85_, s_r_72__84_, s_r_72__83_, s_r_72__82_, s_r_72__81_, s_r_72__80_, s_r_72__79_, s_r_72__78_, s_r_72__77_, s_r_72__76_, s_r_72__75_, s_r_72__74_, s_r_72__73_, s_r_72__72_, s_r_72__71_, s_r_72__70_, s_r_72__69_, s_r_72__68_, s_r_72__67_, s_r_72__66_, s_r_72__65_, s_r_72__64_, s_r_72__63_, s_r_72__62_, s_r_72__61_, s_r_72__60_, s_r_72__59_, s_r_72__58_, s_r_72__57_, s_r_72__56_, s_r_72__55_, s_r_72__54_, s_r_72__53_, s_r_72__52_, s_r_72__51_, s_r_72__50_, s_r_72__49_, s_r_72__48_, s_r_72__47_, s_r_72__46_, s_r_72__45_, s_r_72__44_, s_r_72__43_, s_r_72__42_, s_r_72__41_, s_r_72__40_, s_r_72__39_, s_r_72__38_, s_r_72__37_, s_r_72__36_, s_r_72__35_, s_r_72__34_, s_r_72__33_, s_r_72__32_, s_r_72__31_, s_r_72__30_, s_r_72__29_, s_r_72__28_, s_r_72__27_, s_r_72__26_, s_r_72__25_, s_r_72__24_, s_r_72__23_, s_r_72__22_, s_r_72__21_, s_r_72__20_, s_r_72__19_, s_r_72__18_, s_r_72__17_, s_r_72__16_, s_r_72__15_, s_r_72__14_, s_r_72__13_, s_r_72__12_, s_r_72__11_, s_r_72__10_, s_r_72__9_, s_r_72__8_, s_r_72__7_, s_r_72__6_, s_r_72__5_, s_r_72__4_, s_r_72__3_, s_r_72__2_, s_r_72__1_, s_r_72__0_ }),
    .c_i(c_r[72]),
    .prod_accum_i({ prod_accum_72__73_, prod_accum_72__72_, prod_accum_72__71_, prod_accum_72__70_, prod_accum_72__69_, prod_accum_72__68_, prod_accum_72__67_, prod_accum_72__66_, prod_accum_72__65_, prod_accum_72__64_, prod_accum_72__63_, prod_accum_72__62_, prod_accum_72__61_, prod_accum_72__60_, prod_accum_72__59_, prod_accum_72__58_, prod_accum_72__57_, prod_accum_72__56_, prod_accum_72__55_, prod_accum_72__54_, prod_accum_72__53_, prod_accum_72__52_, prod_accum_72__51_, prod_accum_72__50_, prod_accum_72__49_, prod_accum_72__48_, prod_accum_72__47_, prod_accum_72__46_, prod_accum_72__45_, prod_accum_72__44_, prod_accum_72__43_, prod_accum_72__42_, prod_accum_72__41_, prod_accum_72__40_, prod_accum_72__39_, prod_accum_72__38_, prod_accum_72__37_, prod_accum_72__36_, prod_accum_72__35_, prod_accum_72__34_, prod_accum_72__33_, prod_accum_72__32_, prod_accum_72__31_, prod_accum_72__30_, prod_accum_72__29_, prod_accum_72__28_, prod_accum_72__27_, prod_accum_72__26_, prod_accum_72__25_, prod_accum_72__24_, prod_accum_72__23_, prod_accum_72__22_, prod_accum_72__21_, prod_accum_72__20_, prod_accum_72__19_, prod_accum_72__18_, prod_accum_72__17_, prod_accum_72__16_, prod_accum_72__15_, prod_accum_72__14_, prod_accum_72__13_, prod_accum_72__12_, prod_accum_72__11_, prod_accum_72__10_, prod_accum_72__9_, prod_accum_72__8_, prod_accum_72__7_, prod_accum_72__6_, prod_accum_72__5_, prod_accum_72__4_, prod_accum_72__3_, prod_accum_72__2_, prod_accum_72__1_, prod_accum_72__0_ }),
    .a_o(a_r[9471:9344]),
    .b_o(b_r[9471:9344]),
    .s_o({ s_r_73__127_, s_r_73__126_, s_r_73__125_, s_r_73__124_, s_r_73__123_, s_r_73__122_, s_r_73__121_, s_r_73__120_, s_r_73__119_, s_r_73__118_, s_r_73__117_, s_r_73__116_, s_r_73__115_, s_r_73__114_, s_r_73__113_, s_r_73__112_, s_r_73__111_, s_r_73__110_, s_r_73__109_, s_r_73__108_, s_r_73__107_, s_r_73__106_, s_r_73__105_, s_r_73__104_, s_r_73__103_, s_r_73__102_, s_r_73__101_, s_r_73__100_, s_r_73__99_, s_r_73__98_, s_r_73__97_, s_r_73__96_, s_r_73__95_, s_r_73__94_, s_r_73__93_, s_r_73__92_, s_r_73__91_, s_r_73__90_, s_r_73__89_, s_r_73__88_, s_r_73__87_, s_r_73__86_, s_r_73__85_, s_r_73__84_, s_r_73__83_, s_r_73__82_, s_r_73__81_, s_r_73__80_, s_r_73__79_, s_r_73__78_, s_r_73__77_, s_r_73__76_, s_r_73__75_, s_r_73__74_, s_r_73__73_, s_r_73__72_, s_r_73__71_, s_r_73__70_, s_r_73__69_, s_r_73__68_, s_r_73__67_, s_r_73__66_, s_r_73__65_, s_r_73__64_, s_r_73__63_, s_r_73__62_, s_r_73__61_, s_r_73__60_, s_r_73__59_, s_r_73__58_, s_r_73__57_, s_r_73__56_, s_r_73__55_, s_r_73__54_, s_r_73__53_, s_r_73__52_, s_r_73__51_, s_r_73__50_, s_r_73__49_, s_r_73__48_, s_r_73__47_, s_r_73__46_, s_r_73__45_, s_r_73__44_, s_r_73__43_, s_r_73__42_, s_r_73__41_, s_r_73__40_, s_r_73__39_, s_r_73__38_, s_r_73__37_, s_r_73__36_, s_r_73__35_, s_r_73__34_, s_r_73__33_, s_r_73__32_, s_r_73__31_, s_r_73__30_, s_r_73__29_, s_r_73__28_, s_r_73__27_, s_r_73__26_, s_r_73__25_, s_r_73__24_, s_r_73__23_, s_r_73__22_, s_r_73__21_, s_r_73__20_, s_r_73__19_, s_r_73__18_, s_r_73__17_, s_r_73__16_, s_r_73__15_, s_r_73__14_, s_r_73__13_, s_r_73__12_, s_r_73__11_, s_r_73__10_, s_r_73__9_, s_r_73__8_, s_r_73__7_, s_r_73__6_, s_r_73__5_, s_r_73__4_, s_r_73__3_, s_r_73__2_, s_r_73__1_, s_r_73__0_ }),
    .c_o(c_r[73]),
    .prod_accum_o({ prod_accum_73__74_, prod_accum_73__73_, prod_accum_73__72_, prod_accum_73__71_, prod_accum_73__70_, prod_accum_73__69_, prod_accum_73__68_, prod_accum_73__67_, prod_accum_73__66_, prod_accum_73__65_, prod_accum_73__64_, prod_accum_73__63_, prod_accum_73__62_, prod_accum_73__61_, prod_accum_73__60_, prod_accum_73__59_, prod_accum_73__58_, prod_accum_73__57_, prod_accum_73__56_, prod_accum_73__55_, prod_accum_73__54_, prod_accum_73__53_, prod_accum_73__52_, prod_accum_73__51_, prod_accum_73__50_, prod_accum_73__49_, prod_accum_73__48_, prod_accum_73__47_, prod_accum_73__46_, prod_accum_73__45_, prod_accum_73__44_, prod_accum_73__43_, prod_accum_73__42_, prod_accum_73__41_, prod_accum_73__40_, prod_accum_73__39_, prod_accum_73__38_, prod_accum_73__37_, prod_accum_73__36_, prod_accum_73__35_, prod_accum_73__34_, prod_accum_73__33_, prod_accum_73__32_, prod_accum_73__31_, prod_accum_73__30_, prod_accum_73__29_, prod_accum_73__28_, prod_accum_73__27_, prod_accum_73__26_, prod_accum_73__25_, prod_accum_73__24_, prod_accum_73__23_, prod_accum_73__22_, prod_accum_73__21_, prod_accum_73__20_, prod_accum_73__19_, prod_accum_73__18_, prod_accum_73__17_, prod_accum_73__16_, prod_accum_73__15_, prod_accum_73__14_, prod_accum_73__13_, prod_accum_73__12_, prod_accum_73__11_, prod_accum_73__10_, prod_accum_73__9_, prod_accum_73__8_, prod_accum_73__7_, prod_accum_73__6_, prod_accum_73__5_, prod_accum_73__4_, prod_accum_73__3_, prod_accum_73__2_, prod_accum_73__1_, prod_accum_73__0_ })
  );


  bsg_mul_array_row_128_74_x
  genblk1_74__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[9471:9344]),
    .b_i(b_r[9471:9344]),
    .s_i({ s_r_73__127_, s_r_73__126_, s_r_73__125_, s_r_73__124_, s_r_73__123_, s_r_73__122_, s_r_73__121_, s_r_73__120_, s_r_73__119_, s_r_73__118_, s_r_73__117_, s_r_73__116_, s_r_73__115_, s_r_73__114_, s_r_73__113_, s_r_73__112_, s_r_73__111_, s_r_73__110_, s_r_73__109_, s_r_73__108_, s_r_73__107_, s_r_73__106_, s_r_73__105_, s_r_73__104_, s_r_73__103_, s_r_73__102_, s_r_73__101_, s_r_73__100_, s_r_73__99_, s_r_73__98_, s_r_73__97_, s_r_73__96_, s_r_73__95_, s_r_73__94_, s_r_73__93_, s_r_73__92_, s_r_73__91_, s_r_73__90_, s_r_73__89_, s_r_73__88_, s_r_73__87_, s_r_73__86_, s_r_73__85_, s_r_73__84_, s_r_73__83_, s_r_73__82_, s_r_73__81_, s_r_73__80_, s_r_73__79_, s_r_73__78_, s_r_73__77_, s_r_73__76_, s_r_73__75_, s_r_73__74_, s_r_73__73_, s_r_73__72_, s_r_73__71_, s_r_73__70_, s_r_73__69_, s_r_73__68_, s_r_73__67_, s_r_73__66_, s_r_73__65_, s_r_73__64_, s_r_73__63_, s_r_73__62_, s_r_73__61_, s_r_73__60_, s_r_73__59_, s_r_73__58_, s_r_73__57_, s_r_73__56_, s_r_73__55_, s_r_73__54_, s_r_73__53_, s_r_73__52_, s_r_73__51_, s_r_73__50_, s_r_73__49_, s_r_73__48_, s_r_73__47_, s_r_73__46_, s_r_73__45_, s_r_73__44_, s_r_73__43_, s_r_73__42_, s_r_73__41_, s_r_73__40_, s_r_73__39_, s_r_73__38_, s_r_73__37_, s_r_73__36_, s_r_73__35_, s_r_73__34_, s_r_73__33_, s_r_73__32_, s_r_73__31_, s_r_73__30_, s_r_73__29_, s_r_73__28_, s_r_73__27_, s_r_73__26_, s_r_73__25_, s_r_73__24_, s_r_73__23_, s_r_73__22_, s_r_73__21_, s_r_73__20_, s_r_73__19_, s_r_73__18_, s_r_73__17_, s_r_73__16_, s_r_73__15_, s_r_73__14_, s_r_73__13_, s_r_73__12_, s_r_73__11_, s_r_73__10_, s_r_73__9_, s_r_73__8_, s_r_73__7_, s_r_73__6_, s_r_73__5_, s_r_73__4_, s_r_73__3_, s_r_73__2_, s_r_73__1_, s_r_73__0_ }),
    .c_i(c_r[73]),
    .prod_accum_i({ prod_accum_73__74_, prod_accum_73__73_, prod_accum_73__72_, prod_accum_73__71_, prod_accum_73__70_, prod_accum_73__69_, prod_accum_73__68_, prod_accum_73__67_, prod_accum_73__66_, prod_accum_73__65_, prod_accum_73__64_, prod_accum_73__63_, prod_accum_73__62_, prod_accum_73__61_, prod_accum_73__60_, prod_accum_73__59_, prod_accum_73__58_, prod_accum_73__57_, prod_accum_73__56_, prod_accum_73__55_, prod_accum_73__54_, prod_accum_73__53_, prod_accum_73__52_, prod_accum_73__51_, prod_accum_73__50_, prod_accum_73__49_, prod_accum_73__48_, prod_accum_73__47_, prod_accum_73__46_, prod_accum_73__45_, prod_accum_73__44_, prod_accum_73__43_, prod_accum_73__42_, prod_accum_73__41_, prod_accum_73__40_, prod_accum_73__39_, prod_accum_73__38_, prod_accum_73__37_, prod_accum_73__36_, prod_accum_73__35_, prod_accum_73__34_, prod_accum_73__33_, prod_accum_73__32_, prod_accum_73__31_, prod_accum_73__30_, prod_accum_73__29_, prod_accum_73__28_, prod_accum_73__27_, prod_accum_73__26_, prod_accum_73__25_, prod_accum_73__24_, prod_accum_73__23_, prod_accum_73__22_, prod_accum_73__21_, prod_accum_73__20_, prod_accum_73__19_, prod_accum_73__18_, prod_accum_73__17_, prod_accum_73__16_, prod_accum_73__15_, prod_accum_73__14_, prod_accum_73__13_, prod_accum_73__12_, prod_accum_73__11_, prod_accum_73__10_, prod_accum_73__9_, prod_accum_73__8_, prod_accum_73__7_, prod_accum_73__6_, prod_accum_73__5_, prod_accum_73__4_, prod_accum_73__3_, prod_accum_73__2_, prod_accum_73__1_, prod_accum_73__0_ }),
    .a_o(a_r[9599:9472]),
    .b_o(b_r[9599:9472]),
    .s_o({ s_r_74__127_, s_r_74__126_, s_r_74__125_, s_r_74__124_, s_r_74__123_, s_r_74__122_, s_r_74__121_, s_r_74__120_, s_r_74__119_, s_r_74__118_, s_r_74__117_, s_r_74__116_, s_r_74__115_, s_r_74__114_, s_r_74__113_, s_r_74__112_, s_r_74__111_, s_r_74__110_, s_r_74__109_, s_r_74__108_, s_r_74__107_, s_r_74__106_, s_r_74__105_, s_r_74__104_, s_r_74__103_, s_r_74__102_, s_r_74__101_, s_r_74__100_, s_r_74__99_, s_r_74__98_, s_r_74__97_, s_r_74__96_, s_r_74__95_, s_r_74__94_, s_r_74__93_, s_r_74__92_, s_r_74__91_, s_r_74__90_, s_r_74__89_, s_r_74__88_, s_r_74__87_, s_r_74__86_, s_r_74__85_, s_r_74__84_, s_r_74__83_, s_r_74__82_, s_r_74__81_, s_r_74__80_, s_r_74__79_, s_r_74__78_, s_r_74__77_, s_r_74__76_, s_r_74__75_, s_r_74__74_, s_r_74__73_, s_r_74__72_, s_r_74__71_, s_r_74__70_, s_r_74__69_, s_r_74__68_, s_r_74__67_, s_r_74__66_, s_r_74__65_, s_r_74__64_, s_r_74__63_, s_r_74__62_, s_r_74__61_, s_r_74__60_, s_r_74__59_, s_r_74__58_, s_r_74__57_, s_r_74__56_, s_r_74__55_, s_r_74__54_, s_r_74__53_, s_r_74__52_, s_r_74__51_, s_r_74__50_, s_r_74__49_, s_r_74__48_, s_r_74__47_, s_r_74__46_, s_r_74__45_, s_r_74__44_, s_r_74__43_, s_r_74__42_, s_r_74__41_, s_r_74__40_, s_r_74__39_, s_r_74__38_, s_r_74__37_, s_r_74__36_, s_r_74__35_, s_r_74__34_, s_r_74__33_, s_r_74__32_, s_r_74__31_, s_r_74__30_, s_r_74__29_, s_r_74__28_, s_r_74__27_, s_r_74__26_, s_r_74__25_, s_r_74__24_, s_r_74__23_, s_r_74__22_, s_r_74__21_, s_r_74__20_, s_r_74__19_, s_r_74__18_, s_r_74__17_, s_r_74__16_, s_r_74__15_, s_r_74__14_, s_r_74__13_, s_r_74__12_, s_r_74__11_, s_r_74__10_, s_r_74__9_, s_r_74__8_, s_r_74__7_, s_r_74__6_, s_r_74__5_, s_r_74__4_, s_r_74__3_, s_r_74__2_, s_r_74__1_, s_r_74__0_ }),
    .c_o(c_r[74]),
    .prod_accum_o({ prod_accum_74__75_, prod_accum_74__74_, prod_accum_74__73_, prod_accum_74__72_, prod_accum_74__71_, prod_accum_74__70_, prod_accum_74__69_, prod_accum_74__68_, prod_accum_74__67_, prod_accum_74__66_, prod_accum_74__65_, prod_accum_74__64_, prod_accum_74__63_, prod_accum_74__62_, prod_accum_74__61_, prod_accum_74__60_, prod_accum_74__59_, prod_accum_74__58_, prod_accum_74__57_, prod_accum_74__56_, prod_accum_74__55_, prod_accum_74__54_, prod_accum_74__53_, prod_accum_74__52_, prod_accum_74__51_, prod_accum_74__50_, prod_accum_74__49_, prod_accum_74__48_, prod_accum_74__47_, prod_accum_74__46_, prod_accum_74__45_, prod_accum_74__44_, prod_accum_74__43_, prod_accum_74__42_, prod_accum_74__41_, prod_accum_74__40_, prod_accum_74__39_, prod_accum_74__38_, prod_accum_74__37_, prod_accum_74__36_, prod_accum_74__35_, prod_accum_74__34_, prod_accum_74__33_, prod_accum_74__32_, prod_accum_74__31_, prod_accum_74__30_, prod_accum_74__29_, prod_accum_74__28_, prod_accum_74__27_, prod_accum_74__26_, prod_accum_74__25_, prod_accum_74__24_, prod_accum_74__23_, prod_accum_74__22_, prod_accum_74__21_, prod_accum_74__20_, prod_accum_74__19_, prod_accum_74__18_, prod_accum_74__17_, prod_accum_74__16_, prod_accum_74__15_, prod_accum_74__14_, prod_accum_74__13_, prod_accum_74__12_, prod_accum_74__11_, prod_accum_74__10_, prod_accum_74__9_, prod_accum_74__8_, prod_accum_74__7_, prod_accum_74__6_, prod_accum_74__5_, prod_accum_74__4_, prod_accum_74__3_, prod_accum_74__2_, prod_accum_74__1_, prod_accum_74__0_ })
  );


  bsg_mul_array_row_128_75_x
  genblk1_75__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[9599:9472]),
    .b_i(b_r[9599:9472]),
    .s_i({ s_r_74__127_, s_r_74__126_, s_r_74__125_, s_r_74__124_, s_r_74__123_, s_r_74__122_, s_r_74__121_, s_r_74__120_, s_r_74__119_, s_r_74__118_, s_r_74__117_, s_r_74__116_, s_r_74__115_, s_r_74__114_, s_r_74__113_, s_r_74__112_, s_r_74__111_, s_r_74__110_, s_r_74__109_, s_r_74__108_, s_r_74__107_, s_r_74__106_, s_r_74__105_, s_r_74__104_, s_r_74__103_, s_r_74__102_, s_r_74__101_, s_r_74__100_, s_r_74__99_, s_r_74__98_, s_r_74__97_, s_r_74__96_, s_r_74__95_, s_r_74__94_, s_r_74__93_, s_r_74__92_, s_r_74__91_, s_r_74__90_, s_r_74__89_, s_r_74__88_, s_r_74__87_, s_r_74__86_, s_r_74__85_, s_r_74__84_, s_r_74__83_, s_r_74__82_, s_r_74__81_, s_r_74__80_, s_r_74__79_, s_r_74__78_, s_r_74__77_, s_r_74__76_, s_r_74__75_, s_r_74__74_, s_r_74__73_, s_r_74__72_, s_r_74__71_, s_r_74__70_, s_r_74__69_, s_r_74__68_, s_r_74__67_, s_r_74__66_, s_r_74__65_, s_r_74__64_, s_r_74__63_, s_r_74__62_, s_r_74__61_, s_r_74__60_, s_r_74__59_, s_r_74__58_, s_r_74__57_, s_r_74__56_, s_r_74__55_, s_r_74__54_, s_r_74__53_, s_r_74__52_, s_r_74__51_, s_r_74__50_, s_r_74__49_, s_r_74__48_, s_r_74__47_, s_r_74__46_, s_r_74__45_, s_r_74__44_, s_r_74__43_, s_r_74__42_, s_r_74__41_, s_r_74__40_, s_r_74__39_, s_r_74__38_, s_r_74__37_, s_r_74__36_, s_r_74__35_, s_r_74__34_, s_r_74__33_, s_r_74__32_, s_r_74__31_, s_r_74__30_, s_r_74__29_, s_r_74__28_, s_r_74__27_, s_r_74__26_, s_r_74__25_, s_r_74__24_, s_r_74__23_, s_r_74__22_, s_r_74__21_, s_r_74__20_, s_r_74__19_, s_r_74__18_, s_r_74__17_, s_r_74__16_, s_r_74__15_, s_r_74__14_, s_r_74__13_, s_r_74__12_, s_r_74__11_, s_r_74__10_, s_r_74__9_, s_r_74__8_, s_r_74__7_, s_r_74__6_, s_r_74__5_, s_r_74__4_, s_r_74__3_, s_r_74__2_, s_r_74__1_, s_r_74__0_ }),
    .c_i(c_r[74]),
    .prod_accum_i({ prod_accum_74__75_, prod_accum_74__74_, prod_accum_74__73_, prod_accum_74__72_, prod_accum_74__71_, prod_accum_74__70_, prod_accum_74__69_, prod_accum_74__68_, prod_accum_74__67_, prod_accum_74__66_, prod_accum_74__65_, prod_accum_74__64_, prod_accum_74__63_, prod_accum_74__62_, prod_accum_74__61_, prod_accum_74__60_, prod_accum_74__59_, prod_accum_74__58_, prod_accum_74__57_, prod_accum_74__56_, prod_accum_74__55_, prod_accum_74__54_, prod_accum_74__53_, prod_accum_74__52_, prod_accum_74__51_, prod_accum_74__50_, prod_accum_74__49_, prod_accum_74__48_, prod_accum_74__47_, prod_accum_74__46_, prod_accum_74__45_, prod_accum_74__44_, prod_accum_74__43_, prod_accum_74__42_, prod_accum_74__41_, prod_accum_74__40_, prod_accum_74__39_, prod_accum_74__38_, prod_accum_74__37_, prod_accum_74__36_, prod_accum_74__35_, prod_accum_74__34_, prod_accum_74__33_, prod_accum_74__32_, prod_accum_74__31_, prod_accum_74__30_, prod_accum_74__29_, prod_accum_74__28_, prod_accum_74__27_, prod_accum_74__26_, prod_accum_74__25_, prod_accum_74__24_, prod_accum_74__23_, prod_accum_74__22_, prod_accum_74__21_, prod_accum_74__20_, prod_accum_74__19_, prod_accum_74__18_, prod_accum_74__17_, prod_accum_74__16_, prod_accum_74__15_, prod_accum_74__14_, prod_accum_74__13_, prod_accum_74__12_, prod_accum_74__11_, prod_accum_74__10_, prod_accum_74__9_, prod_accum_74__8_, prod_accum_74__7_, prod_accum_74__6_, prod_accum_74__5_, prod_accum_74__4_, prod_accum_74__3_, prod_accum_74__2_, prod_accum_74__1_, prod_accum_74__0_ }),
    .a_o(a_r[9727:9600]),
    .b_o(b_r[9727:9600]),
    .s_o({ s_r_75__127_, s_r_75__126_, s_r_75__125_, s_r_75__124_, s_r_75__123_, s_r_75__122_, s_r_75__121_, s_r_75__120_, s_r_75__119_, s_r_75__118_, s_r_75__117_, s_r_75__116_, s_r_75__115_, s_r_75__114_, s_r_75__113_, s_r_75__112_, s_r_75__111_, s_r_75__110_, s_r_75__109_, s_r_75__108_, s_r_75__107_, s_r_75__106_, s_r_75__105_, s_r_75__104_, s_r_75__103_, s_r_75__102_, s_r_75__101_, s_r_75__100_, s_r_75__99_, s_r_75__98_, s_r_75__97_, s_r_75__96_, s_r_75__95_, s_r_75__94_, s_r_75__93_, s_r_75__92_, s_r_75__91_, s_r_75__90_, s_r_75__89_, s_r_75__88_, s_r_75__87_, s_r_75__86_, s_r_75__85_, s_r_75__84_, s_r_75__83_, s_r_75__82_, s_r_75__81_, s_r_75__80_, s_r_75__79_, s_r_75__78_, s_r_75__77_, s_r_75__76_, s_r_75__75_, s_r_75__74_, s_r_75__73_, s_r_75__72_, s_r_75__71_, s_r_75__70_, s_r_75__69_, s_r_75__68_, s_r_75__67_, s_r_75__66_, s_r_75__65_, s_r_75__64_, s_r_75__63_, s_r_75__62_, s_r_75__61_, s_r_75__60_, s_r_75__59_, s_r_75__58_, s_r_75__57_, s_r_75__56_, s_r_75__55_, s_r_75__54_, s_r_75__53_, s_r_75__52_, s_r_75__51_, s_r_75__50_, s_r_75__49_, s_r_75__48_, s_r_75__47_, s_r_75__46_, s_r_75__45_, s_r_75__44_, s_r_75__43_, s_r_75__42_, s_r_75__41_, s_r_75__40_, s_r_75__39_, s_r_75__38_, s_r_75__37_, s_r_75__36_, s_r_75__35_, s_r_75__34_, s_r_75__33_, s_r_75__32_, s_r_75__31_, s_r_75__30_, s_r_75__29_, s_r_75__28_, s_r_75__27_, s_r_75__26_, s_r_75__25_, s_r_75__24_, s_r_75__23_, s_r_75__22_, s_r_75__21_, s_r_75__20_, s_r_75__19_, s_r_75__18_, s_r_75__17_, s_r_75__16_, s_r_75__15_, s_r_75__14_, s_r_75__13_, s_r_75__12_, s_r_75__11_, s_r_75__10_, s_r_75__9_, s_r_75__8_, s_r_75__7_, s_r_75__6_, s_r_75__5_, s_r_75__4_, s_r_75__3_, s_r_75__2_, s_r_75__1_, s_r_75__0_ }),
    .c_o(c_r[75]),
    .prod_accum_o({ prod_accum_75__76_, prod_accum_75__75_, prod_accum_75__74_, prod_accum_75__73_, prod_accum_75__72_, prod_accum_75__71_, prod_accum_75__70_, prod_accum_75__69_, prod_accum_75__68_, prod_accum_75__67_, prod_accum_75__66_, prod_accum_75__65_, prod_accum_75__64_, prod_accum_75__63_, prod_accum_75__62_, prod_accum_75__61_, prod_accum_75__60_, prod_accum_75__59_, prod_accum_75__58_, prod_accum_75__57_, prod_accum_75__56_, prod_accum_75__55_, prod_accum_75__54_, prod_accum_75__53_, prod_accum_75__52_, prod_accum_75__51_, prod_accum_75__50_, prod_accum_75__49_, prod_accum_75__48_, prod_accum_75__47_, prod_accum_75__46_, prod_accum_75__45_, prod_accum_75__44_, prod_accum_75__43_, prod_accum_75__42_, prod_accum_75__41_, prod_accum_75__40_, prod_accum_75__39_, prod_accum_75__38_, prod_accum_75__37_, prod_accum_75__36_, prod_accum_75__35_, prod_accum_75__34_, prod_accum_75__33_, prod_accum_75__32_, prod_accum_75__31_, prod_accum_75__30_, prod_accum_75__29_, prod_accum_75__28_, prod_accum_75__27_, prod_accum_75__26_, prod_accum_75__25_, prod_accum_75__24_, prod_accum_75__23_, prod_accum_75__22_, prod_accum_75__21_, prod_accum_75__20_, prod_accum_75__19_, prod_accum_75__18_, prod_accum_75__17_, prod_accum_75__16_, prod_accum_75__15_, prod_accum_75__14_, prod_accum_75__13_, prod_accum_75__12_, prod_accum_75__11_, prod_accum_75__10_, prod_accum_75__9_, prod_accum_75__8_, prod_accum_75__7_, prod_accum_75__6_, prod_accum_75__5_, prod_accum_75__4_, prod_accum_75__3_, prod_accum_75__2_, prod_accum_75__1_, prod_accum_75__0_ })
  );


  bsg_mul_array_row_128_76_x
  genblk1_76__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[9727:9600]),
    .b_i(b_r[9727:9600]),
    .s_i({ s_r_75__127_, s_r_75__126_, s_r_75__125_, s_r_75__124_, s_r_75__123_, s_r_75__122_, s_r_75__121_, s_r_75__120_, s_r_75__119_, s_r_75__118_, s_r_75__117_, s_r_75__116_, s_r_75__115_, s_r_75__114_, s_r_75__113_, s_r_75__112_, s_r_75__111_, s_r_75__110_, s_r_75__109_, s_r_75__108_, s_r_75__107_, s_r_75__106_, s_r_75__105_, s_r_75__104_, s_r_75__103_, s_r_75__102_, s_r_75__101_, s_r_75__100_, s_r_75__99_, s_r_75__98_, s_r_75__97_, s_r_75__96_, s_r_75__95_, s_r_75__94_, s_r_75__93_, s_r_75__92_, s_r_75__91_, s_r_75__90_, s_r_75__89_, s_r_75__88_, s_r_75__87_, s_r_75__86_, s_r_75__85_, s_r_75__84_, s_r_75__83_, s_r_75__82_, s_r_75__81_, s_r_75__80_, s_r_75__79_, s_r_75__78_, s_r_75__77_, s_r_75__76_, s_r_75__75_, s_r_75__74_, s_r_75__73_, s_r_75__72_, s_r_75__71_, s_r_75__70_, s_r_75__69_, s_r_75__68_, s_r_75__67_, s_r_75__66_, s_r_75__65_, s_r_75__64_, s_r_75__63_, s_r_75__62_, s_r_75__61_, s_r_75__60_, s_r_75__59_, s_r_75__58_, s_r_75__57_, s_r_75__56_, s_r_75__55_, s_r_75__54_, s_r_75__53_, s_r_75__52_, s_r_75__51_, s_r_75__50_, s_r_75__49_, s_r_75__48_, s_r_75__47_, s_r_75__46_, s_r_75__45_, s_r_75__44_, s_r_75__43_, s_r_75__42_, s_r_75__41_, s_r_75__40_, s_r_75__39_, s_r_75__38_, s_r_75__37_, s_r_75__36_, s_r_75__35_, s_r_75__34_, s_r_75__33_, s_r_75__32_, s_r_75__31_, s_r_75__30_, s_r_75__29_, s_r_75__28_, s_r_75__27_, s_r_75__26_, s_r_75__25_, s_r_75__24_, s_r_75__23_, s_r_75__22_, s_r_75__21_, s_r_75__20_, s_r_75__19_, s_r_75__18_, s_r_75__17_, s_r_75__16_, s_r_75__15_, s_r_75__14_, s_r_75__13_, s_r_75__12_, s_r_75__11_, s_r_75__10_, s_r_75__9_, s_r_75__8_, s_r_75__7_, s_r_75__6_, s_r_75__5_, s_r_75__4_, s_r_75__3_, s_r_75__2_, s_r_75__1_, s_r_75__0_ }),
    .c_i(c_r[75]),
    .prod_accum_i({ prod_accum_75__76_, prod_accum_75__75_, prod_accum_75__74_, prod_accum_75__73_, prod_accum_75__72_, prod_accum_75__71_, prod_accum_75__70_, prod_accum_75__69_, prod_accum_75__68_, prod_accum_75__67_, prod_accum_75__66_, prod_accum_75__65_, prod_accum_75__64_, prod_accum_75__63_, prod_accum_75__62_, prod_accum_75__61_, prod_accum_75__60_, prod_accum_75__59_, prod_accum_75__58_, prod_accum_75__57_, prod_accum_75__56_, prod_accum_75__55_, prod_accum_75__54_, prod_accum_75__53_, prod_accum_75__52_, prod_accum_75__51_, prod_accum_75__50_, prod_accum_75__49_, prod_accum_75__48_, prod_accum_75__47_, prod_accum_75__46_, prod_accum_75__45_, prod_accum_75__44_, prod_accum_75__43_, prod_accum_75__42_, prod_accum_75__41_, prod_accum_75__40_, prod_accum_75__39_, prod_accum_75__38_, prod_accum_75__37_, prod_accum_75__36_, prod_accum_75__35_, prod_accum_75__34_, prod_accum_75__33_, prod_accum_75__32_, prod_accum_75__31_, prod_accum_75__30_, prod_accum_75__29_, prod_accum_75__28_, prod_accum_75__27_, prod_accum_75__26_, prod_accum_75__25_, prod_accum_75__24_, prod_accum_75__23_, prod_accum_75__22_, prod_accum_75__21_, prod_accum_75__20_, prod_accum_75__19_, prod_accum_75__18_, prod_accum_75__17_, prod_accum_75__16_, prod_accum_75__15_, prod_accum_75__14_, prod_accum_75__13_, prod_accum_75__12_, prod_accum_75__11_, prod_accum_75__10_, prod_accum_75__9_, prod_accum_75__8_, prod_accum_75__7_, prod_accum_75__6_, prod_accum_75__5_, prod_accum_75__4_, prod_accum_75__3_, prod_accum_75__2_, prod_accum_75__1_, prod_accum_75__0_ }),
    .a_o(a_r[9855:9728]),
    .b_o(b_r[9855:9728]),
    .s_o({ s_r_76__127_, s_r_76__126_, s_r_76__125_, s_r_76__124_, s_r_76__123_, s_r_76__122_, s_r_76__121_, s_r_76__120_, s_r_76__119_, s_r_76__118_, s_r_76__117_, s_r_76__116_, s_r_76__115_, s_r_76__114_, s_r_76__113_, s_r_76__112_, s_r_76__111_, s_r_76__110_, s_r_76__109_, s_r_76__108_, s_r_76__107_, s_r_76__106_, s_r_76__105_, s_r_76__104_, s_r_76__103_, s_r_76__102_, s_r_76__101_, s_r_76__100_, s_r_76__99_, s_r_76__98_, s_r_76__97_, s_r_76__96_, s_r_76__95_, s_r_76__94_, s_r_76__93_, s_r_76__92_, s_r_76__91_, s_r_76__90_, s_r_76__89_, s_r_76__88_, s_r_76__87_, s_r_76__86_, s_r_76__85_, s_r_76__84_, s_r_76__83_, s_r_76__82_, s_r_76__81_, s_r_76__80_, s_r_76__79_, s_r_76__78_, s_r_76__77_, s_r_76__76_, s_r_76__75_, s_r_76__74_, s_r_76__73_, s_r_76__72_, s_r_76__71_, s_r_76__70_, s_r_76__69_, s_r_76__68_, s_r_76__67_, s_r_76__66_, s_r_76__65_, s_r_76__64_, s_r_76__63_, s_r_76__62_, s_r_76__61_, s_r_76__60_, s_r_76__59_, s_r_76__58_, s_r_76__57_, s_r_76__56_, s_r_76__55_, s_r_76__54_, s_r_76__53_, s_r_76__52_, s_r_76__51_, s_r_76__50_, s_r_76__49_, s_r_76__48_, s_r_76__47_, s_r_76__46_, s_r_76__45_, s_r_76__44_, s_r_76__43_, s_r_76__42_, s_r_76__41_, s_r_76__40_, s_r_76__39_, s_r_76__38_, s_r_76__37_, s_r_76__36_, s_r_76__35_, s_r_76__34_, s_r_76__33_, s_r_76__32_, s_r_76__31_, s_r_76__30_, s_r_76__29_, s_r_76__28_, s_r_76__27_, s_r_76__26_, s_r_76__25_, s_r_76__24_, s_r_76__23_, s_r_76__22_, s_r_76__21_, s_r_76__20_, s_r_76__19_, s_r_76__18_, s_r_76__17_, s_r_76__16_, s_r_76__15_, s_r_76__14_, s_r_76__13_, s_r_76__12_, s_r_76__11_, s_r_76__10_, s_r_76__9_, s_r_76__8_, s_r_76__7_, s_r_76__6_, s_r_76__5_, s_r_76__4_, s_r_76__3_, s_r_76__2_, s_r_76__1_, s_r_76__0_ }),
    .c_o(c_r[76]),
    .prod_accum_o({ prod_accum_76__77_, prod_accum_76__76_, prod_accum_76__75_, prod_accum_76__74_, prod_accum_76__73_, prod_accum_76__72_, prod_accum_76__71_, prod_accum_76__70_, prod_accum_76__69_, prod_accum_76__68_, prod_accum_76__67_, prod_accum_76__66_, prod_accum_76__65_, prod_accum_76__64_, prod_accum_76__63_, prod_accum_76__62_, prod_accum_76__61_, prod_accum_76__60_, prod_accum_76__59_, prod_accum_76__58_, prod_accum_76__57_, prod_accum_76__56_, prod_accum_76__55_, prod_accum_76__54_, prod_accum_76__53_, prod_accum_76__52_, prod_accum_76__51_, prod_accum_76__50_, prod_accum_76__49_, prod_accum_76__48_, prod_accum_76__47_, prod_accum_76__46_, prod_accum_76__45_, prod_accum_76__44_, prod_accum_76__43_, prod_accum_76__42_, prod_accum_76__41_, prod_accum_76__40_, prod_accum_76__39_, prod_accum_76__38_, prod_accum_76__37_, prod_accum_76__36_, prod_accum_76__35_, prod_accum_76__34_, prod_accum_76__33_, prod_accum_76__32_, prod_accum_76__31_, prod_accum_76__30_, prod_accum_76__29_, prod_accum_76__28_, prod_accum_76__27_, prod_accum_76__26_, prod_accum_76__25_, prod_accum_76__24_, prod_accum_76__23_, prod_accum_76__22_, prod_accum_76__21_, prod_accum_76__20_, prod_accum_76__19_, prod_accum_76__18_, prod_accum_76__17_, prod_accum_76__16_, prod_accum_76__15_, prod_accum_76__14_, prod_accum_76__13_, prod_accum_76__12_, prod_accum_76__11_, prod_accum_76__10_, prod_accum_76__9_, prod_accum_76__8_, prod_accum_76__7_, prod_accum_76__6_, prod_accum_76__5_, prod_accum_76__4_, prod_accum_76__3_, prod_accum_76__2_, prod_accum_76__1_, prod_accum_76__0_ })
  );


  bsg_mul_array_row_128_77_x
  genblk1_77__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[9855:9728]),
    .b_i(b_r[9855:9728]),
    .s_i({ s_r_76__127_, s_r_76__126_, s_r_76__125_, s_r_76__124_, s_r_76__123_, s_r_76__122_, s_r_76__121_, s_r_76__120_, s_r_76__119_, s_r_76__118_, s_r_76__117_, s_r_76__116_, s_r_76__115_, s_r_76__114_, s_r_76__113_, s_r_76__112_, s_r_76__111_, s_r_76__110_, s_r_76__109_, s_r_76__108_, s_r_76__107_, s_r_76__106_, s_r_76__105_, s_r_76__104_, s_r_76__103_, s_r_76__102_, s_r_76__101_, s_r_76__100_, s_r_76__99_, s_r_76__98_, s_r_76__97_, s_r_76__96_, s_r_76__95_, s_r_76__94_, s_r_76__93_, s_r_76__92_, s_r_76__91_, s_r_76__90_, s_r_76__89_, s_r_76__88_, s_r_76__87_, s_r_76__86_, s_r_76__85_, s_r_76__84_, s_r_76__83_, s_r_76__82_, s_r_76__81_, s_r_76__80_, s_r_76__79_, s_r_76__78_, s_r_76__77_, s_r_76__76_, s_r_76__75_, s_r_76__74_, s_r_76__73_, s_r_76__72_, s_r_76__71_, s_r_76__70_, s_r_76__69_, s_r_76__68_, s_r_76__67_, s_r_76__66_, s_r_76__65_, s_r_76__64_, s_r_76__63_, s_r_76__62_, s_r_76__61_, s_r_76__60_, s_r_76__59_, s_r_76__58_, s_r_76__57_, s_r_76__56_, s_r_76__55_, s_r_76__54_, s_r_76__53_, s_r_76__52_, s_r_76__51_, s_r_76__50_, s_r_76__49_, s_r_76__48_, s_r_76__47_, s_r_76__46_, s_r_76__45_, s_r_76__44_, s_r_76__43_, s_r_76__42_, s_r_76__41_, s_r_76__40_, s_r_76__39_, s_r_76__38_, s_r_76__37_, s_r_76__36_, s_r_76__35_, s_r_76__34_, s_r_76__33_, s_r_76__32_, s_r_76__31_, s_r_76__30_, s_r_76__29_, s_r_76__28_, s_r_76__27_, s_r_76__26_, s_r_76__25_, s_r_76__24_, s_r_76__23_, s_r_76__22_, s_r_76__21_, s_r_76__20_, s_r_76__19_, s_r_76__18_, s_r_76__17_, s_r_76__16_, s_r_76__15_, s_r_76__14_, s_r_76__13_, s_r_76__12_, s_r_76__11_, s_r_76__10_, s_r_76__9_, s_r_76__8_, s_r_76__7_, s_r_76__6_, s_r_76__5_, s_r_76__4_, s_r_76__3_, s_r_76__2_, s_r_76__1_, s_r_76__0_ }),
    .c_i(c_r[76]),
    .prod_accum_i({ prod_accum_76__77_, prod_accum_76__76_, prod_accum_76__75_, prod_accum_76__74_, prod_accum_76__73_, prod_accum_76__72_, prod_accum_76__71_, prod_accum_76__70_, prod_accum_76__69_, prod_accum_76__68_, prod_accum_76__67_, prod_accum_76__66_, prod_accum_76__65_, prod_accum_76__64_, prod_accum_76__63_, prod_accum_76__62_, prod_accum_76__61_, prod_accum_76__60_, prod_accum_76__59_, prod_accum_76__58_, prod_accum_76__57_, prod_accum_76__56_, prod_accum_76__55_, prod_accum_76__54_, prod_accum_76__53_, prod_accum_76__52_, prod_accum_76__51_, prod_accum_76__50_, prod_accum_76__49_, prod_accum_76__48_, prod_accum_76__47_, prod_accum_76__46_, prod_accum_76__45_, prod_accum_76__44_, prod_accum_76__43_, prod_accum_76__42_, prod_accum_76__41_, prod_accum_76__40_, prod_accum_76__39_, prod_accum_76__38_, prod_accum_76__37_, prod_accum_76__36_, prod_accum_76__35_, prod_accum_76__34_, prod_accum_76__33_, prod_accum_76__32_, prod_accum_76__31_, prod_accum_76__30_, prod_accum_76__29_, prod_accum_76__28_, prod_accum_76__27_, prod_accum_76__26_, prod_accum_76__25_, prod_accum_76__24_, prod_accum_76__23_, prod_accum_76__22_, prod_accum_76__21_, prod_accum_76__20_, prod_accum_76__19_, prod_accum_76__18_, prod_accum_76__17_, prod_accum_76__16_, prod_accum_76__15_, prod_accum_76__14_, prod_accum_76__13_, prod_accum_76__12_, prod_accum_76__11_, prod_accum_76__10_, prod_accum_76__9_, prod_accum_76__8_, prod_accum_76__7_, prod_accum_76__6_, prod_accum_76__5_, prod_accum_76__4_, prod_accum_76__3_, prod_accum_76__2_, prod_accum_76__1_, prod_accum_76__0_ }),
    .a_o(a_r[9983:9856]),
    .b_o(b_r[9983:9856]),
    .s_o({ s_r_77__127_, s_r_77__126_, s_r_77__125_, s_r_77__124_, s_r_77__123_, s_r_77__122_, s_r_77__121_, s_r_77__120_, s_r_77__119_, s_r_77__118_, s_r_77__117_, s_r_77__116_, s_r_77__115_, s_r_77__114_, s_r_77__113_, s_r_77__112_, s_r_77__111_, s_r_77__110_, s_r_77__109_, s_r_77__108_, s_r_77__107_, s_r_77__106_, s_r_77__105_, s_r_77__104_, s_r_77__103_, s_r_77__102_, s_r_77__101_, s_r_77__100_, s_r_77__99_, s_r_77__98_, s_r_77__97_, s_r_77__96_, s_r_77__95_, s_r_77__94_, s_r_77__93_, s_r_77__92_, s_r_77__91_, s_r_77__90_, s_r_77__89_, s_r_77__88_, s_r_77__87_, s_r_77__86_, s_r_77__85_, s_r_77__84_, s_r_77__83_, s_r_77__82_, s_r_77__81_, s_r_77__80_, s_r_77__79_, s_r_77__78_, s_r_77__77_, s_r_77__76_, s_r_77__75_, s_r_77__74_, s_r_77__73_, s_r_77__72_, s_r_77__71_, s_r_77__70_, s_r_77__69_, s_r_77__68_, s_r_77__67_, s_r_77__66_, s_r_77__65_, s_r_77__64_, s_r_77__63_, s_r_77__62_, s_r_77__61_, s_r_77__60_, s_r_77__59_, s_r_77__58_, s_r_77__57_, s_r_77__56_, s_r_77__55_, s_r_77__54_, s_r_77__53_, s_r_77__52_, s_r_77__51_, s_r_77__50_, s_r_77__49_, s_r_77__48_, s_r_77__47_, s_r_77__46_, s_r_77__45_, s_r_77__44_, s_r_77__43_, s_r_77__42_, s_r_77__41_, s_r_77__40_, s_r_77__39_, s_r_77__38_, s_r_77__37_, s_r_77__36_, s_r_77__35_, s_r_77__34_, s_r_77__33_, s_r_77__32_, s_r_77__31_, s_r_77__30_, s_r_77__29_, s_r_77__28_, s_r_77__27_, s_r_77__26_, s_r_77__25_, s_r_77__24_, s_r_77__23_, s_r_77__22_, s_r_77__21_, s_r_77__20_, s_r_77__19_, s_r_77__18_, s_r_77__17_, s_r_77__16_, s_r_77__15_, s_r_77__14_, s_r_77__13_, s_r_77__12_, s_r_77__11_, s_r_77__10_, s_r_77__9_, s_r_77__8_, s_r_77__7_, s_r_77__6_, s_r_77__5_, s_r_77__4_, s_r_77__3_, s_r_77__2_, s_r_77__1_, s_r_77__0_ }),
    .c_o(c_r[77]),
    .prod_accum_o({ prod_accum_77__78_, prod_accum_77__77_, prod_accum_77__76_, prod_accum_77__75_, prod_accum_77__74_, prod_accum_77__73_, prod_accum_77__72_, prod_accum_77__71_, prod_accum_77__70_, prod_accum_77__69_, prod_accum_77__68_, prod_accum_77__67_, prod_accum_77__66_, prod_accum_77__65_, prod_accum_77__64_, prod_accum_77__63_, prod_accum_77__62_, prod_accum_77__61_, prod_accum_77__60_, prod_accum_77__59_, prod_accum_77__58_, prod_accum_77__57_, prod_accum_77__56_, prod_accum_77__55_, prod_accum_77__54_, prod_accum_77__53_, prod_accum_77__52_, prod_accum_77__51_, prod_accum_77__50_, prod_accum_77__49_, prod_accum_77__48_, prod_accum_77__47_, prod_accum_77__46_, prod_accum_77__45_, prod_accum_77__44_, prod_accum_77__43_, prod_accum_77__42_, prod_accum_77__41_, prod_accum_77__40_, prod_accum_77__39_, prod_accum_77__38_, prod_accum_77__37_, prod_accum_77__36_, prod_accum_77__35_, prod_accum_77__34_, prod_accum_77__33_, prod_accum_77__32_, prod_accum_77__31_, prod_accum_77__30_, prod_accum_77__29_, prod_accum_77__28_, prod_accum_77__27_, prod_accum_77__26_, prod_accum_77__25_, prod_accum_77__24_, prod_accum_77__23_, prod_accum_77__22_, prod_accum_77__21_, prod_accum_77__20_, prod_accum_77__19_, prod_accum_77__18_, prod_accum_77__17_, prod_accum_77__16_, prod_accum_77__15_, prod_accum_77__14_, prod_accum_77__13_, prod_accum_77__12_, prod_accum_77__11_, prod_accum_77__10_, prod_accum_77__9_, prod_accum_77__8_, prod_accum_77__7_, prod_accum_77__6_, prod_accum_77__5_, prod_accum_77__4_, prod_accum_77__3_, prod_accum_77__2_, prod_accum_77__1_, prod_accum_77__0_ })
  );


  bsg_mul_array_row_128_78_x
  genblk1_78__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[9983:9856]),
    .b_i(b_r[9983:9856]),
    .s_i({ s_r_77__127_, s_r_77__126_, s_r_77__125_, s_r_77__124_, s_r_77__123_, s_r_77__122_, s_r_77__121_, s_r_77__120_, s_r_77__119_, s_r_77__118_, s_r_77__117_, s_r_77__116_, s_r_77__115_, s_r_77__114_, s_r_77__113_, s_r_77__112_, s_r_77__111_, s_r_77__110_, s_r_77__109_, s_r_77__108_, s_r_77__107_, s_r_77__106_, s_r_77__105_, s_r_77__104_, s_r_77__103_, s_r_77__102_, s_r_77__101_, s_r_77__100_, s_r_77__99_, s_r_77__98_, s_r_77__97_, s_r_77__96_, s_r_77__95_, s_r_77__94_, s_r_77__93_, s_r_77__92_, s_r_77__91_, s_r_77__90_, s_r_77__89_, s_r_77__88_, s_r_77__87_, s_r_77__86_, s_r_77__85_, s_r_77__84_, s_r_77__83_, s_r_77__82_, s_r_77__81_, s_r_77__80_, s_r_77__79_, s_r_77__78_, s_r_77__77_, s_r_77__76_, s_r_77__75_, s_r_77__74_, s_r_77__73_, s_r_77__72_, s_r_77__71_, s_r_77__70_, s_r_77__69_, s_r_77__68_, s_r_77__67_, s_r_77__66_, s_r_77__65_, s_r_77__64_, s_r_77__63_, s_r_77__62_, s_r_77__61_, s_r_77__60_, s_r_77__59_, s_r_77__58_, s_r_77__57_, s_r_77__56_, s_r_77__55_, s_r_77__54_, s_r_77__53_, s_r_77__52_, s_r_77__51_, s_r_77__50_, s_r_77__49_, s_r_77__48_, s_r_77__47_, s_r_77__46_, s_r_77__45_, s_r_77__44_, s_r_77__43_, s_r_77__42_, s_r_77__41_, s_r_77__40_, s_r_77__39_, s_r_77__38_, s_r_77__37_, s_r_77__36_, s_r_77__35_, s_r_77__34_, s_r_77__33_, s_r_77__32_, s_r_77__31_, s_r_77__30_, s_r_77__29_, s_r_77__28_, s_r_77__27_, s_r_77__26_, s_r_77__25_, s_r_77__24_, s_r_77__23_, s_r_77__22_, s_r_77__21_, s_r_77__20_, s_r_77__19_, s_r_77__18_, s_r_77__17_, s_r_77__16_, s_r_77__15_, s_r_77__14_, s_r_77__13_, s_r_77__12_, s_r_77__11_, s_r_77__10_, s_r_77__9_, s_r_77__8_, s_r_77__7_, s_r_77__6_, s_r_77__5_, s_r_77__4_, s_r_77__3_, s_r_77__2_, s_r_77__1_, s_r_77__0_ }),
    .c_i(c_r[77]),
    .prod_accum_i({ prod_accum_77__78_, prod_accum_77__77_, prod_accum_77__76_, prod_accum_77__75_, prod_accum_77__74_, prod_accum_77__73_, prod_accum_77__72_, prod_accum_77__71_, prod_accum_77__70_, prod_accum_77__69_, prod_accum_77__68_, prod_accum_77__67_, prod_accum_77__66_, prod_accum_77__65_, prod_accum_77__64_, prod_accum_77__63_, prod_accum_77__62_, prod_accum_77__61_, prod_accum_77__60_, prod_accum_77__59_, prod_accum_77__58_, prod_accum_77__57_, prod_accum_77__56_, prod_accum_77__55_, prod_accum_77__54_, prod_accum_77__53_, prod_accum_77__52_, prod_accum_77__51_, prod_accum_77__50_, prod_accum_77__49_, prod_accum_77__48_, prod_accum_77__47_, prod_accum_77__46_, prod_accum_77__45_, prod_accum_77__44_, prod_accum_77__43_, prod_accum_77__42_, prod_accum_77__41_, prod_accum_77__40_, prod_accum_77__39_, prod_accum_77__38_, prod_accum_77__37_, prod_accum_77__36_, prod_accum_77__35_, prod_accum_77__34_, prod_accum_77__33_, prod_accum_77__32_, prod_accum_77__31_, prod_accum_77__30_, prod_accum_77__29_, prod_accum_77__28_, prod_accum_77__27_, prod_accum_77__26_, prod_accum_77__25_, prod_accum_77__24_, prod_accum_77__23_, prod_accum_77__22_, prod_accum_77__21_, prod_accum_77__20_, prod_accum_77__19_, prod_accum_77__18_, prod_accum_77__17_, prod_accum_77__16_, prod_accum_77__15_, prod_accum_77__14_, prod_accum_77__13_, prod_accum_77__12_, prod_accum_77__11_, prod_accum_77__10_, prod_accum_77__9_, prod_accum_77__8_, prod_accum_77__7_, prod_accum_77__6_, prod_accum_77__5_, prod_accum_77__4_, prod_accum_77__3_, prod_accum_77__2_, prod_accum_77__1_, prod_accum_77__0_ }),
    .a_o(a_r[10111:9984]),
    .b_o(b_r[10111:9984]),
    .s_o({ s_r_78__127_, s_r_78__126_, s_r_78__125_, s_r_78__124_, s_r_78__123_, s_r_78__122_, s_r_78__121_, s_r_78__120_, s_r_78__119_, s_r_78__118_, s_r_78__117_, s_r_78__116_, s_r_78__115_, s_r_78__114_, s_r_78__113_, s_r_78__112_, s_r_78__111_, s_r_78__110_, s_r_78__109_, s_r_78__108_, s_r_78__107_, s_r_78__106_, s_r_78__105_, s_r_78__104_, s_r_78__103_, s_r_78__102_, s_r_78__101_, s_r_78__100_, s_r_78__99_, s_r_78__98_, s_r_78__97_, s_r_78__96_, s_r_78__95_, s_r_78__94_, s_r_78__93_, s_r_78__92_, s_r_78__91_, s_r_78__90_, s_r_78__89_, s_r_78__88_, s_r_78__87_, s_r_78__86_, s_r_78__85_, s_r_78__84_, s_r_78__83_, s_r_78__82_, s_r_78__81_, s_r_78__80_, s_r_78__79_, s_r_78__78_, s_r_78__77_, s_r_78__76_, s_r_78__75_, s_r_78__74_, s_r_78__73_, s_r_78__72_, s_r_78__71_, s_r_78__70_, s_r_78__69_, s_r_78__68_, s_r_78__67_, s_r_78__66_, s_r_78__65_, s_r_78__64_, s_r_78__63_, s_r_78__62_, s_r_78__61_, s_r_78__60_, s_r_78__59_, s_r_78__58_, s_r_78__57_, s_r_78__56_, s_r_78__55_, s_r_78__54_, s_r_78__53_, s_r_78__52_, s_r_78__51_, s_r_78__50_, s_r_78__49_, s_r_78__48_, s_r_78__47_, s_r_78__46_, s_r_78__45_, s_r_78__44_, s_r_78__43_, s_r_78__42_, s_r_78__41_, s_r_78__40_, s_r_78__39_, s_r_78__38_, s_r_78__37_, s_r_78__36_, s_r_78__35_, s_r_78__34_, s_r_78__33_, s_r_78__32_, s_r_78__31_, s_r_78__30_, s_r_78__29_, s_r_78__28_, s_r_78__27_, s_r_78__26_, s_r_78__25_, s_r_78__24_, s_r_78__23_, s_r_78__22_, s_r_78__21_, s_r_78__20_, s_r_78__19_, s_r_78__18_, s_r_78__17_, s_r_78__16_, s_r_78__15_, s_r_78__14_, s_r_78__13_, s_r_78__12_, s_r_78__11_, s_r_78__10_, s_r_78__9_, s_r_78__8_, s_r_78__7_, s_r_78__6_, s_r_78__5_, s_r_78__4_, s_r_78__3_, s_r_78__2_, s_r_78__1_, s_r_78__0_ }),
    .c_o(c_r[78]),
    .prod_accum_o({ prod_accum_78__79_, prod_accum_78__78_, prod_accum_78__77_, prod_accum_78__76_, prod_accum_78__75_, prod_accum_78__74_, prod_accum_78__73_, prod_accum_78__72_, prod_accum_78__71_, prod_accum_78__70_, prod_accum_78__69_, prod_accum_78__68_, prod_accum_78__67_, prod_accum_78__66_, prod_accum_78__65_, prod_accum_78__64_, prod_accum_78__63_, prod_accum_78__62_, prod_accum_78__61_, prod_accum_78__60_, prod_accum_78__59_, prod_accum_78__58_, prod_accum_78__57_, prod_accum_78__56_, prod_accum_78__55_, prod_accum_78__54_, prod_accum_78__53_, prod_accum_78__52_, prod_accum_78__51_, prod_accum_78__50_, prod_accum_78__49_, prod_accum_78__48_, prod_accum_78__47_, prod_accum_78__46_, prod_accum_78__45_, prod_accum_78__44_, prod_accum_78__43_, prod_accum_78__42_, prod_accum_78__41_, prod_accum_78__40_, prod_accum_78__39_, prod_accum_78__38_, prod_accum_78__37_, prod_accum_78__36_, prod_accum_78__35_, prod_accum_78__34_, prod_accum_78__33_, prod_accum_78__32_, prod_accum_78__31_, prod_accum_78__30_, prod_accum_78__29_, prod_accum_78__28_, prod_accum_78__27_, prod_accum_78__26_, prod_accum_78__25_, prod_accum_78__24_, prod_accum_78__23_, prod_accum_78__22_, prod_accum_78__21_, prod_accum_78__20_, prod_accum_78__19_, prod_accum_78__18_, prod_accum_78__17_, prod_accum_78__16_, prod_accum_78__15_, prod_accum_78__14_, prod_accum_78__13_, prod_accum_78__12_, prod_accum_78__11_, prod_accum_78__10_, prod_accum_78__9_, prod_accum_78__8_, prod_accum_78__7_, prod_accum_78__6_, prod_accum_78__5_, prod_accum_78__4_, prod_accum_78__3_, prod_accum_78__2_, prod_accum_78__1_, prod_accum_78__0_ })
  );


  bsg_mul_array_row_128_79_x
  genblk1_79__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[10111:9984]),
    .b_i(b_r[10111:9984]),
    .s_i({ s_r_78__127_, s_r_78__126_, s_r_78__125_, s_r_78__124_, s_r_78__123_, s_r_78__122_, s_r_78__121_, s_r_78__120_, s_r_78__119_, s_r_78__118_, s_r_78__117_, s_r_78__116_, s_r_78__115_, s_r_78__114_, s_r_78__113_, s_r_78__112_, s_r_78__111_, s_r_78__110_, s_r_78__109_, s_r_78__108_, s_r_78__107_, s_r_78__106_, s_r_78__105_, s_r_78__104_, s_r_78__103_, s_r_78__102_, s_r_78__101_, s_r_78__100_, s_r_78__99_, s_r_78__98_, s_r_78__97_, s_r_78__96_, s_r_78__95_, s_r_78__94_, s_r_78__93_, s_r_78__92_, s_r_78__91_, s_r_78__90_, s_r_78__89_, s_r_78__88_, s_r_78__87_, s_r_78__86_, s_r_78__85_, s_r_78__84_, s_r_78__83_, s_r_78__82_, s_r_78__81_, s_r_78__80_, s_r_78__79_, s_r_78__78_, s_r_78__77_, s_r_78__76_, s_r_78__75_, s_r_78__74_, s_r_78__73_, s_r_78__72_, s_r_78__71_, s_r_78__70_, s_r_78__69_, s_r_78__68_, s_r_78__67_, s_r_78__66_, s_r_78__65_, s_r_78__64_, s_r_78__63_, s_r_78__62_, s_r_78__61_, s_r_78__60_, s_r_78__59_, s_r_78__58_, s_r_78__57_, s_r_78__56_, s_r_78__55_, s_r_78__54_, s_r_78__53_, s_r_78__52_, s_r_78__51_, s_r_78__50_, s_r_78__49_, s_r_78__48_, s_r_78__47_, s_r_78__46_, s_r_78__45_, s_r_78__44_, s_r_78__43_, s_r_78__42_, s_r_78__41_, s_r_78__40_, s_r_78__39_, s_r_78__38_, s_r_78__37_, s_r_78__36_, s_r_78__35_, s_r_78__34_, s_r_78__33_, s_r_78__32_, s_r_78__31_, s_r_78__30_, s_r_78__29_, s_r_78__28_, s_r_78__27_, s_r_78__26_, s_r_78__25_, s_r_78__24_, s_r_78__23_, s_r_78__22_, s_r_78__21_, s_r_78__20_, s_r_78__19_, s_r_78__18_, s_r_78__17_, s_r_78__16_, s_r_78__15_, s_r_78__14_, s_r_78__13_, s_r_78__12_, s_r_78__11_, s_r_78__10_, s_r_78__9_, s_r_78__8_, s_r_78__7_, s_r_78__6_, s_r_78__5_, s_r_78__4_, s_r_78__3_, s_r_78__2_, s_r_78__1_, s_r_78__0_ }),
    .c_i(c_r[78]),
    .prod_accum_i({ prod_accum_78__79_, prod_accum_78__78_, prod_accum_78__77_, prod_accum_78__76_, prod_accum_78__75_, prod_accum_78__74_, prod_accum_78__73_, prod_accum_78__72_, prod_accum_78__71_, prod_accum_78__70_, prod_accum_78__69_, prod_accum_78__68_, prod_accum_78__67_, prod_accum_78__66_, prod_accum_78__65_, prod_accum_78__64_, prod_accum_78__63_, prod_accum_78__62_, prod_accum_78__61_, prod_accum_78__60_, prod_accum_78__59_, prod_accum_78__58_, prod_accum_78__57_, prod_accum_78__56_, prod_accum_78__55_, prod_accum_78__54_, prod_accum_78__53_, prod_accum_78__52_, prod_accum_78__51_, prod_accum_78__50_, prod_accum_78__49_, prod_accum_78__48_, prod_accum_78__47_, prod_accum_78__46_, prod_accum_78__45_, prod_accum_78__44_, prod_accum_78__43_, prod_accum_78__42_, prod_accum_78__41_, prod_accum_78__40_, prod_accum_78__39_, prod_accum_78__38_, prod_accum_78__37_, prod_accum_78__36_, prod_accum_78__35_, prod_accum_78__34_, prod_accum_78__33_, prod_accum_78__32_, prod_accum_78__31_, prod_accum_78__30_, prod_accum_78__29_, prod_accum_78__28_, prod_accum_78__27_, prod_accum_78__26_, prod_accum_78__25_, prod_accum_78__24_, prod_accum_78__23_, prod_accum_78__22_, prod_accum_78__21_, prod_accum_78__20_, prod_accum_78__19_, prod_accum_78__18_, prod_accum_78__17_, prod_accum_78__16_, prod_accum_78__15_, prod_accum_78__14_, prod_accum_78__13_, prod_accum_78__12_, prod_accum_78__11_, prod_accum_78__10_, prod_accum_78__9_, prod_accum_78__8_, prod_accum_78__7_, prod_accum_78__6_, prod_accum_78__5_, prod_accum_78__4_, prod_accum_78__3_, prod_accum_78__2_, prod_accum_78__1_, prod_accum_78__0_ }),
    .a_o(a_r[10239:10112]),
    .b_o(b_r[10239:10112]),
    .s_o({ s_r_79__127_, s_r_79__126_, s_r_79__125_, s_r_79__124_, s_r_79__123_, s_r_79__122_, s_r_79__121_, s_r_79__120_, s_r_79__119_, s_r_79__118_, s_r_79__117_, s_r_79__116_, s_r_79__115_, s_r_79__114_, s_r_79__113_, s_r_79__112_, s_r_79__111_, s_r_79__110_, s_r_79__109_, s_r_79__108_, s_r_79__107_, s_r_79__106_, s_r_79__105_, s_r_79__104_, s_r_79__103_, s_r_79__102_, s_r_79__101_, s_r_79__100_, s_r_79__99_, s_r_79__98_, s_r_79__97_, s_r_79__96_, s_r_79__95_, s_r_79__94_, s_r_79__93_, s_r_79__92_, s_r_79__91_, s_r_79__90_, s_r_79__89_, s_r_79__88_, s_r_79__87_, s_r_79__86_, s_r_79__85_, s_r_79__84_, s_r_79__83_, s_r_79__82_, s_r_79__81_, s_r_79__80_, s_r_79__79_, s_r_79__78_, s_r_79__77_, s_r_79__76_, s_r_79__75_, s_r_79__74_, s_r_79__73_, s_r_79__72_, s_r_79__71_, s_r_79__70_, s_r_79__69_, s_r_79__68_, s_r_79__67_, s_r_79__66_, s_r_79__65_, s_r_79__64_, s_r_79__63_, s_r_79__62_, s_r_79__61_, s_r_79__60_, s_r_79__59_, s_r_79__58_, s_r_79__57_, s_r_79__56_, s_r_79__55_, s_r_79__54_, s_r_79__53_, s_r_79__52_, s_r_79__51_, s_r_79__50_, s_r_79__49_, s_r_79__48_, s_r_79__47_, s_r_79__46_, s_r_79__45_, s_r_79__44_, s_r_79__43_, s_r_79__42_, s_r_79__41_, s_r_79__40_, s_r_79__39_, s_r_79__38_, s_r_79__37_, s_r_79__36_, s_r_79__35_, s_r_79__34_, s_r_79__33_, s_r_79__32_, s_r_79__31_, s_r_79__30_, s_r_79__29_, s_r_79__28_, s_r_79__27_, s_r_79__26_, s_r_79__25_, s_r_79__24_, s_r_79__23_, s_r_79__22_, s_r_79__21_, s_r_79__20_, s_r_79__19_, s_r_79__18_, s_r_79__17_, s_r_79__16_, s_r_79__15_, s_r_79__14_, s_r_79__13_, s_r_79__12_, s_r_79__11_, s_r_79__10_, s_r_79__9_, s_r_79__8_, s_r_79__7_, s_r_79__6_, s_r_79__5_, s_r_79__4_, s_r_79__3_, s_r_79__2_, s_r_79__1_, s_r_79__0_ }),
    .c_o(c_r[79]),
    .prod_accum_o({ prod_accum_79__80_, prod_accum_79__79_, prod_accum_79__78_, prod_accum_79__77_, prod_accum_79__76_, prod_accum_79__75_, prod_accum_79__74_, prod_accum_79__73_, prod_accum_79__72_, prod_accum_79__71_, prod_accum_79__70_, prod_accum_79__69_, prod_accum_79__68_, prod_accum_79__67_, prod_accum_79__66_, prod_accum_79__65_, prod_accum_79__64_, prod_accum_79__63_, prod_accum_79__62_, prod_accum_79__61_, prod_accum_79__60_, prod_accum_79__59_, prod_accum_79__58_, prod_accum_79__57_, prod_accum_79__56_, prod_accum_79__55_, prod_accum_79__54_, prod_accum_79__53_, prod_accum_79__52_, prod_accum_79__51_, prod_accum_79__50_, prod_accum_79__49_, prod_accum_79__48_, prod_accum_79__47_, prod_accum_79__46_, prod_accum_79__45_, prod_accum_79__44_, prod_accum_79__43_, prod_accum_79__42_, prod_accum_79__41_, prod_accum_79__40_, prod_accum_79__39_, prod_accum_79__38_, prod_accum_79__37_, prod_accum_79__36_, prod_accum_79__35_, prod_accum_79__34_, prod_accum_79__33_, prod_accum_79__32_, prod_accum_79__31_, prod_accum_79__30_, prod_accum_79__29_, prod_accum_79__28_, prod_accum_79__27_, prod_accum_79__26_, prod_accum_79__25_, prod_accum_79__24_, prod_accum_79__23_, prod_accum_79__22_, prod_accum_79__21_, prod_accum_79__20_, prod_accum_79__19_, prod_accum_79__18_, prod_accum_79__17_, prod_accum_79__16_, prod_accum_79__15_, prod_accum_79__14_, prod_accum_79__13_, prod_accum_79__12_, prod_accum_79__11_, prod_accum_79__10_, prod_accum_79__9_, prod_accum_79__8_, prod_accum_79__7_, prod_accum_79__6_, prod_accum_79__5_, prod_accum_79__4_, prod_accum_79__3_, prod_accum_79__2_, prod_accum_79__1_, prod_accum_79__0_ })
  );


  bsg_mul_array_row_128_80_x
  genblk1_80__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[10239:10112]),
    .b_i(b_r[10239:10112]),
    .s_i({ s_r_79__127_, s_r_79__126_, s_r_79__125_, s_r_79__124_, s_r_79__123_, s_r_79__122_, s_r_79__121_, s_r_79__120_, s_r_79__119_, s_r_79__118_, s_r_79__117_, s_r_79__116_, s_r_79__115_, s_r_79__114_, s_r_79__113_, s_r_79__112_, s_r_79__111_, s_r_79__110_, s_r_79__109_, s_r_79__108_, s_r_79__107_, s_r_79__106_, s_r_79__105_, s_r_79__104_, s_r_79__103_, s_r_79__102_, s_r_79__101_, s_r_79__100_, s_r_79__99_, s_r_79__98_, s_r_79__97_, s_r_79__96_, s_r_79__95_, s_r_79__94_, s_r_79__93_, s_r_79__92_, s_r_79__91_, s_r_79__90_, s_r_79__89_, s_r_79__88_, s_r_79__87_, s_r_79__86_, s_r_79__85_, s_r_79__84_, s_r_79__83_, s_r_79__82_, s_r_79__81_, s_r_79__80_, s_r_79__79_, s_r_79__78_, s_r_79__77_, s_r_79__76_, s_r_79__75_, s_r_79__74_, s_r_79__73_, s_r_79__72_, s_r_79__71_, s_r_79__70_, s_r_79__69_, s_r_79__68_, s_r_79__67_, s_r_79__66_, s_r_79__65_, s_r_79__64_, s_r_79__63_, s_r_79__62_, s_r_79__61_, s_r_79__60_, s_r_79__59_, s_r_79__58_, s_r_79__57_, s_r_79__56_, s_r_79__55_, s_r_79__54_, s_r_79__53_, s_r_79__52_, s_r_79__51_, s_r_79__50_, s_r_79__49_, s_r_79__48_, s_r_79__47_, s_r_79__46_, s_r_79__45_, s_r_79__44_, s_r_79__43_, s_r_79__42_, s_r_79__41_, s_r_79__40_, s_r_79__39_, s_r_79__38_, s_r_79__37_, s_r_79__36_, s_r_79__35_, s_r_79__34_, s_r_79__33_, s_r_79__32_, s_r_79__31_, s_r_79__30_, s_r_79__29_, s_r_79__28_, s_r_79__27_, s_r_79__26_, s_r_79__25_, s_r_79__24_, s_r_79__23_, s_r_79__22_, s_r_79__21_, s_r_79__20_, s_r_79__19_, s_r_79__18_, s_r_79__17_, s_r_79__16_, s_r_79__15_, s_r_79__14_, s_r_79__13_, s_r_79__12_, s_r_79__11_, s_r_79__10_, s_r_79__9_, s_r_79__8_, s_r_79__7_, s_r_79__6_, s_r_79__5_, s_r_79__4_, s_r_79__3_, s_r_79__2_, s_r_79__1_, s_r_79__0_ }),
    .c_i(c_r[79]),
    .prod_accum_i({ prod_accum_79__80_, prod_accum_79__79_, prod_accum_79__78_, prod_accum_79__77_, prod_accum_79__76_, prod_accum_79__75_, prod_accum_79__74_, prod_accum_79__73_, prod_accum_79__72_, prod_accum_79__71_, prod_accum_79__70_, prod_accum_79__69_, prod_accum_79__68_, prod_accum_79__67_, prod_accum_79__66_, prod_accum_79__65_, prod_accum_79__64_, prod_accum_79__63_, prod_accum_79__62_, prod_accum_79__61_, prod_accum_79__60_, prod_accum_79__59_, prod_accum_79__58_, prod_accum_79__57_, prod_accum_79__56_, prod_accum_79__55_, prod_accum_79__54_, prod_accum_79__53_, prod_accum_79__52_, prod_accum_79__51_, prod_accum_79__50_, prod_accum_79__49_, prod_accum_79__48_, prod_accum_79__47_, prod_accum_79__46_, prod_accum_79__45_, prod_accum_79__44_, prod_accum_79__43_, prod_accum_79__42_, prod_accum_79__41_, prod_accum_79__40_, prod_accum_79__39_, prod_accum_79__38_, prod_accum_79__37_, prod_accum_79__36_, prod_accum_79__35_, prod_accum_79__34_, prod_accum_79__33_, prod_accum_79__32_, prod_accum_79__31_, prod_accum_79__30_, prod_accum_79__29_, prod_accum_79__28_, prod_accum_79__27_, prod_accum_79__26_, prod_accum_79__25_, prod_accum_79__24_, prod_accum_79__23_, prod_accum_79__22_, prod_accum_79__21_, prod_accum_79__20_, prod_accum_79__19_, prod_accum_79__18_, prod_accum_79__17_, prod_accum_79__16_, prod_accum_79__15_, prod_accum_79__14_, prod_accum_79__13_, prod_accum_79__12_, prod_accum_79__11_, prod_accum_79__10_, prod_accum_79__9_, prod_accum_79__8_, prod_accum_79__7_, prod_accum_79__6_, prod_accum_79__5_, prod_accum_79__4_, prod_accum_79__3_, prod_accum_79__2_, prod_accum_79__1_, prod_accum_79__0_ }),
    .a_o(a_r[10367:10240]),
    .b_o(b_r[10367:10240]),
    .s_o({ s_r_80__127_, s_r_80__126_, s_r_80__125_, s_r_80__124_, s_r_80__123_, s_r_80__122_, s_r_80__121_, s_r_80__120_, s_r_80__119_, s_r_80__118_, s_r_80__117_, s_r_80__116_, s_r_80__115_, s_r_80__114_, s_r_80__113_, s_r_80__112_, s_r_80__111_, s_r_80__110_, s_r_80__109_, s_r_80__108_, s_r_80__107_, s_r_80__106_, s_r_80__105_, s_r_80__104_, s_r_80__103_, s_r_80__102_, s_r_80__101_, s_r_80__100_, s_r_80__99_, s_r_80__98_, s_r_80__97_, s_r_80__96_, s_r_80__95_, s_r_80__94_, s_r_80__93_, s_r_80__92_, s_r_80__91_, s_r_80__90_, s_r_80__89_, s_r_80__88_, s_r_80__87_, s_r_80__86_, s_r_80__85_, s_r_80__84_, s_r_80__83_, s_r_80__82_, s_r_80__81_, s_r_80__80_, s_r_80__79_, s_r_80__78_, s_r_80__77_, s_r_80__76_, s_r_80__75_, s_r_80__74_, s_r_80__73_, s_r_80__72_, s_r_80__71_, s_r_80__70_, s_r_80__69_, s_r_80__68_, s_r_80__67_, s_r_80__66_, s_r_80__65_, s_r_80__64_, s_r_80__63_, s_r_80__62_, s_r_80__61_, s_r_80__60_, s_r_80__59_, s_r_80__58_, s_r_80__57_, s_r_80__56_, s_r_80__55_, s_r_80__54_, s_r_80__53_, s_r_80__52_, s_r_80__51_, s_r_80__50_, s_r_80__49_, s_r_80__48_, s_r_80__47_, s_r_80__46_, s_r_80__45_, s_r_80__44_, s_r_80__43_, s_r_80__42_, s_r_80__41_, s_r_80__40_, s_r_80__39_, s_r_80__38_, s_r_80__37_, s_r_80__36_, s_r_80__35_, s_r_80__34_, s_r_80__33_, s_r_80__32_, s_r_80__31_, s_r_80__30_, s_r_80__29_, s_r_80__28_, s_r_80__27_, s_r_80__26_, s_r_80__25_, s_r_80__24_, s_r_80__23_, s_r_80__22_, s_r_80__21_, s_r_80__20_, s_r_80__19_, s_r_80__18_, s_r_80__17_, s_r_80__16_, s_r_80__15_, s_r_80__14_, s_r_80__13_, s_r_80__12_, s_r_80__11_, s_r_80__10_, s_r_80__9_, s_r_80__8_, s_r_80__7_, s_r_80__6_, s_r_80__5_, s_r_80__4_, s_r_80__3_, s_r_80__2_, s_r_80__1_, s_r_80__0_ }),
    .c_o(c_r[80]),
    .prod_accum_o({ prod_accum_80__81_, prod_accum_80__80_, prod_accum_80__79_, prod_accum_80__78_, prod_accum_80__77_, prod_accum_80__76_, prod_accum_80__75_, prod_accum_80__74_, prod_accum_80__73_, prod_accum_80__72_, prod_accum_80__71_, prod_accum_80__70_, prod_accum_80__69_, prod_accum_80__68_, prod_accum_80__67_, prod_accum_80__66_, prod_accum_80__65_, prod_accum_80__64_, prod_accum_80__63_, prod_accum_80__62_, prod_accum_80__61_, prod_accum_80__60_, prod_accum_80__59_, prod_accum_80__58_, prod_accum_80__57_, prod_accum_80__56_, prod_accum_80__55_, prod_accum_80__54_, prod_accum_80__53_, prod_accum_80__52_, prod_accum_80__51_, prod_accum_80__50_, prod_accum_80__49_, prod_accum_80__48_, prod_accum_80__47_, prod_accum_80__46_, prod_accum_80__45_, prod_accum_80__44_, prod_accum_80__43_, prod_accum_80__42_, prod_accum_80__41_, prod_accum_80__40_, prod_accum_80__39_, prod_accum_80__38_, prod_accum_80__37_, prod_accum_80__36_, prod_accum_80__35_, prod_accum_80__34_, prod_accum_80__33_, prod_accum_80__32_, prod_accum_80__31_, prod_accum_80__30_, prod_accum_80__29_, prod_accum_80__28_, prod_accum_80__27_, prod_accum_80__26_, prod_accum_80__25_, prod_accum_80__24_, prod_accum_80__23_, prod_accum_80__22_, prod_accum_80__21_, prod_accum_80__20_, prod_accum_80__19_, prod_accum_80__18_, prod_accum_80__17_, prod_accum_80__16_, prod_accum_80__15_, prod_accum_80__14_, prod_accum_80__13_, prod_accum_80__12_, prod_accum_80__11_, prod_accum_80__10_, prod_accum_80__9_, prod_accum_80__8_, prod_accum_80__7_, prod_accum_80__6_, prod_accum_80__5_, prod_accum_80__4_, prod_accum_80__3_, prod_accum_80__2_, prod_accum_80__1_, prod_accum_80__0_ })
  );


  bsg_mul_array_row_128_81_x
  genblk1_81__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[10367:10240]),
    .b_i(b_r[10367:10240]),
    .s_i({ s_r_80__127_, s_r_80__126_, s_r_80__125_, s_r_80__124_, s_r_80__123_, s_r_80__122_, s_r_80__121_, s_r_80__120_, s_r_80__119_, s_r_80__118_, s_r_80__117_, s_r_80__116_, s_r_80__115_, s_r_80__114_, s_r_80__113_, s_r_80__112_, s_r_80__111_, s_r_80__110_, s_r_80__109_, s_r_80__108_, s_r_80__107_, s_r_80__106_, s_r_80__105_, s_r_80__104_, s_r_80__103_, s_r_80__102_, s_r_80__101_, s_r_80__100_, s_r_80__99_, s_r_80__98_, s_r_80__97_, s_r_80__96_, s_r_80__95_, s_r_80__94_, s_r_80__93_, s_r_80__92_, s_r_80__91_, s_r_80__90_, s_r_80__89_, s_r_80__88_, s_r_80__87_, s_r_80__86_, s_r_80__85_, s_r_80__84_, s_r_80__83_, s_r_80__82_, s_r_80__81_, s_r_80__80_, s_r_80__79_, s_r_80__78_, s_r_80__77_, s_r_80__76_, s_r_80__75_, s_r_80__74_, s_r_80__73_, s_r_80__72_, s_r_80__71_, s_r_80__70_, s_r_80__69_, s_r_80__68_, s_r_80__67_, s_r_80__66_, s_r_80__65_, s_r_80__64_, s_r_80__63_, s_r_80__62_, s_r_80__61_, s_r_80__60_, s_r_80__59_, s_r_80__58_, s_r_80__57_, s_r_80__56_, s_r_80__55_, s_r_80__54_, s_r_80__53_, s_r_80__52_, s_r_80__51_, s_r_80__50_, s_r_80__49_, s_r_80__48_, s_r_80__47_, s_r_80__46_, s_r_80__45_, s_r_80__44_, s_r_80__43_, s_r_80__42_, s_r_80__41_, s_r_80__40_, s_r_80__39_, s_r_80__38_, s_r_80__37_, s_r_80__36_, s_r_80__35_, s_r_80__34_, s_r_80__33_, s_r_80__32_, s_r_80__31_, s_r_80__30_, s_r_80__29_, s_r_80__28_, s_r_80__27_, s_r_80__26_, s_r_80__25_, s_r_80__24_, s_r_80__23_, s_r_80__22_, s_r_80__21_, s_r_80__20_, s_r_80__19_, s_r_80__18_, s_r_80__17_, s_r_80__16_, s_r_80__15_, s_r_80__14_, s_r_80__13_, s_r_80__12_, s_r_80__11_, s_r_80__10_, s_r_80__9_, s_r_80__8_, s_r_80__7_, s_r_80__6_, s_r_80__5_, s_r_80__4_, s_r_80__3_, s_r_80__2_, s_r_80__1_, s_r_80__0_ }),
    .c_i(c_r[80]),
    .prod_accum_i({ prod_accum_80__81_, prod_accum_80__80_, prod_accum_80__79_, prod_accum_80__78_, prod_accum_80__77_, prod_accum_80__76_, prod_accum_80__75_, prod_accum_80__74_, prod_accum_80__73_, prod_accum_80__72_, prod_accum_80__71_, prod_accum_80__70_, prod_accum_80__69_, prod_accum_80__68_, prod_accum_80__67_, prod_accum_80__66_, prod_accum_80__65_, prod_accum_80__64_, prod_accum_80__63_, prod_accum_80__62_, prod_accum_80__61_, prod_accum_80__60_, prod_accum_80__59_, prod_accum_80__58_, prod_accum_80__57_, prod_accum_80__56_, prod_accum_80__55_, prod_accum_80__54_, prod_accum_80__53_, prod_accum_80__52_, prod_accum_80__51_, prod_accum_80__50_, prod_accum_80__49_, prod_accum_80__48_, prod_accum_80__47_, prod_accum_80__46_, prod_accum_80__45_, prod_accum_80__44_, prod_accum_80__43_, prod_accum_80__42_, prod_accum_80__41_, prod_accum_80__40_, prod_accum_80__39_, prod_accum_80__38_, prod_accum_80__37_, prod_accum_80__36_, prod_accum_80__35_, prod_accum_80__34_, prod_accum_80__33_, prod_accum_80__32_, prod_accum_80__31_, prod_accum_80__30_, prod_accum_80__29_, prod_accum_80__28_, prod_accum_80__27_, prod_accum_80__26_, prod_accum_80__25_, prod_accum_80__24_, prod_accum_80__23_, prod_accum_80__22_, prod_accum_80__21_, prod_accum_80__20_, prod_accum_80__19_, prod_accum_80__18_, prod_accum_80__17_, prod_accum_80__16_, prod_accum_80__15_, prod_accum_80__14_, prod_accum_80__13_, prod_accum_80__12_, prod_accum_80__11_, prod_accum_80__10_, prod_accum_80__9_, prod_accum_80__8_, prod_accum_80__7_, prod_accum_80__6_, prod_accum_80__5_, prod_accum_80__4_, prod_accum_80__3_, prod_accum_80__2_, prod_accum_80__1_, prod_accum_80__0_ }),
    .a_o(a_r[10495:10368]),
    .b_o(b_r[10495:10368]),
    .s_o({ s_r_81__127_, s_r_81__126_, s_r_81__125_, s_r_81__124_, s_r_81__123_, s_r_81__122_, s_r_81__121_, s_r_81__120_, s_r_81__119_, s_r_81__118_, s_r_81__117_, s_r_81__116_, s_r_81__115_, s_r_81__114_, s_r_81__113_, s_r_81__112_, s_r_81__111_, s_r_81__110_, s_r_81__109_, s_r_81__108_, s_r_81__107_, s_r_81__106_, s_r_81__105_, s_r_81__104_, s_r_81__103_, s_r_81__102_, s_r_81__101_, s_r_81__100_, s_r_81__99_, s_r_81__98_, s_r_81__97_, s_r_81__96_, s_r_81__95_, s_r_81__94_, s_r_81__93_, s_r_81__92_, s_r_81__91_, s_r_81__90_, s_r_81__89_, s_r_81__88_, s_r_81__87_, s_r_81__86_, s_r_81__85_, s_r_81__84_, s_r_81__83_, s_r_81__82_, s_r_81__81_, s_r_81__80_, s_r_81__79_, s_r_81__78_, s_r_81__77_, s_r_81__76_, s_r_81__75_, s_r_81__74_, s_r_81__73_, s_r_81__72_, s_r_81__71_, s_r_81__70_, s_r_81__69_, s_r_81__68_, s_r_81__67_, s_r_81__66_, s_r_81__65_, s_r_81__64_, s_r_81__63_, s_r_81__62_, s_r_81__61_, s_r_81__60_, s_r_81__59_, s_r_81__58_, s_r_81__57_, s_r_81__56_, s_r_81__55_, s_r_81__54_, s_r_81__53_, s_r_81__52_, s_r_81__51_, s_r_81__50_, s_r_81__49_, s_r_81__48_, s_r_81__47_, s_r_81__46_, s_r_81__45_, s_r_81__44_, s_r_81__43_, s_r_81__42_, s_r_81__41_, s_r_81__40_, s_r_81__39_, s_r_81__38_, s_r_81__37_, s_r_81__36_, s_r_81__35_, s_r_81__34_, s_r_81__33_, s_r_81__32_, s_r_81__31_, s_r_81__30_, s_r_81__29_, s_r_81__28_, s_r_81__27_, s_r_81__26_, s_r_81__25_, s_r_81__24_, s_r_81__23_, s_r_81__22_, s_r_81__21_, s_r_81__20_, s_r_81__19_, s_r_81__18_, s_r_81__17_, s_r_81__16_, s_r_81__15_, s_r_81__14_, s_r_81__13_, s_r_81__12_, s_r_81__11_, s_r_81__10_, s_r_81__9_, s_r_81__8_, s_r_81__7_, s_r_81__6_, s_r_81__5_, s_r_81__4_, s_r_81__3_, s_r_81__2_, s_r_81__1_, s_r_81__0_ }),
    .c_o(c_r[81]),
    .prod_accum_o({ prod_accum_81__82_, prod_accum_81__81_, prod_accum_81__80_, prod_accum_81__79_, prod_accum_81__78_, prod_accum_81__77_, prod_accum_81__76_, prod_accum_81__75_, prod_accum_81__74_, prod_accum_81__73_, prod_accum_81__72_, prod_accum_81__71_, prod_accum_81__70_, prod_accum_81__69_, prod_accum_81__68_, prod_accum_81__67_, prod_accum_81__66_, prod_accum_81__65_, prod_accum_81__64_, prod_accum_81__63_, prod_accum_81__62_, prod_accum_81__61_, prod_accum_81__60_, prod_accum_81__59_, prod_accum_81__58_, prod_accum_81__57_, prod_accum_81__56_, prod_accum_81__55_, prod_accum_81__54_, prod_accum_81__53_, prod_accum_81__52_, prod_accum_81__51_, prod_accum_81__50_, prod_accum_81__49_, prod_accum_81__48_, prod_accum_81__47_, prod_accum_81__46_, prod_accum_81__45_, prod_accum_81__44_, prod_accum_81__43_, prod_accum_81__42_, prod_accum_81__41_, prod_accum_81__40_, prod_accum_81__39_, prod_accum_81__38_, prod_accum_81__37_, prod_accum_81__36_, prod_accum_81__35_, prod_accum_81__34_, prod_accum_81__33_, prod_accum_81__32_, prod_accum_81__31_, prod_accum_81__30_, prod_accum_81__29_, prod_accum_81__28_, prod_accum_81__27_, prod_accum_81__26_, prod_accum_81__25_, prod_accum_81__24_, prod_accum_81__23_, prod_accum_81__22_, prod_accum_81__21_, prod_accum_81__20_, prod_accum_81__19_, prod_accum_81__18_, prod_accum_81__17_, prod_accum_81__16_, prod_accum_81__15_, prod_accum_81__14_, prod_accum_81__13_, prod_accum_81__12_, prod_accum_81__11_, prod_accum_81__10_, prod_accum_81__9_, prod_accum_81__8_, prod_accum_81__7_, prod_accum_81__6_, prod_accum_81__5_, prod_accum_81__4_, prod_accum_81__3_, prod_accum_81__2_, prod_accum_81__1_, prod_accum_81__0_ })
  );


  bsg_mul_array_row_128_82_x
  genblk1_82__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[10495:10368]),
    .b_i(b_r[10495:10368]),
    .s_i({ s_r_81__127_, s_r_81__126_, s_r_81__125_, s_r_81__124_, s_r_81__123_, s_r_81__122_, s_r_81__121_, s_r_81__120_, s_r_81__119_, s_r_81__118_, s_r_81__117_, s_r_81__116_, s_r_81__115_, s_r_81__114_, s_r_81__113_, s_r_81__112_, s_r_81__111_, s_r_81__110_, s_r_81__109_, s_r_81__108_, s_r_81__107_, s_r_81__106_, s_r_81__105_, s_r_81__104_, s_r_81__103_, s_r_81__102_, s_r_81__101_, s_r_81__100_, s_r_81__99_, s_r_81__98_, s_r_81__97_, s_r_81__96_, s_r_81__95_, s_r_81__94_, s_r_81__93_, s_r_81__92_, s_r_81__91_, s_r_81__90_, s_r_81__89_, s_r_81__88_, s_r_81__87_, s_r_81__86_, s_r_81__85_, s_r_81__84_, s_r_81__83_, s_r_81__82_, s_r_81__81_, s_r_81__80_, s_r_81__79_, s_r_81__78_, s_r_81__77_, s_r_81__76_, s_r_81__75_, s_r_81__74_, s_r_81__73_, s_r_81__72_, s_r_81__71_, s_r_81__70_, s_r_81__69_, s_r_81__68_, s_r_81__67_, s_r_81__66_, s_r_81__65_, s_r_81__64_, s_r_81__63_, s_r_81__62_, s_r_81__61_, s_r_81__60_, s_r_81__59_, s_r_81__58_, s_r_81__57_, s_r_81__56_, s_r_81__55_, s_r_81__54_, s_r_81__53_, s_r_81__52_, s_r_81__51_, s_r_81__50_, s_r_81__49_, s_r_81__48_, s_r_81__47_, s_r_81__46_, s_r_81__45_, s_r_81__44_, s_r_81__43_, s_r_81__42_, s_r_81__41_, s_r_81__40_, s_r_81__39_, s_r_81__38_, s_r_81__37_, s_r_81__36_, s_r_81__35_, s_r_81__34_, s_r_81__33_, s_r_81__32_, s_r_81__31_, s_r_81__30_, s_r_81__29_, s_r_81__28_, s_r_81__27_, s_r_81__26_, s_r_81__25_, s_r_81__24_, s_r_81__23_, s_r_81__22_, s_r_81__21_, s_r_81__20_, s_r_81__19_, s_r_81__18_, s_r_81__17_, s_r_81__16_, s_r_81__15_, s_r_81__14_, s_r_81__13_, s_r_81__12_, s_r_81__11_, s_r_81__10_, s_r_81__9_, s_r_81__8_, s_r_81__7_, s_r_81__6_, s_r_81__5_, s_r_81__4_, s_r_81__3_, s_r_81__2_, s_r_81__1_, s_r_81__0_ }),
    .c_i(c_r[81]),
    .prod_accum_i({ prod_accum_81__82_, prod_accum_81__81_, prod_accum_81__80_, prod_accum_81__79_, prod_accum_81__78_, prod_accum_81__77_, prod_accum_81__76_, prod_accum_81__75_, prod_accum_81__74_, prod_accum_81__73_, prod_accum_81__72_, prod_accum_81__71_, prod_accum_81__70_, prod_accum_81__69_, prod_accum_81__68_, prod_accum_81__67_, prod_accum_81__66_, prod_accum_81__65_, prod_accum_81__64_, prod_accum_81__63_, prod_accum_81__62_, prod_accum_81__61_, prod_accum_81__60_, prod_accum_81__59_, prod_accum_81__58_, prod_accum_81__57_, prod_accum_81__56_, prod_accum_81__55_, prod_accum_81__54_, prod_accum_81__53_, prod_accum_81__52_, prod_accum_81__51_, prod_accum_81__50_, prod_accum_81__49_, prod_accum_81__48_, prod_accum_81__47_, prod_accum_81__46_, prod_accum_81__45_, prod_accum_81__44_, prod_accum_81__43_, prod_accum_81__42_, prod_accum_81__41_, prod_accum_81__40_, prod_accum_81__39_, prod_accum_81__38_, prod_accum_81__37_, prod_accum_81__36_, prod_accum_81__35_, prod_accum_81__34_, prod_accum_81__33_, prod_accum_81__32_, prod_accum_81__31_, prod_accum_81__30_, prod_accum_81__29_, prod_accum_81__28_, prod_accum_81__27_, prod_accum_81__26_, prod_accum_81__25_, prod_accum_81__24_, prod_accum_81__23_, prod_accum_81__22_, prod_accum_81__21_, prod_accum_81__20_, prod_accum_81__19_, prod_accum_81__18_, prod_accum_81__17_, prod_accum_81__16_, prod_accum_81__15_, prod_accum_81__14_, prod_accum_81__13_, prod_accum_81__12_, prod_accum_81__11_, prod_accum_81__10_, prod_accum_81__9_, prod_accum_81__8_, prod_accum_81__7_, prod_accum_81__6_, prod_accum_81__5_, prod_accum_81__4_, prod_accum_81__3_, prod_accum_81__2_, prod_accum_81__1_, prod_accum_81__0_ }),
    .a_o(a_r[10623:10496]),
    .b_o(b_r[10623:10496]),
    .s_o({ s_r_82__127_, s_r_82__126_, s_r_82__125_, s_r_82__124_, s_r_82__123_, s_r_82__122_, s_r_82__121_, s_r_82__120_, s_r_82__119_, s_r_82__118_, s_r_82__117_, s_r_82__116_, s_r_82__115_, s_r_82__114_, s_r_82__113_, s_r_82__112_, s_r_82__111_, s_r_82__110_, s_r_82__109_, s_r_82__108_, s_r_82__107_, s_r_82__106_, s_r_82__105_, s_r_82__104_, s_r_82__103_, s_r_82__102_, s_r_82__101_, s_r_82__100_, s_r_82__99_, s_r_82__98_, s_r_82__97_, s_r_82__96_, s_r_82__95_, s_r_82__94_, s_r_82__93_, s_r_82__92_, s_r_82__91_, s_r_82__90_, s_r_82__89_, s_r_82__88_, s_r_82__87_, s_r_82__86_, s_r_82__85_, s_r_82__84_, s_r_82__83_, s_r_82__82_, s_r_82__81_, s_r_82__80_, s_r_82__79_, s_r_82__78_, s_r_82__77_, s_r_82__76_, s_r_82__75_, s_r_82__74_, s_r_82__73_, s_r_82__72_, s_r_82__71_, s_r_82__70_, s_r_82__69_, s_r_82__68_, s_r_82__67_, s_r_82__66_, s_r_82__65_, s_r_82__64_, s_r_82__63_, s_r_82__62_, s_r_82__61_, s_r_82__60_, s_r_82__59_, s_r_82__58_, s_r_82__57_, s_r_82__56_, s_r_82__55_, s_r_82__54_, s_r_82__53_, s_r_82__52_, s_r_82__51_, s_r_82__50_, s_r_82__49_, s_r_82__48_, s_r_82__47_, s_r_82__46_, s_r_82__45_, s_r_82__44_, s_r_82__43_, s_r_82__42_, s_r_82__41_, s_r_82__40_, s_r_82__39_, s_r_82__38_, s_r_82__37_, s_r_82__36_, s_r_82__35_, s_r_82__34_, s_r_82__33_, s_r_82__32_, s_r_82__31_, s_r_82__30_, s_r_82__29_, s_r_82__28_, s_r_82__27_, s_r_82__26_, s_r_82__25_, s_r_82__24_, s_r_82__23_, s_r_82__22_, s_r_82__21_, s_r_82__20_, s_r_82__19_, s_r_82__18_, s_r_82__17_, s_r_82__16_, s_r_82__15_, s_r_82__14_, s_r_82__13_, s_r_82__12_, s_r_82__11_, s_r_82__10_, s_r_82__9_, s_r_82__8_, s_r_82__7_, s_r_82__6_, s_r_82__5_, s_r_82__4_, s_r_82__3_, s_r_82__2_, s_r_82__1_, s_r_82__0_ }),
    .c_o(c_r[82]),
    .prod_accum_o({ prod_accum_82__83_, prod_accum_82__82_, prod_accum_82__81_, prod_accum_82__80_, prod_accum_82__79_, prod_accum_82__78_, prod_accum_82__77_, prod_accum_82__76_, prod_accum_82__75_, prod_accum_82__74_, prod_accum_82__73_, prod_accum_82__72_, prod_accum_82__71_, prod_accum_82__70_, prod_accum_82__69_, prod_accum_82__68_, prod_accum_82__67_, prod_accum_82__66_, prod_accum_82__65_, prod_accum_82__64_, prod_accum_82__63_, prod_accum_82__62_, prod_accum_82__61_, prod_accum_82__60_, prod_accum_82__59_, prod_accum_82__58_, prod_accum_82__57_, prod_accum_82__56_, prod_accum_82__55_, prod_accum_82__54_, prod_accum_82__53_, prod_accum_82__52_, prod_accum_82__51_, prod_accum_82__50_, prod_accum_82__49_, prod_accum_82__48_, prod_accum_82__47_, prod_accum_82__46_, prod_accum_82__45_, prod_accum_82__44_, prod_accum_82__43_, prod_accum_82__42_, prod_accum_82__41_, prod_accum_82__40_, prod_accum_82__39_, prod_accum_82__38_, prod_accum_82__37_, prod_accum_82__36_, prod_accum_82__35_, prod_accum_82__34_, prod_accum_82__33_, prod_accum_82__32_, prod_accum_82__31_, prod_accum_82__30_, prod_accum_82__29_, prod_accum_82__28_, prod_accum_82__27_, prod_accum_82__26_, prod_accum_82__25_, prod_accum_82__24_, prod_accum_82__23_, prod_accum_82__22_, prod_accum_82__21_, prod_accum_82__20_, prod_accum_82__19_, prod_accum_82__18_, prod_accum_82__17_, prod_accum_82__16_, prod_accum_82__15_, prod_accum_82__14_, prod_accum_82__13_, prod_accum_82__12_, prod_accum_82__11_, prod_accum_82__10_, prod_accum_82__9_, prod_accum_82__8_, prod_accum_82__7_, prod_accum_82__6_, prod_accum_82__5_, prod_accum_82__4_, prod_accum_82__3_, prod_accum_82__2_, prod_accum_82__1_, prod_accum_82__0_ })
  );


  bsg_mul_array_row_128_83_x
  genblk1_83__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[10623:10496]),
    .b_i(b_r[10623:10496]),
    .s_i({ s_r_82__127_, s_r_82__126_, s_r_82__125_, s_r_82__124_, s_r_82__123_, s_r_82__122_, s_r_82__121_, s_r_82__120_, s_r_82__119_, s_r_82__118_, s_r_82__117_, s_r_82__116_, s_r_82__115_, s_r_82__114_, s_r_82__113_, s_r_82__112_, s_r_82__111_, s_r_82__110_, s_r_82__109_, s_r_82__108_, s_r_82__107_, s_r_82__106_, s_r_82__105_, s_r_82__104_, s_r_82__103_, s_r_82__102_, s_r_82__101_, s_r_82__100_, s_r_82__99_, s_r_82__98_, s_r_82__97_, s_r_82__96_, s_r_82__95_, s_r_82__94_, s_r_82__93_, s_r_82__92_, s_r_82__91_, s_r_82__90_, s_r_82__89_, s_r_82__88_, s_r_82__87_, s_r_82__86_, s_r_82__85_, s_r_82__84_, s_r_82__83_, s_r_82__82_, s_r_82__81_, s_r_82__80_, s_r_82__79_, s_r_82__78_, s_r_82__77_, s_r_82__76_, s_r_82__75_, s_r_82__74_, s_r_82__73_, s_r_82__72_, s_r_82__71_, s_r_82__70_, s_r_82__69_, s_r_82__68_, s_r_82__67_, s_r_82__66_, s_r_82__65_, s_r_82__64_, s_r_82__63_, s_r_82__62_, s_r_82__61_, s_r_82__60_, s_r_82__59_, s_r_82__58_, s_r_82__57_, s_r_82__56_, s_r_82__55_, s_r_82__54_, s_r_82__53_, s_r_82__52_, s_r_82__51_, s_r_82__50_, s_r_82__49_, s_r_82__48_, s_r_82__47_, s_r_82__46_, s_r_82__45_, s_r_82__44_, s_r_82__43_, s_r_82__42_, s_r_82__41_, s_r_82__40_, s_r_82__39_, s_r_82__38_, s_r_82__37_, s_r_82__36_, s_r_82__35_, s_r_82__34_, s_r_82__33_, s_r_82__32_, s_r_82__31_, s_r_82__30_, s_r_82__29_, s_r_82__28_, s_r_82__27_, s_r_82__26_, s_r_82__25_, s_r_82__24_, s_r_82__23_, s_r_82__22_, s_r_82__21_, s_r_82__20_, s_r_82__19_, s_r_82__18_, s_r_82__17_, s_r_82__16_, s_r_82__15_, s_r_82__14_, s_r_82__13_, s_r_82__12_, s_r_82__11_, s_r_82__10_, s_r_82__9_, s_r_82__8_, s_r_82__7_, s_r_82__6_, s_r_82__5_, s_r_82__4_, s_r_82__3_, s_r_82__2_, s_r_82__1_, s_r_82__0_ }),
    .c_i(c_r[82]),
    .prod_accum_i({ prod_accum_82__83_, prod_accum_82__82_, prod_accum_82__81_, prod_accum_82__80_, prod_accum_82__79_, prod_accum_82__78_, prod_accum_82__77_, prod_accum_82__76_, prod_accum_82__75_, prod_accum_82__74_, prod_accum_82__73_, prod_accum_82__72_, prod_accum_82__71_, prod_accum_82__70_, prod_accum_82__69_, prod_accum_82__68_, prod_accum_82__67_, prod_accum_82__66_, prod_accum_82__65_, prod_accum_82__64_, prod_accum_82__63_, prod_accum_82__62_, prod_accum_82__61_, prod_accum_82__60_, prod_accum_82__59_, prod_accum_82__58_, prod_accum_82__57_, prod_accum_82__56_, prod_accum_82__55_, prod_accum_82__54_, prod_accum_82__53_, prod_accum_82__52_, prod_accum_82__51_, prod_accum_82__50_, prod_accum_82__49_, prod_accum_82__48_, prod_accum_82__47_, prod_accum_82__46_, prod_accum_82__45_, prod_accum_82__44_, prod_accum_82__43_, prod_accum_82__42_, prod_accum_82__41_, prod_accum_82__40_, prod_accum_82__39_, prod_accum_82__38_, prod_accum_82__37_, prod_accum_82__36_, prod_accum_82__35_, prod_accum_82__34_, prod_accum_82__33_, prod_accum_82__32_, prod_accum_82__31_, prod_accum_82__30_, prod_accum_82__29_, prod_accum_82__28_, prod_accum_82__27_, prod_accum_82__26_, prod_accum_82__25_, prod_accum_82__24_, prod_accum_82__23_, prod_accum_82__22_, prod_accum_82__21_, prod_accum_82__20_, prod_accum_82__19_, prod_accum_82__18_, prod_accum_82__17_, prod_accum_82__16_, prod_accum_82__15_, prod_accum_82__14_, prod_accum_82__13_, prod_accum_82__12_, prod_accum_82__11_, prod_accum_82__10_, prod_accum_82__9_, prod_accum_82__8_, prod_accum_82__7_, prod_accum_82__6_, prod_accum_82__5_, prod_accum_82__4_, prod_accum_82__3_, prod_accum_82__2_, prod_accum_82__1_, prod_accum_82__0_ }),
    .a_o(a_r[10751:10624]),
    .b_o(b_r[10751:10624]),
    .s_o({ s_r_83__127_, s_r_83__126_, s_r_83__125_, s_r_83__124_, s_r_83__123_, s_r_83__122_, s_r_83__121_, s_r_83__120_, s_r_83__119_, s_r_83__118_, s_r_83__117_, s_r_83__116_, s_r_83__115_, s_r_83__114_, s_r_83__113_, s_r_83__112_, s_r_83__111_, s_r_83__110_, s_r_83__109_, s_r_83__108_, s_r_83__107_, s_r_83__106_, s_r_83__105_, s_r_83__104_, s_r_83__103_, s_r_83__102_, s_r_83__101_, s_r_83__100_, s_r_83__99_, s_r_83__98_, s_r_83__97_, s_r_83__96_, s_r_83__95_, s_r_83__94_, s_r_83__93_, s_r_83__92_, s_r_83__91_, s_r_83__90_, s_r_83__89_, s_r_83__88_, s_r_83__87_, s_r_83__86_, s_r_83__85_, s_r_83__84_, s_r_83__83_, s_r_83__82_, s_r_83__81_, s_r_83__80_, s_r_83__79_, s_r_83__78_, s_r_83__77_, s_r_83__76_, s_r_83__75_, s_r_83__74_, s_r_83__73_, s_r_83__72_, s_r_83__71_, s_r_83__70_, s_r_83__69_, s_r_83__68_, s_r_83__67_, s_r_83__66_, s_r_83__65_, s_r_83__64_, s_r_83__63_, s_r_83__62_, s_r_83__61_, s_r_83__60_, s_r_83__59_, s_r_83__58_, s_r_83__57_, s_r_83__56_, s_r_83__55_, s_r_83__54_, s_r_83__53_, s_r_83__52_, s_r_83__51_, s_r_83__50_, s_r_83__49_, s_r_83__48_, s_r_83__47_, s_r_83__46_, s_r_83__45_, s_r_83__44_, s_r_83__43_, s_r_83__42_, s_r_83__41_, s_r_83__40_, s_r_83__39_, s_r_83__38_, s_r_83__37_, s_r_83__36_, s_r_83__35_, s_r_83__34_, s_r_83__33_, s_r_83__32_, s_r_83__31_, s_r_83__30_, s_r_83__29_, s_r_83__28_, s_r_83__27_, s_r_83__26_, s_r_83__25_, s_r_83__24_, s_r_83__23_, s_r_83__22_, s_r_83__21_, s_r_83__20_, s_r_83__19_, s_r_83__18_, s_r_83__17_, s_r_83__16_, s_r_83__15_, s_r_83__14_, s_r_83__13_, s_r_83__12_, s_r_83__11_, s_r_83__10_, s_r_83__9_, s_r_83__8_, s_r_83__7_, s_r_83__6_, s_r_83__5_, s_r_83__4_, s_r_83__3_, s_r_83__2_, s_r_83__1_, s_r_83__0_ }),
    .c_o(c_r[83]),
    .prod_accum_o({ prod_accum_83__84_, prod_accum_83__83_, prod_accum_83__82_, prod_accum_83__81_, prod_accum_83__80_, prod_accum_83__79_, prod_accum_83__78_, prod_accum_83__77_, prod_accum_83__76_, prod_accum_83__75_, prod_accum_83__74_, prod_accum_83__73_, prod_accum_83__72_, prod_accum_83__71_, prod_accum_83__70_, prod_accum_83__69_, prod_accum_83__68_, prod_accum_83__67_, prod_accum_83__66_, prod_accum_83__65_, prod_accum_83__64_, prod_accum_83__63_, prod_accum_83__62_, prod_accum_83__61_, prod_accum_83__60_, prod_accum_83__59_, prod_accum_83__58_, prod_accum_83__57_, prod_accum_83__56_, prod_accum_83__55_, prod_accum_83__54_, prod_accum_83__53_, prod_accum_83__52_, prod_accum_83__51_, prod_accum_83__50_, prod_accum_83__49_, prod_accum_83__48_, prod_accum_83__47_, prod_accum_83__46_, prod_accum_83__45_, prod_accum_83__44_, prod_accum_83__43_, prod_accum_83__42_, prod_accum_83__41_, prod_accum_83__40_, prod_accum_83__39_, prod_accum_83__38_, prod_accum_83__37_, prod_accum_83__36_, prod_accum_83__35_, prod_accum_83__34_, prod_accum_83__33_, prod_accum_83__32_, prod_accum_83__31_, prod_accum_83__30_, prod_accum_83__29_, prod_accum_83__28_, prod_accum_83__27_, prod_accum_83__26_, prod_accum_83__25_, prod_accum_83__24_, prod_accum_83__23_, prod_accum_83__22_, prod_accum_83__21_, prod_accum_83__20_, prod_accum_83__19_, prod_accum_83__18_, prod_accum_83__17_, prod_accum_83__16_, prod_accum_83__15_, prod_accum_83__14_, prod_accum_83__13_, prod_accum_83__12_, prod_accum_83__11_, prod_accum_83__10_, prod_accum_83__9_, prod_accum_83__8_, prod_accum_83__7_, prod_accum_83__6_, prod_accum_83__5_, prod_accum_83__4_, prod_accum_83__3_, prod_accum_83__2_, prod_accum_83__1_, prod_accum_83__0_ })
  );


  bsg_mul_array_row_128_84_x
  genblk1_84__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[10751:10624]),
    .b_i(b_r[10751:10624]),
    .s_i({ s_r_83__127_, s_r_83__126_, s_r_83__125_, s_r_83__124_, s_r_83__123_, s_r_83__122_, s_r_83__121_, s_r_83__120_, s_r_83__119_, s_r_83__118_, s_r_83__117_, s_r_83__116_, s_r_83__115_, s_r_83__114_, s_r_83__113_, s_r_83__112_, s_r_83__111_, s_r_83__110_, s_r_83__109_, s_r_83__108_, s_r_83__107_, s_r_83__106_, s_r_83__105_, s_r_83__104_, s_r_83__103_, s_r_83__102_, s_r_83__101_, s_r_83__100_, s_r_83__99_, s_r_83__98_, s_r_83__97_, s_r_83__96_, s_r_83__95_, s_r_83__94_, s_r_83__93_, s_r_83__92_, s_r_83__91_, s_r_83__90_, s_r_83__89_, s_r_83__88_, s_r_83__87_, s_r_83__86_, s_r_83__85_, s_r_83__84_, s_r_83__83_, s_r_83__82_, s_r_83__81_, s_r_83__80_, s_r_83__79_, s_r_83__78_, s_r_83__77_, s_r_83__76_, s_r_83__75_, s_r_83__74_, s_r_83__73_, s_r_83__72_, s_r_83__71_, s_r_83__70_, s_r_83__69_, s_r_83__68_, s_r_83__67_, s_r_83__66_, s_r_83__65_, s_r_83__64_, s_r_83__63_, s_r_83__62_, s_r_83__61_, s_r_83__60_, s_r_83__59_, s_r_83__58_, s_r_83__57_, s_r_83__56_, s_r_83__55_, s_r_83__54_, s_r_83__53_, s_r_83__52_, s_r_83__51_, s_r_83__50_, s_r_83__49_, s_r_83__48_, s_r_83__47_, s_r_83__46_, s_r_83__45_, s_r_83__44_, s_r_83__43_, s_r_83__42_, s_r_83__41_, s_r_83__40_, s_r_83__39_, s_r_83__38_, s_r_83__37_, s_r_83__36_, s_r_83__35_, s_r_83__34_, s_r_83__33_, s_r_83__32_, s_r_83__31_, s_r_83__30_, s_r_83__29_, s_r_83__28_, s_r_83__27_, s_r_83__26_, s_r_83__25_, s_r_83__24_, s_r_83__23_, s_r_83__22_, s_r_83__21_, s_r_83__20_, s_r_83__19_, s_r_83__18_, s_r_83__17_, s_r_83__16_, s_r_83__15_, s_r_83__14_, s_r_83__13_, s_r_83__12_, s_r_83__11_, s_r_83__10_, s_r_83__9_, s_r_83__8_, s_r_83__7_, s_r_83__6_, s_r_83__5_, s_r_83__4_, s_r_83__3_, s_r_83__2_, s_r_83__1_, s_r_83__0_ }),
    .c_i(c_r[83]),
    .prod_accum_i({ prod_accum_83__84_, prod_accum_83__83_, prod_accum_83__82_, prod_accum_83__81_, prod_accum_83__80_, prod_accum_83__79_, prod_accum_83__78_, prod_accum_83__77_, prod_accum_83__76_, prod_accum_83__75_, prod_accum_83__74_, prod_accum_83__73_, prod_accum_83__72_, prod_accum_83__71_, prod_accum_83__70_, prod_accum_83__69_, prod_accum_83__68_, prod_accum_83__67_, prod_accum_83__66_, prod_accum_83__65_, prod_accum_83__64_, prod_accum_83__63_, prod_accum_83__62_, prod_accum_83__61_, prod_accum_83__60_, prod_accum_83__59_, prod_accum_83__58_, prod_accum_83__57_, prod_accum_83__56_, prod_accum_83__55_, prod_accum_83__54_, prod_accum_83__53_, prod_accum_83__52_, prod_accum_83__51_, prod_accum_83__50_, prod_accum_83__49_, prod_accum_83__48_, prod_accum_83__47_, prod_accum_83__46_, prod_accum_83__45_, prod_accum_83__44_, prod_accum_83__43_, prod_accum_83__42_, prod_accum_83__41_, prod_accum_83__40_, prod_accum_83__39_, prod_accum_83__38_, prod_accum_83__37_, prod_accum_83__36_, prod_accum_83__35_, prod_accum_83__34_, prod_accum_83__33_, prod_accum_83__32_, prod_accum_83__31_, prod_accum_83__30_, prod_accum_83__29_, prod_accum_83__28_, prod_accum_83__27_, prod_accum_83__26_, prod_accum_83__25_, prod_accum_83__24_, prod_accum_83__23_, prod_accum_83__22_, prod_accum_83__21_, prod_accum_83__20_, prod_accum_83__19_, prod_accum_83__18_, prod_accum_83__17_, prod_accum_83__16_, prod_accum_83__15_, prod_accum_83__14_, prod_accum_83__13_, prod_accum_83__12_, prod_accum_83__11_, prod_accum_83__10_, prod_accum_83__9_, prod_accum_83__8_, prod_accum_83__7_, prod_accum_83__6_, prod_accum_83__5_, prod_accum_83__4_, prod_accum_83__3_, prod_accum_83__2_, prod_accum_83__1_, prod_accum_83__0_ }),
    .a_o(a_r[10879:10752]),
    .b_o(b_r[10879:10752]),
    .s_o({ s_r_84__127_, s_r_84__126_, s_r_84__125_, s_r_84__124_, s_r_84__123_, s_r_84__122_, s_r_84__121_, s_r_84__120_, s_r_84__119_, s_r_84__118_, s_r_84__117_, s_r_84__116_, s_r_84__115_, s_r_84__114_, s_r_84__113_, s_r_84__112_, s_r_84__111_, s_r_84__110_, s_r_84__109_, s_r_84__108_, s_r_84__107_, s_r_84__106_, s_r_84__105_, s_r_84__104_, s_r_84__103_, s_r_84__102_, s_r_84__101_, s_r_84__100_, s_r_84__99_, s_r_84__98_, s_r_84__97_, s_r_84__96_, s_r_84__95_, s_r_84__94_, s_r_84__93_, s_r_84__92_, s_r_84__91_, s_r_84__90_, s_r_84__89_, s_r_84__88_, s_r_84__87_, s_r_84__86_, s_r_84__85_, s_r_84__84_, s_r_84__83_, s_r_84__82_, s_r_84__81_, s_r_84__80_, s_r_84__79_, s_r_84__78_, s_r_84__77_, s_r_84__76_, s_r_84__75_, s_r_84__74_, s_r_84__73_, s_r_84__72_, s_r_84__71_, s_r_84__70_, s_r_84__69_, s_r_84__68_, s_r_84__67_, s_r_84__66_, s_r_84__65_, s_r_84__64_, s_r_84__63_, s_r_84__62_, s_r_84__61_, s_r_84__60_, s_r_84__59_, s_r_84__58_, s_r_84__57_, s_r_84__56_, s_r_84__55_, s_r_84__54_, s_r_84__53_, s_r_84__52_, s_r_84__51_, s_r_84__50_, s_r_84__49_, s_r_84__48_, s_r_84__47_, s_r_84__46_, s_r_84__45_, s_r_84__44_, s_r_84__43_, s_r_84__42_, s_r_84__41_, s_r_84__40_, s_r_84__39_, s_r_84__38_, s_r_84__37_, s_r_84__36_, s_r_84__35_, s_r_84__34_, s_r_84__33_, s_r_84__32_, s_r_84__31_, s_r_84__30_, s_r_84__29_, s_r_84__28_, s_r_84__27_, s_r_84__26_, s_r_84__25_, s_r_84__24_, s_r_84__23_, s_r_84__22_, s_r_84__21_, s_r_84__20_, s_r_84__19_, s_r_84__18_, s_r_84__17_, s_r_84__16_, s_r_84__15_, s_r_84__14_, s_r_84__13_, s_r_84__12_, s_r_84__11_, s_r_84__10_, s_r_84__9_, s_r_84__8_, s_r_84__7_, s_r_84__6_, s_r_84__5_, s_r_84__4_, s_r_84__3_, s_r_84__2_, s_r_84__1_, s_r_84__0_ }),
    .c_o(c_r[84]),
    .prod_accum_o({ prod_accum_84__85_, prod_accum_84__84_, prod_accum_84__83_, prod_accum_84__82_, prod_accum_84__81_, prod_accum_84__80_, prod_accum_84__79_, prod_accum_84__78_, prod_accum_84__77_, prod_accum_84__76_, prod_accum_84__75_, prod_accum_84__74_, prod_accum_84__73_, prod_accum_84__72_, prod_accum_84__71_, prod_accum_84__70_, prod_accum_84__69_, prod_accum_84__68_, prod_accum_84__67_, prod_accum_84__66_, prod_accum_84__65_, prod_accum_84__64_, prod_accum_84__63_, prod_accum_84__62_, prod_accum_84__61_, prod_accum_84__60_, prod_accum_84__59_, prod_accum_84__58_, prod_accum_84__57_, prod_accum_84__56_, prod_accum_84__55_, prod_accum_84__54_, prod_accum_84__53_, prod_accum_84__52_, prod_accum_84__51_, prod_accum_84__50_, prod_accum_84__49_, prod_accum_84__48_, prod_accum_84__47_, prod_accum_84__46_, prod_accum_84__45_, prod_accum_84__44_, prod_accum_84__43_, prod_accum_84__42_, prod_accum_84__41_, prod_accum_84__40_, prod_accum_84__39_, prod_accum_84__38_, prod_accum_84__37_, prod_accum_84__36_, prod_accum_84__35_, prod_accum_84__34_, prod_accum_84__33_, prod_accum_84__32_, prod_accum_84__31_, prod_accum_84__30_, prod_accum_84__29_, prod_accum_84__28_, prod_accum_84__27_, prod_accum_84__26_, prod_accum_84__25_, prod_accum_84__24_, prod_accum_84__23_, prod_accum_84__22_, prod_accum_84__21_, prod_accum_84__20_, prod_accum_84__19_, prod_accum_84__18_, prod_accum_84__17_, prod_accum_84__16_, prod_accum_84__15_, prod_accum_84__14_, prod_accum_84__13_, prod_accum_84__12_, prod_accum_84__11_, prod_accum_84__10_, prod_accum_84__9_, prod_accum_84__8_, prod_accum_84__7_, prod_accum_84__6_, prod_accum_84__5_, prod_accum_84__4_, prod_accum_84__3_, prod_accum_84__2_, prod_accum_84__1_, prod_accum_84__0_ })
  );


  bsg_mul_array_row_128_85_x
  genblk1_85__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[10879:10752]),
    .b_i(b_r[10879:10752]),
    .s_i({ s_r_84__127_, s_r_84__126_, s_r_84__125_, s_r_84__124_, s_r_84__123_, s_r_84__122_, s_r_84__121_, s_r_84__120_, s_r_84__119_, s_r_84__118_, s_r_84__117_, s_r_84__116_, s_r_84__115_, s_r_84__114_, s_r_84__113_, s_r_84__112_, s_r_84__111_, s_r_84__110_, s_r_84__109_, s_r_84__108_, s_r_84__107_, s_r_84__106_, s_r_84__105_, s_r_84__104_, s_r_84__103_, s_r_84__102_, s_r_84__101_, s_r_84__100_, s_r_84__99_, s_r_84__98_, s_r_84__97_, s_r_84__96_, s_r_84__95_, s_r_84__94_, s_r_84__93_, s_r_84__92_, s_r_84__91_, s_r_84__90_, s_r_84__89_, s_r_84__88_, s_r_84__87_, s_r_84__86_, s_r_84__85_, s_r_84__84_, s_r_84__83_, s_r_84__82_, s_r_84__81_, s_r_84__80_, s_r_84__79_, s_r_84__78_, s_r_84__77_, s_r_84__76_, s_r_84__75_, s_r_84__74_, s_r_84__73_, s_r_84__72_, s_r_84__71_, s_r_84__70_, s_r_84__69_, s_r_84__68_, s_r_84__67_, s_r_84__66_, s_r_84__65_, s_r_84__64_, s_r_84__63_, s_r_84__62_, s_r_84__61_, s_r_84__60_, s_r_84__59_, s_r_84__58_, s_r_84__57_, s_r_84__56_, s_r_84__55_, s_r_84__54_, s_r_84__53_, s_r_84__52_, s_r_84__51_, s_r_84__50_, s_r_84__49_, s_r_84__48_, s_r_84__47_, s_r_84__46_, s_r_84__45_, s_r_84__44_, s_r_84__43_, s_r_84__42_, s_r_84__41_, s_r_84__40_, s_r_84__39_, s_r_84__38_, s_r_84__37_, s_r_84__36_, s_r_84__35_, s_r_84__34_, s_r_84__33_, s_r_84__32_, s_r_84__31_, s_r_84__30_, s_r_84__29_, s_r_84__28_, s_r_84__27_, s_r_84__26_, s_r_84__25_, s_r_84__24_, s_r_84__23_, s_r_84__22_, s_r_84__21_, s_r_84__20_, s_r_84__19_, s_r_84__18_, s_r_84__17_, s_r_84__16_, s_r_84__15_, s_r_84__14_, s_r_84__13_, s_r_84__12_, s_r_84__11_, s_r_84__10_, s_r_84__9_, s_r_84__8_, s_r_84__7_, s_r_84__6_, s_r_84__5_, s_r_84__4_, s_r_84__3_, s_r_84__2_, s_r_84__1_, s_r_84__0_ }),
    .c_i(c_r[84]),
    .prod_accum_i({ prod_accum_84__85_, prod_accum_84__84_, prod_accum_84__83_, prod_accum_84__82_, prod_accum_84__81_, prod_accum_84__80_, prod_accum_84__79_, prod_accum_84__78_, prod_accum_84__77_, prod_accum_84__76_, prod_accum_84__75_, prod_accum_84__74_, prod_accum_84__73_, prod_accum_84__72_, prod_accum_84__71_, prod_accum_84__70_, prod_accum_84__69_, prod_accum_84__68_, prod_accum_84__67_, prod_accum_84__66_, prod_accum_84__65_, prod_accum_84__64_, prod_accum_84__63_, prod_accum_84__62_, prod_accum_84__61_, prod_accum_84__60_, prod_accum_84__59_, prod_accum_84__58_, prod_accum_84__57_, prod_accum_84__56_, prod_accum_84__55_, prod_accum_84__54_, prod_accum_84__53_, prod_accum_84__52_, prod_accum_84__51_, prod_accum_84__50_, prod_accum_84__49_, prod_accum_84__48_, prod_accum_84__47_, prod_accum_84__46_, prod_accum_84__45_, prod_accum_84__44_, prod_accum_84__43_, prod_accum_84__42_, prod_accum_84__41_, prod_accum_84__40_, prod_accum_84__39_, prod_accum_84__38_, prod_accum_84__37_, prod_accum_84__36_, prod_accum_84__35_, prod_accum_84__34_, prod_accum_84__33_, prod_accum_84__32_, prod_accum_84__31_, prod_accum_84__30_, prod_accum_84__29_, prod_accum_84__28_, prod_accum_84__27_, prod_accum_84__26_, prod_accum_84__25_, prod_accum_84__24_, prod_accum_84__23_, prod_accum_84__22_, prod_accum_84__21_, prod_accum_84__20_, prod_accum_84__19_, prod_accum_84__18_, prod_accum_84__17_, prod_accum_84__16_, prod_accum_84__15_, prod_accum_84__14_, prod_accum_84__13_, prod_accum_84__12_, prod_accum_84__11_, prod_accum_84__10_, prod_accum_84__9_, prod_accum_84__8_, prod_accum_84__7_, prod_accum_84__6_, prod_accum_84__5_, prod_accum_84__4_, prod_accum_84__3_, prod_accum_84__2_, prod_accum_84__1_, prod_accum_84__0_ }),
    .a_o(a_r[11007:10880]),
    .b_o(b_r[11007:10880]),
    .s_o({ s_r_85__127_, s_r_85__126_, s_r_85__125_, s_r_85__124_, s_r_85__123_, s_r_85__122_, s_r_85__121_, s_r_85__120_, s_r_85__119_, s_r_85__118_, s_r_85__117_, s_r_85__116_, s_r_85__115_, s_r_85__114_, s_r_85__113_, s_r_85__112_, s_r_85__111_, s_r_85__110_, s_r_85__109_, s_r_85__108_, s_r_85__107_, s_r_85__106_, s_r_85__105_, s_r_85__104_, s_r_85__103_, s_r_85__102_, s_r_85__101_, s_r_85__100_, s_r_85__99_, s_r_85__98_, s_r_85__97_, s_r_85__96_, s_r_85__95_, s_r_85__94_, s_r_85__93_, s_r_85__92_, s_r_85__91_, s_r_85__90_, s_r_85__89_, s_r_85__88_, s_r_85__87_, s_r_85__86_, s_r_85__85_, s_r_85__84_, s_r_85__83_, s_r_85__82_, s_r_85__81_, s_r_85__80_, s_r_85__79_, s_r_85__78_, s_r_85__77_, s_r_85__76_, s_r_85__75_, s_r_85__74_, s_r_85__73_, s_r_85__72_, s_r_85__71_, s_r_85__70_, s_r_85__69_, s_r_85__68_, s_r_85__67_, s_r_85__66_, s_r_85__65_, s_r_85__64_, s_r_85__63_, s_r_85__62_, s_r_85__61_, s_r_85__60_, s_r_85__59_, s_r_85__58_, s_r_85__57_, s_r_85__56_, s_r_85__55_, s_r_85__54_, s_r_85__53_, s_r_85__52_, s_r_85__51_, s_r_85__50_, s_r_85__49_, s_r_85__48_, s_r_85__47_, s_r_85__46_, s_r_85__45_, s_r_85__44_, s_r_85__43_, s_r_85__42_, s_r_85__41_, s_r_85__40_, s_r_85__39_, s_r_85__38_, s_r_85__37_, s_r_85__36_, s_r_85__35_, s_r_85__34_, s_r_85__33_, s_r_85__32_, s_r_85__31_, s_r_85__30_, s_r_85__29_, s_r_85__28_, s_r_85__27_, s_r_85__26_, s_r_85__25_, s_r_85__24_, s_r_85__23_, s_r_85__22_, s_r_85__21_, s_r_85__20_, s_r_85__19_, s_r_85__18_, s_r_85__17_, s_r_85__16_, s_r_85__15_, s_r_85__14_, s_r_85__13_, s_r_85__12_, s_r_85__11_, s_r_85__10_, s_r_85__9_, s_r_85__8_, s_r_85__7_, s_r_85__6_, s_r_85__5_, s_r_85__4_, s_r_85__3_, s_r_85__2_, s_r_85__1_, s_r_85__0_ }),
    .c_o(c_r[85]),
    .prod_accum_o({ prod_accum_85__86_, prod_accum_85__85_, prod_accum_85__84_, prod_accum_85__83_, prod_accum_85__82_, prod_accum_85__81_, prod_accum_85__80_, prod_accum_85__79_, prod_accum_85__78_, prod_accum_85__77_, prod_accum_85__76_, prod_accum_85__75_, prod_accum_85__74_, prod_accum_85__73_, prod_accum_85__72_, prod_accum_85__71_, prod_accum_85__70_, prod_accum_85__69_, prod_accum_85__68_, prod_accum_85__67_, prod_accum_85__66_, prod_accum_85__65_, prod_accum_85__64_, prod_accum_85__63_, prod_accum_85__62_, prod_accum_85__61_, prod_accum_85__60_, prod_accum_85__59_, prod_accum_85__58_, prod_accum_85__57_, prod_accum_85__56_, prod_accum_85__55_, prod_accum_85__54_, prod_accum_85__53_, prod_accum_85__52_, prod_accum_85__51_, prod_accum_85__50_, prod_accum_85__49_, prod_accum_85__48_, prod_accum_85__47_, prod_accum_85__46_, prod_accum_85__45_, prod_accum_85__44_, prod_accum_85__43_, prod_accum_85__42_, prod_accum_85__41_, prod_accum_85__40_, prod_accum_85__39_, prod_accum_85__38_, prod_accum_85__37_, prod_accum_85__36_, prod_accum_85__35_, prod_accum_85__34_, prod_accum_85__33_, prod_accum_85__32_, prod_accum_85__31_, prod_accum_85__30_, prod_accum_85__29_, prod_accum_85__28_, prod_accum_85__27_, prod_accum_85__26_, prod_accum_85__25_, prod_accum_85__24_, prod_accum_85__23_, prod_accum_85__22_, prod_accum_85__21_, prod_accum_85__20_, prod_accum_85__19_, prod_accum_85__18_, prod_accum_85__17_, prod_accum_85__16_, prod_accum_85__15_, prod_accum_85__14_, prod_accum_85__13_, prod_accum_85__12_, prod_accum_85__11_, prod_accum_85__10_, prod_accum_85__9_, prod_accum_85__8_, prod_accum_85__7_, prod_accum_85__6_, prod_accum_85__5_, prod_accum_85__4_, prod_accum_85__3_, prod_accum_85__2_, prod_accum_85__1_, prod_accum_85__0_ })
  );


  bsg_mul_array_row_128_86_x
  genblk1_86__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[11007:10880]),
    .b_i(b_r[11007:10880]),
    .s_i({ s_r_85__127_, s_r_85__126_, s_r_85__125_, s_r_85__124_, s_r_85__123_, s_r_85__122_, s_r_85__121_, s_r_85__120_, s_r_85__119_, s_r_85__118_, s_r_85__117_, s_r_85__116_, s_r_85__115_, s_r_85__114_, s_r_85__113_, s_r_85__112_, s_r_85__111_, s_r_85__110_, s_r_85__109_, s_r_85__108_, s_r_85__107_, s_r_85__106_, s_r_85__105_, s_r_85__104_, s_r_85__103_, s_r_85__102_, s_r_85__101_, s_r_85__100_, s_r_85__99_, s_r_85__98_, s_r_85__97_, s_r_85__96_, s_r_85__95_, s_r_85__94_, s_r_85__93_, s_r_85__92_, s_r_85__91_, s_r_85__90_, s_r_85__89_, s_r_85__88_, s_r_85__87_, s_r_85__86_, s_r_85__85_, s_r_85__84_, s_r_85__83_, s_r_85__82_, s_r_85__81_, s_r_85__80_, s_r_85__79_, s_r_85__78_, s_r_85__77_, s_r_85__76_, s_r_85__75_, s_r_85__74_, s_r_85__73_, s_r_85__72_, s_r_85__71_, s_r_85__70_, s_r_85__69_, s_r_85__68_, s_r_85__67_, s_r_85__66_, s_r_85__65_, s_r_85__64_, s_r_85__63_, s_r_85__62_, s_r_85__61_, s_r_85__60_, s_r_85__59_, s_r_85__58_, s_r_85__57_, s_r_85__56_, s_r_85__55_, s_r_85__54_, s_r_85__53_, s_r_85__52_, s_r_85__51_, s_r_85__50_, s_r_85__49_, s_r_85__48_, s_r_85__47_, s_r_85__46_, s_r_85__45_, s_r_85__44_, s_r_85__43_, s_r_85__42_, s_r_85__41_, s_r_85__40_, s_r_85__39_, s_r_85__38_, s_r_85__37_, s_r_85__36_, s_r_85__35_, s_r_85__34_, s_r_85__33_, s_r_85__32_, s_r_85__31_, s_r_85__30_, s_r_85__29_, s_r_85__28_, s_r_85__27_, s_r_85__26_, s_r_85__25_, s_r_85__24_, s_r_85__23_, s_r_85__22_, s_r_85__21_, s_r_85__20_, s_r_85__19_, s_r_85__18_, s_r_85__17_, s_r_85__16_, s_r_85__15_, s_r_85__14_, s_r_85__13_, s_r_85__12_, s_r_85__11_, s_r_85__10_, s_r_85__9_, s_r_85__8_, s_r_85__7_, s_r_85__6_, s_r_85__5_, s_r_85__4_, s_r_85__3_, s_r_85__2_, s_r_85__1_, s_r_85__0_ }),
    .c_i(c_r[85]),
    .prod_accum_i({ prod_accum_85__86_, prod_accum_85__85_, prod_accum_85__84_, prod_accum_85__83_, prod_accum_85__82_, prod_accum_85__81_, prod_accum_85__80_, prod_accum_85__79_, prod_accum_85__78_, prod_accum_85__77_, prod_accum_85__76_, prod_accum_85__75_, prod_accum_85__74_, prod_accum_85__73_, prod_accum_85__72_, prod_accum_85__71_, prod_accum_85__70_, prod_accum_85__69_, prod_accum_85__68_, prod_accum_85__67_, prod_accum_85__66_, prod_accum_85__65_, prod_accum_85__64_, prod_accum_85__63_, prod_accum_85__62_, prod_accum_85__61_, prod_accum_85__60_, prod_accum_85__59_, prod_accum_85__58_, prod_accum_85__57_, prod_accum_85__56_, prod_accum_85__55_, prod_accum_85__54_, prod_accum_85__53_, prod_accum_85__52_, prod_accum_85__51_, prod_accum_85__50_, prod_accum_85__49_, prod_accum_85__48_, prod_accum_85__47_, prod_accum_85__46_, prod_accum_85__45_, prod_accum_85__44_, prod_accum_85__43_, prod_accum_85__42_, prod_accum_85__41_, prod_accum_85__40_, prod_accum_85__39_, prod_accum_85__38_, prod_accum_85__37_, prod_accum_85__36_, prod_accum_85__35_, prod_accum_85__34_, prod_accum_85__33_, prod_accum_85__32_, prod_accum_85__31_, prod_accum_85__30_, prod_accum_85__29_, prod_accum_85__28_, prod_accum_85__27_, prod_accum_85__26_, prod_accum_85__25_, prod_accum_85__24_, prod_accum_85__23_, prod_accum_85__22_, prod_accum_85__21_, prod_accum_85__20_, prod_accum_85__19_, prod_accum_85__18_, prod_accum_85__17_, prod_accum_85__16_, prod_accum_85__15_, prod_accum_85__14_, prod_accum_85__13_, prod_accum_85__12_, prod_accum_85__11_, prod_accum_85__10_, prod_accum_85__9_, prod_accum_85__8_, prod_accum_85__7_, prod_accum_85__6_, prod_accum_85__5_, prod_accum_85__4_, prod_accum_85__3_, prod_accum_85__2_, prod_accum_85__1_, prod_accum_85__0_ }),
    .a_o(a_r[11135:11008]),
    .b_o(b_r[11135:11008]),
    .s_o({ s_r_86__127_, s_r_86__126_, s_r_86__125_, s_r_86__124_, s_r_86__123_, s_r_86__122_, s_r_86__121_, s_r_86__120_, s_r_86__119_, s_r_86__118_, s_r_86__117_, s_r_86__116_, s_r_86__115_, s_r_86__114_, s_r_86__113_, s_r_86__112_, s_r_86__111_, s_r_86__110_, s_r_86__109_, s_r_86__108_, s_r_86__107_, s_r_86__106_, s_r_86__105_, s_r_86__104_, s_r_86__103_, s_r_86__102_, s_r_86__101_, s_r_86__100_, s_r_86__99_, s_r_86__98_, s_r_86__97_, s_r_86__96_, s_r_86__95_, s_r_86__94_, s_r_86__93_, s_r_86__92_, s_r_86__91_, s_r_86__90_, s_r_86__89_, s_r_86__88_, s_r_86__87_, s_r_86__86_, s_r_86__85_, s_r_86__84_, s_r_86__83_, s_r_86__82_, s_r_86__81_, s_r_86__80_, s_r_86__79_, s_r_86__78_, s_r_86__77_, s_r_86__76_, s_r_86__75_, s_r_86__74_, s_r_86__73_, s_r_86__72_, s_r_86__71_, s_r_86__70_, s_r_86__69_, s_r_86__68_, s_r_86__67_, s_r_86__66_, s_r_86__65_, s_r_86__64_, s_r_86__63_, s_r_86__62_, s_r_86__61_, s_r_86__60_, s_r_86__59_, s_r_86__58_, s_r_86__57_, s_r_86__56_, s_r_86__55_, s_r_86__54_, s_r_86__53_, s_r_86__52_, s_r_86__51_, s_r_86__50_, s_r_86__49_, s_r_86__48_, s_r_86__47_, s_r_86__46_, s_r_86__45_, s_r_86__44_, s_r_86__43_, s_r_86__42_, s_r_86__41_, s_r_86__40_, s_r_86__39_, s_r_86__38_, s_r_86__37_, s_r_86__36_, s_r_86__35_, s_r_86__34_, s_r_86__33_, s_r_86__32_, s_r_86__31_, s_r_86__30_, s_r_86__29_, s_r_86__28_, s_r_86__27_, s_r_86__26_, s_r_86__25_, s_r_86__24_, s_r_86__23_, s_r_86__22_, s_r_86__21_, s_r_86__20_, s_r_86__19_, s_r_86__18_, s_r_86__17_, s_r_86__16_, s_r_86__15_, s_r_86__14_, s_r_86__13_, s_r_86__12_, s_r_86__11_, s_r_86__10_, s_r_86__9_, s_r_86__8_, s_r_86__7_, s_r_86__6_, s_r_86__5_, s_r_86__4_, s_r_86__3_, s_r_86__2_, s_r_86__1_, s_r_86__0_ }),
    .c_o(c_r[86]),
    .prod_accum_o({ prod_accum_86__87_, prod_accum_86__86_, prod_accum_86__85_, prod_accum_86__84_, prod_accum_86__83_, prod_accum_86__82_, prod_accum_86__81_, prod_accum_86__80_, prod_accum_86__79_, prod_accum_86__78_, prod_accum_86__77_, prod_accum_86__76_, prod_accum_86__75_, prod_accum_86__74_, prod_accum_86__73_, prod_accum_86__72_, prod_accum_86__71_, prod_accum_86__70_, prod_accum_86__69_, prod_accum_86__68_, prod_accum_86__67_, prod_accum_86__66_, prod_accum_86__65_, prod_accum_86__64_, prod_accum_86__63_, prod_accum_86__62_, prod_accum_86__61_, prod_accum_86__60_, prod_accum_86__59_, prod_accum_86__58_, prod_accum_86__57_, prod_accum_86__56_, prod_accum_86__55_, prod_accum_86__54_, prod_accum_86__53_, prod_accum_86__52_, prod_accum_86__51_, prod_accum_86__50_, prod_accum_86__49_, prod_accum_86__48_, prod_accum_86__47_, prod_accum_86__46_, prod_accum_86__45_, prod_accum_86__44_, prod_accum_86__43_, prod_accum_86__42_, prod_accum_86__41_, prod_accum_86__40_, prod_accum_86__39_, prod_accum_86__38_, prod_accum_86__37_, prod_accum_86__36_, prod_accum_86__35_, prod_accum_86__34_, prod_accum_86__33_, prod_accum_86__32_, prod_accum_86__31_, prod_accum_86__30_, prod_accum_86__29_, prod_accum_86__28_, prod_accum_86__27_, prod_accum_86__26_, prod_accum_86__25_, prod_accum_86__24_, prod_accum_86__23_, prod_accum_86__22_, prod_accum_86__21_, prod_accum_86__20_, prod_accum_86__19_, prod_accum_86__18_, prod_accum_86__17_, prod_accum_86__16_, prod_accum_86__15_, prod_accum_86__14_, prod_accum_86__13_, prod_accum_86__12_, prod_accum_86__11_, prod_accum_86__10_, prod_accum_86__9_, prod_accum_86__8_, prod_accum_86__7_, prod_accum_86__6_, prod_accum_86__5_, prod_accum_86__4_, prod_accum_86__3_, prod_accum_86__2_, prod_accum_86__1_, prod_accum_86__0_ })
  );


  bsg_mul_array_row_128_87_x
  genblk1_87__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[11135:11008]),
    .b_i(b_r[11135:11008]),
    .s_i({ s_r_86__127_, s_r_86__126_, s_r_86__125_, s_r_86__124_, s_r_86__123_, s_r_86__122_, s_r_86__121_, s_r_86__120_, s_r_86__119_, s_r_86__118_, s_r_86__117_, s_r_86__116_, s_r_86__115_, s_r_86__114_, s_r_86__113_, s_r_86__112_, s_r_86__111_, s_r_86__110_, s_r_86__109_, s_r_86__108_, s_r_86__107_, s_r_86__106_, s_r_86__105_, s_r_86__104_, s_r_86__103_, s_r_86__102_, s_r_86__101_, s_r_86__100_, s_r_86__99_, s_r_86__98_, s_r_86__97_, s_r_86__96_, s_r_86__95_, s_r_86__94_, s_r_86__93_, s_r_86__92_, s_r_86__91_, s_r_86__90_, s_r_86__89_, s_r_86__88_, s_r_86__87_, s_r_86__86_, s_r_86__85_, s_r_86__84_, s_r_86__83_, s_r_86__82_, s_r_86__81_, s_r_86__80_, s_r_86__79_, s_r_86__78_, s_r_86__77_, s_r_86__76_, s_r_86__75_, s_r_86__74_, s_r_86__73_, s_r_86__72_, s_r_86__71_, s_r_86__70_, s_r_86__69_, s_r_86__68_, s_r_86__67_, s_r_86__66_, s_r_86__65_, s_r_86__64_, s_r_86__63_, s_r_86__62_, s_r_86__61_, s_r_86__60_, s_r_86__59_, s_r_86__58_, s_r_86__57_, s_r_86__56_, s_r_86__55_, s_r_86__54_, s_r_86__53_, s_r_86__52_, s_r_86__51_, s_r_86__50_, s_r_86__49_, s_r_86__48_, s_r_86__47_, s_r_86__46_, s_r_86__45_, s_r_86__44_, s_r_86__43_, s_r_86__42_, s_r_86__41_, s_r_86__40_, s_r_86__39_, s_r_86__38_, s_r_86__37_, s_r_86__36_, s_r_86__35_, s_r_86__34_, s_r_86__33_, s_r_86__32_, s_r_86__31_, s_r_86__30_, s_r_86__29_, s_r_86__28_, s_r_86__27_, s_r_86__26_, s_r_86__25_, s_r_86__24_, s_r_86__23_, s_r_86__22_, s_r_86__21_, s_r_86__20_, s_r_86__19_, s_r_86__18_, s_r_86__17_, s_r_86__16_, s_r_86__15_, s_r_86__14_, s_r_86__13_, s_r_86__12_, s_r_86__11_, s_r_86__10_, s_r_86__9_, s_r_86__8_, s_r_86__7_, s_r_86__6_, s_r_86__5_, s_r_86__4_, s_r_86__3_, s_r_86__2_, s_r_86__1_, s_r_86__0_ }),
    .c_i(c_r[86]),
    .prod_accum_i({ prod_accum_86__87_, prod_accum_86__86_, prod_accum_86__85_, prod_accum_86__84_, prod_accum_86__83_, prod_accum_86__82_, prod_accum_86__81_, prod_accum_86__80_, prod_accum_86__79_, prod_accum_86__78_, prod_accum_86__77_, prod_accum_86__76_, prod_accum_86__75_, prod_accum_86__74_, prod_accum_86__73_, prod_accum_86__72_, prod_accum_86__71_, prod_accum_86__70_, prod_accum_86__69_, prod_accum_86__68_, prod_accum_86__67_, prod_accum_86__66_, prod_accum_86__65_, prod_accum_86__64_, prod_accum_86__63_, prod_accum_86__62_, prod_accum_86__61_, prod_accum_86__60_, prod_accum_86__59_, prod_accum_86__58_, prod_accum_86__57_, prod_accum_86__56_, prod_accum_86__55_, prod_accum_86__54_, prod_accum_86__53_, prod_accum_86__52_, prod_accum_86__51_, prod_accum_86__50_, prod_accum_86__49_, prod_accum_86__48_, prod_accum_86__47_, prod_accum_86__46_, prod_accum_86__45_, prod_accum_86__44_, prod_accum_86__43_, prod_accum_86__42_, prod_accum_86__41_, prod_accum_86__40_, prod_accum_86__39_, prod_accum_86__38_, prod_accum_86__37_, prod_accum_86__36_, prod_accum_86__35_, prod_accum_86__34_, prod_accum_86__33_, prod_accum_86__32_, prod_accum_86__31_, prod_accum_86__30_, prod_accum_86__29_, prod_accum_86__28_, prod_accum_86__27_, prod_accum_86__26_, prod_accum_86__25_, prod_accum_86__24_, prod_accum_86__23_, prod_accum_86__22_, prod_accum_86__21_, prod_accum_86__20_, prod_accum_86__19_, prod_accum_86__18_, prod_accum_86__17_, prod_accum_86__16_, prod_accum_86__15_, prod_accum_86__14_, prod_accum_86__13_, prod_accum_86__12_, prod_accum_86__11_, prod_accum_86__10_, prod_accum_86__9_, prod_accum_86__8_, prod_accum_86__7_, prod_accum_86__6_, prod_accum_86__5_, prod_accum_86__4_, prod_accum_86__3_, prod_accum_86__2_, prod_accum_86__1_, prod_accum_86__0_ }),
    .a_o(a_r[11263:11136]),
    .b_o(b_r[11263:11136]),
    .s_o({ s_r_87__127_, s_r_87__126_, s_r_87__125_, s_r_87__124_, s_r_87__123_, s_r_87__122_, s_r_87__121_, s_r_87__120_, s_r_87__119_, s_r_87__118_, s_r_87__117_, s_r_87__116_, s_r_87__115_, s_r_87__114_, s_r_87__113_, s_r_87__112_, s_r_87__111_, s_r_87__110_, s_r_87__109_, s_r_87__108_, s_r_87__107_, s_r_87__106_, s_r_87__105_, s_r_87__104_, s_r_87__103_, s_r_87__102_, s_r_87__101_, s_r_87__100_, s_r_87__99_, s_r_87__98_, s_r_87__97_, s_r_87__96_, s_r_87__95_, s_r_87__94_, s_r_87__93_, s_r_87__92_, s_r_87__91_, s_r_87__90_, s_r_87__89_, s_r_87__88_, s_r_87__87_, s_r_87__86_, s_r_87__85_, s_r_87__84_, s_r_87__83_, s_r_87__82_, s_r_87__81_, s_r_87__80_, s_r_87__79_, s_r_87__78_, s_r_87__77_, s_r_87__76_, s_r_87__75_, s_r_87__74_, s_r_87__73_, s_r_87__72_, s_r_87__71_, s_r_87__70_, s_r_87__69_, s_r_87__68_, s_r_87__67_, s_r_87__66_, s_r_87__65_, s_r_87__64_, s_r_87__63_, s_r_87__62_, s_r_87__61_, s_r_87__60_, s_r_87__59_, s_r_87__58_, s_r_87__57_, s_r_87__56_, s_r_87__55_, s_r_87__54_, s_r_87__53_, s_r_87__52_, s_r_87__51_, s_r_87__50_, s_r_87__49_, s_r_87__48_, s_r_87__47_, s_r_87__46_, s_r_87__45_, s_r_87__44_, s_r_87__43_, s_r_87__42_, s_r_87__41_, s_r_87__40_, s_r_87__39_, s_r_87__38_, s_r_87__37_, s_r_87__36_, s_r_87__35_, s_r_87__34_, s_r_87__33_, s_r_87__32_, s_r_87__31_, s_r_87__30_, s_r_87__29_, s_r_87__28_, s_r_87__27_, s_r_87__26_, s_r_87__25_, s_r_87__24_, s_r_87__23_, s_r_87__22_, s_r_87__21_, s_r_87__20_, s_r_87__19_, s_r_87__18_, s_r_87__17_, s_r_87__16_, s_r_87__15_, s_r_87__14_, s_r_87__13_, s_r_87__12_, s_r_87__11_, s_r_87__10_, s_r_87__9_, s_r_87__8_, s_r_87__7_, s_r_87__6_, s_r_87__5_, s_r_87__4_, s_r_87__3_, s_r_87__2_, s_r_87__1_, s_r_87__0_ }),
    .c_o(c_r[87]),
    .prod_accum_o({ prod_accum_87__88_, prod_accum_87__87_, prod_accum_87__86_, prod_accum_87__85_, prod_accum_87__84_, prod_accum_87__83_, prod_accum_87__82_, prod_accum_87__81_, prod_accum_87__80_, prod_accum_87__79_, prod_accum_87__78_, prod_accum_87__77_, prod_accum_87__76_, prod_accum_87__75_, prod_accum_87__74_, prod_accum_87__73_, prod_accum_87__72_, prod_accum_87__71_, prod_accum_87__70_, prod_accum_87__69_, prod_accum_87__68_, prod_accum_87__67_, prod_accum_87__66_, prod_accum_87__65_, prod_accum_87__64_, prod_accum_87__63_, prod_accum_87__62_, prod_accum_87__61_, prod_accum_87__60_, prod_accum_87__59_, prod_accum_87__58_, prod_accum_87__57_, prod_accum_87__56_, prod_accum_87__55_, prod_accum_87__54_, prod_accum_87__53_, prod_accum_87__52_, prod_accum_87__51_, prod_accum_87__50_, prod_accum_87__49_, prod_accum_87__48_, prod_accum_87__47_, prod_accum_87__46_, prod_accum_87__45_, prod_accum_87__44_, prod_accum_87__43_, prod_accum_87__42_, prod_accum_87__41_, prod_accum_87__40_, prod_accum_87__39_, prod_accum_87__38_, prod_accum_87__37_, prod_accum_87__36_, prod_accum_87__35_, prod_accum_87__34_, prod_accum_87__33_, prod_accum_87__32_, prod_accum_87__31_, prod_accum_87__30_, prod_accum_87__29_, prod_accum_87__28_, prod_accum_87__27_, prod_accum_87__26_, prod_accum_87__25_, prod_accum_87__24_, prod_accum_87__23_, prod_accum_87__22_, prod_accum_87__21_, prod_accum_87__20_, prod_accum_87__19_, prod_accum_87__18_, prod_accum_87__17_, prod_accum_87__16_, prod_accum_87__15_, prod_accum_87__14_, prod_accum_87__13_, prod_accum_87__12_, prod_accum_87__11_, prod_accum_87__10_, prod_accum_87__9_, prod_accum_87__8_, prod_accum_87__7_, prod_accum_87__6_, prod_accum_87__5_, prod_accum_87__4_, prod_accum_87__3_, prod_accum_87__2_, prod_accum_87__1_, prod_accum_87__0_ })
  );


  bsg_mul_array_row_128_88_x
  genblk1_88__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[11263:11136]),
    .b_i(b_r[11263:11136]),
    .s_i({ s_r_87__127_, s_r_87__126_, s_r_87__125_, s_r_87__124_, s_r_87__123_, s_r_87__122_, s_r_87__121_, s_r_87__120_, s_r_87__119_, s_r_87__118_, s_r_87__117_, s_r_87__116_, s_r_87__115_, s_r_87__114_, s_r_87__113_, s_r_87__112_, s_r_87__111_, s_r_87__110_, s_r_87__109_, s_r_87__108_, s_r_87__107_, s_r_87__106_, s_r_87__105_, s_r_87__104_, s_r_87__103_, s_r_87__102_, s_r_87__101_, s_r_87__100_, s_r_87__99_, s_r_87__98_, s_r_87__97_, s_r_87__96_, s_r_87__95_, s_r_87__94_, s_r_87__93_, s_r_87__92_, s_r_87__91_, s_r_87__90_, s_r_87__89_, s_r_87__88_, s_r_87__87_, s_r_87__86_, s_r_87__85_, s_r_87__84_, s_r_87__83_, s_r_87__82_, s_r_87__81_, s_r_87__80_, s_r_87__79_, s_r_87__78_, s_r_87__77_, s_r_87__76_, s_r_87__75_, s_r_87__74_, s_r_87__73_, s_r_87__72_, s_r_87__71_, s_r_87__70_, s_r_87__69_, s_r_87__68_, s_r_87__67_, s_r_87__66_, s_r_87__65_, s_r_87__64_, s_r_87__63_, s_r_87__62_, s_r_87__61_, s_r_87__60_, s_r_87__59_, s_r_87__58_, s_r_87__57_, s_r_87__56_, s_r_87__55_, s_r_87__54_, s_r_87__53_, s_r_87__52_, s_r_87__51_, s_r_87__50_, s_r_87__49_, s_r_87__48_, s_r_87__47_, s_r_87__46_, s_r_87__45_, s_r_87__44_, s_r_87__43_, s_r_87__42_, s_r_87__41_, s_r_87__40_, s_r_87__39_, s_r_87__38_, s_r_87__37_, s_r_87__36_, s_r_87__35_, s_r_87__34_, s_r_87__33_, s_r_87__32_, s_r_87__31_, s_r_87__30_, s_r_87__29_, s_r_87__28_, s_r_87__27_, s_r_87__26_, s_r_87__25_, s_r_87__24_, s_r_87__23_, s_r_87__22_, s_r_87__21_, s_r_87__20_, s_r_87__19_, s_r_87__18_, s_r_87__17_, s_r_87__16_, s_r_87__15_, s_r_87__14_, s_r_87__13_, s_r_87__12_, s_r_87__11_, s_r_87__10_, s_r_87__9_, s_r_87__8_, s_r_87__7_, s_r_87__6_, s_r_87__5_, s_r_87__4_, s_r_87__3_, s_r_87__2_, s_r_87__1_, s_r_87__0_ }),
    .c_i(c_r[87]),
    .prod_accum_i({ prod_accum_87__88_, prod_accum_87__87_, prod_accum_87__86_, prod_accum_87__85_, prod_accum_87__84_, prod_accum_87__83_, prod_accum_87__82_, prod_accum_87__81_, prod_accum_87__80_, prod_accum_87__79_, prod_accum_87__78_, prod_accum_87__77_, prod_accum_87__76_, prod_accum_87__75_, prod_accum_87__74_, prod_accum_87__73_, prod_accum_87__72_, prod_accum_87__71_, prod_accum_87__70_, prod_accum_87__69_, prod_accum_87__68_, prod_accum_87__67_, prod_accum_87__66_, prod_accum_87__65_, prod_accum_87__64_, prod_accum_87__63_, prod_accum_87__62_, prod_accum_87__61_, prod_accum_87__60_, prod_accum_87__59_, prod_accum_87__58_, prod_accum_87__57_, prod_accum_87__56_, prod_accum_87__55_, prod_accum_87__54_, prod_accum_87__53_, prod_accum_87__52_, prod_accum_87__51_, prod_accum_87__50_, prod_accum_87__49_, prod_accum_87__48_, prod_accum_87__47_, prod_accum_87__46_, prod_accum_87__45_, prod_accum_87__44_, prod_accum_87__43_, prod_accum_87__42_, prod_accum_87__41_, prod_accum_87__40_, prod_accum_87__39_, prod_accum_87__38_, prod_accum_87__37_, prod_accum_87__36_, prod_accum_87__35_, prod_accum_87__34_, prod_accum_87__33_, prod_accum_87__32_, prod_accum_87__31_, prod_accum_87__30_, prod_accum_87__29_, prod_accum_87__28_, prod_accum_87__27_, prod_accum_87__26_, prod_accum_87__25_, prod_accum_87__24_, prod_accum_87__23_, prod_accum_87__22_, prod_accum_87__21_, prod_accum_87__20_, prod_accum_87__19_, prod_accum_87__18_, prod_accum_87__17_, prod_accum_87__16_, prod_accum_87__15_, prod_accum_87__14_, prod_accum_87__13_, prod_accum_87__12_, prod_accum_87__11_, prod_accum_87__10_, prod_accum_87__9_, prod_accum_87__8_, prod_accum_87__7_, prod_accum_87__6_, prod_accum_87__5_, prod_accum_87__4_, prod_accum_87__3_, prod_accum_87__2_, prod_accum_87__1_, prod_accum_87__0_ }),
    .a_o(a_r[11391:11264]),
    .b_o(b_r[11391:11264]),
    .s_o({ s_r_88__127_, s_r_88__126_, s_r_88__125_, s_r_88__124_, s_r_88__123_, s_r_88__122_, s_r_88__121_, s_r_88__120_, s_r_88__119_, s_r_88__118_, s_r_88__117_, s_r_88__116_, s_r_88__115_, s_r_88__114_, s_r_88__113_, s_r_88__112_, s_r_88__111_, s_r_88__110_, s_r_88__109_, s_r_88__108_, s_r_88__107_, s_r_88__106_, s_r_88__105_, s_r_88__104_, s_r_88__103_, s_r_88__102_, s_r_88__101_, s_r_88__100_, s_r_88__99_, s_r_88__98_, s_r_88__97_, s_r_88__96_, s_r_88__95_, s_r_88__94_, s_r_88__93_, s_r_88__92_, s_r_88__91_, s_r_88__90_, s_r_88__89_, s_r_88__88_, s_r_88__87_, s_r_88__86_, s_r_88__85_, s_r_88__84_, s_r_88__83_, s_r_88__82_, s_r_88__81_, s_r_88__80_, s_r_88__79_, s_r_88__78_, s_r_88__77_, s_r_88__76_, s_r_88__75_, s_r_88__74_, s_r_88__73_, s_r_88__72_, s_r_88__71_, s_r_88__70_, s_r_88__69_, s_r_88__68_, s_r_88__67_, s_r_88__66_, s_r_88__65_, s_r_88__64_, s_r_88__63_, s_r_88__62_, s_r_88__61_, s_r_88__60_, s_r_88__59_, s_r_88__58_, s_r_88__57_, s_r_88__56_, s_r_88__55_, s_r_88__54_, s_r_88__53_, s_r_88__52_, s_r_88__51_, s_r_88__50_, s_r_88__49_, s_r_88__48_, s_r_88__47_, s_r_88__46_, s_r_88__45_, s_r_88__44_, s_r_88__43_, s_r_88__42_, s_r_88__41_, s_r_88__40_, s_r_88__39_, s_r_88__38_, s_r_88__37_, s_r_88__36_, s_r_88__35_, s_r_88__34_, s_r_88__33_, s_r_88__32_, s_r_88__31_, s_r_88__30_, s_r_88__29_, s_r_88__28_, s_r_88__27_, s_r_88__26_, s_r_88__25_, s_r_88__24_, s_r_88__23_, s_r_88__22_, s_r_88__21_, s_r_88__20_, s_r_88__19_, s_r_88__18_, s_r_88__17_, s_r_88__16_, s_r_88__15_, s_r_88__14_, s_r_88__13_, s_r_88__12_, s_r_88__11_, s_r_88__10_, s_r_88__9_, s_r_88__8_, s_r_88__7_, s_r_88__6_, s_r_88__5_, s_r_88__4_, s_r_88__3_, s_r_88__2_, s_r_88__1_, s_r_88__0_ }),
    .c_o(c_r[88]),
    .prod_accum_o({ prod_accum_88__89_, prod_accum_88__88_, prod_accum_88__87_, prod_accum_88__86_, prod_accum_88__85_, prod_accum_88__84_, prod_accum_88__83_, prod_accum_88__82_, prod_accum_88__81_, prod_accum_88__80_, prod_accum_88__79_, prod_accum_88__78_, prod_accum_88__77_, prod_accum_88__76_, prod_accum_88__75_, prod_accum_88__74_, prod_accum_88__73_, prod_accum_88__72_, prod_accum_88__71_, prod_accum_88__70_, prod_accum_88__69_, prod_accum_88__68_, prod_accum_88__67_, prod_accum_88__66_, prod_accum_88__65_, prod_accum_88__64_, prod_accum_88__63_, prod_accum_88__62_, prod_accum_88__61_, prod_accum_88__60_, prod_accum_88__59_, prod_accum_88__58_, prod_accum_88__57_, prod_accum_88__56_, prod_accum_88__55_, prod_accum_88__54_, prod_accum_88__53_, prod_accum_88__52_, prod_accum_88__51_, prod_accum_88__50_, prod_accum_88__49_, prod_accum_88__48_, prod_accum_88__47_, prod_accum_88__46_, prod_accum_88__45_, prod_accum_88__44_, prod_accum_88__43_, prod_accum_88__42_, prod_accum_88__41_, prod_accum_88__40_, prod_accum_88__39_, prod_accum_88__38_, prod_accum_88__37_, prod_accum_88__36_, prod_accum_88__35_, prod_accum_88__34_, prod_accum_88__33_, prod_accum_88__32_, prod_accum_88__31_, prod_accum_88__30_, prod_accum_88__29_, prod_accum_88__28_, prod_accum_88__27_, prod_accum_88__26_, prod_accum_88__25_, prod_accum_88__24_, prod_accum_88__23_, prod_accum_88__22_, prod_accum_88__21_, prod_accum_88__20_, prod_accum_88__19_, prod_accum_88__18_, prod_accum_88__17_, prod_accum_88__16_, prod_accum_88__15_, prod_accum_88__14_, prod_accum_88__13_, prod_accum_88__12_, prod_accum_88__11_, prod_accum_88__10_, prod_accum_88__9_, prod_accum_88__8_, prod_accum_88__7_, prod_accum_88__6_, prod_accum_88__5_, prod_accum_88__4_, prod_accum_88__3_, prod_accum_88__2_, prod_accum_88__1_, prod_accum_88__0_ })
  );


  bsg_mul_array_row_128_89_x
  genblk1_89__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[11391:11264]),
    .b_i(b_r[11391:11264]),
    .s_i({ s_r_88__127_, s_r_88__126_, s_r_88__125_, s_r_88__124_, s_r_88__123_, s_r_88__122_, s_r_88__121_, s_r_88__120_, s_r_88__119_, s_r_88__118_, s_r_88__117_, s_r_88__116_, s_r_88__115_, s_r_88__114_, s_r_88__113_, s_r_88__112_, s_r_88__111_, s_r_88__110_, s_r_88__109_, s_r_88__108_, s_r_88__107_, s_r_88__106_, s_r_88__105_, s_r_88__104_, s_r_88__103_, s_r_88__102_, s_r_88__101_, s_r_88__100_, s_r_88__99_, s_r_88__98_, s_r_88__97_, s_r_88__96_, s_r_88__95_, s_r_88__94_, s_r_88__93_, s_r_88__92_, s_r_88__91_, s_r_88__90_, s_r_88__89_, s_r_88__88_, s_r_88__87_, s_r_88__86_, s_r_88__85_, s_r_88__84_, s_r_88__83_, s_r_88__82_, s_r_88__81_, s_r_88__80_, s_r_88__79_, s_r_88__78_, s_r_88__77_, s_r_88__76_, s_r_88__75_, s_r_88__74_, s_r_88__73_, s_r_88__72_, s_r_88__71_, s_r_88__70_, s_r_88__69_, s_r_88__68_, s_r_88__67_, s_r_88__66_, s_r_88__65_, s_r_88__64_, s_r_88__63_, s_r_88__62_, s_r_88__61_, s_r_88__60_, s_r_88__59_, s_r_88__58_, s_r_88__57_, s_r_88__56_, s_r_88__55_, s_r_88__54_, s_r_88__53_, s_r_88__52_, s_r_88__51_, s_r_88__50_, s_r_88__49_, s_r_88__48_, s_r_88__47_, s_r_88__46_, s_r_88__45_, s_r_88__44_, s_r_88__43_, s_r_88__42_, s_r_88__41_, s_r_88__40_, s_r_88__39_, s_r_88__38_, s_r_88__37_, s_r_88__36_, s_r_88__35_, s_r_88__34_, s_r_88__33_, s_r_88__32_, s_r_88__31_, s_r_88__30_, s_r_88__29_, s_r_88__28_, s_r_88__27_, s_r_88__26_, s_r_88__25_, s_r_88__24_, s_r_88__23_, s_r_88__22_, s_r_88__21_, s_r_88__20_, s_r_88__19_, s_r_88__18_, s_r_88__17_, s_r_88__16_, s_r_88__15_, s_r_88__14_, s_r_88__13_, s_r_88__12_, s_r_88__11_, s_r_88__10_, s_r_88__9_, s_r_88__8_, s_r_88__7_, s_r_88__6_, s_r_88__5_, s_r_88__4_, s_r_88__3_, s_r_88__2_, s_r_88__1_, s_r_88__0_ }),
    .c_i(c_r[88]),
    .prod_accum_i({ prod_accum_88__89_, prod_accum_88__88_, prod_accum_88__87_, prod_accum_88__86_, prod_accum_88__85_, prod_accum_88__84_, prod_accum_88__83_, prod_accum_88__82_, prod_accum_88__81_, prod_accum_88__80_, prod_accum_88__79_, prod_accum_88__78_, prod_accum_88__77_, prod_accum_88__76_, prod_accum_88__75_, prod_accum_88__74_, prod_accum_88__73_, prod_accum_88__72_, prod_accum_88__71_, prod_accum_88__70_, prod_accum_88__69_, prod_accum_88__68_, prod_accum_88__67_, prod_accum_88__66_, prod_accum_88__65_, prod_accum_88__64_, prod_accum_88__63_, prod_accum_88__62_, prod_accum_88__61_, prod_accum_88__60_, prod_accum_88__59_, prod_accum_88__58_, prod_accum_88__57_, prod_accum_88__56_, prod_accum_88__55_, prod_accum_88__54_, prod_accum_88__53_, prod_accum_88__52_, prod_accum_88__51_, prod_accum_88__50_, prod_accum_88__49_, prod_accum_88__48_, prod_accum_88__47_, prod_accum_88__46_, prod_accum_88__45_, prod_accum_88__44_, prod_accum_88__43_, prod_accum_88__42_, prod_accum_88__41_, prod_accum_88__40_, prod_accum_88__39_, prod_accum_88__38_, prod_accum_88__37_, prod_accum_88__36_, prod_accum_88__35_, prod_accum_88__34_, prod_accum_88__33_, prod_accum_88__32_, prod_accum_88__31_, prod_accum_88__30_, prod_accum_88__29_, prod_accum_88__28_, prod_accum_88__27_, prod_accum_88__26_, prod_accum_88__25_, prod_accum_88__24_, prod_accum_88__23_, prod_accum_88__22_, prod_accum_88__21_, prod_accum_88__20_, prod_accum_88__19_, prod_accum_88__18_, prod_accum_88__17_, prod_accum_88__16_, prod_accum_88__15_, prod_accum_88__14_, prod_accum_88__13_, prod_accum_88__12_, prod_accum_88__11_, prod_accum_88__10_, prod_accum_88__9_, prod_accum_88__8_, prod_accum_88__7_, prod_accum_88__6_, prod_accum_88__5_, prod_accum_88__4_, prod_accum_88__3_, prod_accum_88__2_, prod_accum_88__1_, prod_accum_88__0_ }),
    .a_o(a_r[11519:11392]),
    .b_o(b_r[11519:11392]),
    .s_o({ s_r_89__127_, s_r_89__126_, s_r_89__125_, s_r_89__124_, s_r_89__123_, s_r_89__122_, s_r_89__121_, s_r_89__120_, s_r_89__119_, s_r_89__118_, s_r_89__117_, s_r_89__116_, s_r_89__115_, s_r_89__114_, s_r_89__113_, s_r_89__112_, s_r_89__111_, s_r_89__110_, s_r_89__109_, s_r_89__108_, s_r_89__107_, s_r_89__106_, s_r_89__105_, s_r_89__104_, s_r_89__103_, s_r_89__102_, s_r_89__101_, s_r_89__100_, s_r_89__99_, s_r_89__98_, s_r_89__97_, s_r_89__96_, s_r_89__95_, s_r_89__94_, s_r_89__93_, s_r_89__92_, s_r_89__91_, s_r_89__90_, s_r_89__89_, s_r_89__88_, s_r_89__87_, s_r_89__86_, s_r_89__85_, s_r_89__84_, s_r_89__83_, s_r_89__82_, s_r_89__81_, s_r_89__80_, s_r_89__79_, s_r_89__78_, s_r_89__77_, s_r_89__76_, s_r_89__75_, s_r_89__74_, s_r_89__73_, s_r_89__72_, s_r_89__71_, s_r_89__70_, s_r_89__69_, s_r_89__68_, s_r_89__67_, s_r_89__66_, s_r_89__65_, s_r_89__64_, s_r_89__63_, s_r_89__62_, s_r_89__61_, s_r_89__60_, s_r_89__59_, s_r_89__58_, s_r_89__57_, s_r_89__56_, s_r_89__55_, s_r_89__54_, s_r_89__53_, s_r_89__52_, s_r_89__51_, s_r_89__50_, s_r_89__49_, s_r_89__48_, s_r_89__47_, s_r_89__46_, s_r_89__45_, s_r_89__44_, s_r_89__43_, s_r_89__42_, s_r_89__41_, s_r_89__40_, s_r_89__39_, s_r_89__38_, s_r_89__37_, s_r_89__36_, s_r_89__35_, s_r_89__34_, s_r_89__33_, s_r_89__32_, s_r_89__31_, s_r_89__30_, s_r_89__29_, s_r_89__28_, s_r_89__27_, s_r_89__26_, s_r_89__25_, s_r_89__24_, s_r_89__23_, s_r_89__22_, s_r_89__21_, s_r_89__20_, s_r_89__19_, s_r_89__18_, s_r_89__17_, s_r_89__16_, s_r_89__15_, s_r_89__14_, s_r_89__13_, s_r_89__12_, s_r_89__11_, s_r_89__10_, s_r_89__9_, s_r_89__8_, s_r_89__7_, s_r_89__6_, s_r_89__5_, s_r_89__4_, s_r_89__3_, s_r_89__2_, s_r_89__1_, s_r_89__0_ }),
    .c_o(c_r[89]),
    .prod_accum_o({ prod_accum_89__90_, prod_accum_89__89_, prod_accum_89__88_, prod_accum_89__87_, prod_accum_89__86_, prod_accum_89__85_, prod_accum_89__84_, prod_accum_89__83_, prod_accum_89__82_, prod_accum_89__81_, prod_accum_89__80_, prod_accum_89__79_, prod_accum_89__78_, prod_accum_89__77_, prod_accum_89__76_, prod_accum_89__75_, prod_accum_89__74_, prod_accum_89__73_, prod_accum_89__72_, prod_accum_89__71_, prod_accum_89__70_, prod_accum_89__69_, prod_accum_89__68_, prod_accum_89__67_, prod_accum_89__66_, prod_accum_89__65_, prod_accum_89__64_, prod_accum_89__63_, prod_accum_89__62_, prod_accum_89__61_, prod_accum_89__60_, prod_accum_89__59_, prod_accum_89__58_, prod_accum_89__57_, prod_accum_89__56_, prod_accum_89__55_, prod_accum_89__54_, prod_accum_89__53_, prod_accum_89__52_, prod_accum_89__51_, prod_accum_89__50_, prod_accum_89__49_, prod_accum_89__48_, prod_accum_89__47_, prod_accum_89__46_, prod_accum_89__45_, prod_accum_89__44_, prod_accum_89__43_, prod_accum_89__42_, prod_accum_89__41_, prod_accum_89__40_, prod_accum_89__39_, prod_accum_89__38_, prod_accum_89__37_, prod_accum_89__36_, prod_accum_89__35_, prod_accum_89__34_, prod_accum_89__33_, prod_accum_89__32_, prod_accum_89__31_, prod_accum_89__30_, prod_accum_89__29_, prod_accum_89__28_, prod_accum_89__27_, prod_accum_89__26_, prod_accum_89__25_, prod_accum_89__24_, prod_accum_89__23_, prod_accum_89__22_, prod_accum_89__21_, prod_accum_89__20_, prod_accum_89__19_, prod_accum_89__18_, prod_accum_89__17_, prod_accum_89__16_, prod_accum_89__15_, prod_accum_89__14_, prod_accum_89__13_, prod_accum_89__12_, prod_accum_89__11_, prod_accum_89__10_, prod_accum_89__9_, prod_accum_89__8_, prod_accum_89__7_, prod_accum_89__6_, prod_accum_89__5_, prod_accum_89__4_, prod_accum_89__3_, prod_accum_89__2_, prod_accum_89__1_, prod_accum_89__0_ })
  );


  bsg_mul_array_row_128_90_x
  genblk1_90__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[11519:11392]),
    .b_i(b_r[11519:11392]),
    .s_i({ s_r_89__127_, s_r_89__126_, s_r_89__125_, s_r_89__124_, s_r_89__123_, s_r_89__122_, s_r_89__121_, s_r_89__120_, s_r_89__119_, s_r_89__118_, s_r_89__117_, s_r_89__116_, s_r_89__115_, s_r_89__114_, s_r_89__113_, s_r_89__112_, s_r_89__111_, s_r_89__110_, s_r_89__109_, s_r_89__108_, s_r_89__107_, s_r_89__106_, s_r_89__105_, s_r_89__104_, s_r_89__103_, s_r_89__102_, s_r_89__101_, s_r_89__100_, s_r_89__99_, s_r_89__98_, s_r_89__97_, s_r_89__96_, s_r_89__95_, s_r_89__94_, s_r_89__93_, s_r_89__92_, s_r_89__91_, s_r_89__90_, s_r_89__89_, s_r_89__88_, s_r_89__87_, s_r_89__86_, s_r_89__85_, s_r_89__84_, s_r_89__83_, s_r_89__82_, s_r_89__81_, s_r_89__80_, s_r_89__79_, s_r_89__78_, s_r_89__77_, s_r_89__76_, s_r_89__75_, s_r_89__74_, s_r_89__73_, s_r_89__72_, s_r_89__71_, s_r_89__70_, s_r_89__69_, s_r_89__68_, s_r_89__67_, s_r_89__66_, s_r_89__65_, s_r_89__64_, s_r_89__63_, s_r_89__62_, s_r_89__61_, s_r_89__60_, s_r_89__59_, s_r_89__58_, s_r_89__57_, s_r_89__56_, s_r_89__55_, s_r_89__54_, s_r_89__53_, s_r_89__52_, s_r_89__51_, s_r_89__50_, s_r_89__49_, s_r_89__48_, s_r_89__47_, s_r_89__46_, s_r_89__45_, s_r_89__44_, s_r_89__43_, s_r_89__42_, s_r_89__41_, s_r_89__40_, s_r_89__39_, s_r_89__38_, s_r_89__37_, s_r_89__36_, s_r_89__35_, s_r_89__34_, s_r_89__33_, s_r_89__32_, s_r_89__31_, s_r_89__30_, s_r_89__29_, s_r_89__28_, s_r_89__27_, s_r_89__26_, s_r_89__25_, s_r_89__24_, s_r_89__23_, s_r_89__22_, s_r_89__21_, s_r_89__20_, s_r_89__19_, s_r_89__18_, s_r_89__17_, s_r_89__16_, s_r_89__15_, s_r_89__14_, s_r_89__13_, s_r_89__12_, s_r_89__11_, s_r_89__10_, s_r_89__9_, s_r_89__8_, s_r_89__7_, s_r_89__6_, s_r_89__5_, s_r_89__4_, s_r_89__3_, s_r_89__2_, s_r_89__1_, s_r_89__0_ }),
    .c_i(c_r[89]),
    .prod_accum_i({ prod_accum_89__90_, prod_accum_89__89_, prod_accum_89__88_, prod_accum_89__87_, prod_accum_89__86_, prod_accum_89__85_, prod_accum_89__84_, prod_accum_89__83_, prod_accum_89__82_, prod_accum_89__81_, prod_accum_89__80_, prod_accum_89__79_, prod_accum_89__78_, prod_accum_89__77_, prod_accum_89__76_, prod_accum_89__75_, prod_accum_89__74_, prod_accum_89__73_, prod_accum_89__72_, prod_accum_89__71_, prod_accum_89__70_, prod_accum_89__69_, prod_accum_89__68_, prod_accum_89__67_, prod_accum_89__66_, prod_accum_89__65_, prod_accum_89__64_, prod_accum_89__63_, prod_accum_89__62_, prod_accum_89__61_, prod_accum_89__60_, prod_accum_89__59_, prod_accum_89__58_, prod_accum_89__57_, prod_accum_89__56_, prod_accum_89__55_, prod_accum_89__54_, prod_accum_89__53_, prod_accum_89__52_, prod_accum_89__51_, prod_accum_89__50_, prod_accum_89__49_, prod_accum_89__48_, prod_accum_89__47_, prod_accum_89__46_, prod_accum_89__45_, prod_accum_89__44_, prod_accum_89__43_, prod_accum_89__42_, prod_accum_89__41_, prod_accum_89__40_, prod_accum_89__39_, prod_accum_89__38_, prod_accum_89__37_, prod_accum_89__36_, prod_accum_89__35_, prod_accum_89__34_, prod_accum_89__33_, prod_accum_89__32_, prod_accum_89__31_, prod_accum_89__30_, prod_accum_89__29_, prod_accum_89__28_, prod_accum_89__27_, prod_accum_89__26_, prod_accum_89__25_, prod_accum_89__24_, prod_accum_89__23_, prod_accum_89__22_, prod_accum_89__21_, prod_accum_89__20_, prod_accum_89__19_, prod_accum_89__18_, prod_accum_89__17_, prod_accum_89__16_, prod_accum_89__15_, prod_accum_89__14_, prod_accum_89__13_, prod_accum_89__12_, prod_accum_89__11_, prod_accum_89__10_, prod_accum_89__9_, prod_accum_89__8_, prod_accum_89__7_, prod_accum_89__6_, prod_accum_89__5_, prod_accum_89__4_, prod_accum_89__3_, prod_accum_89__2_, prod_accum_89__1_, prod_accum_89__0_ }),
    .a_o(a_r[11647:11520]),
    .b_o(b_r[11647:11520]),
    .s_o({ s_r_90__127_, s_r_90__126_, s_r_90__125_, s_r_90__124_, s_r_90__123_, s_r_90__122_, s_r_90__121_, s_r_90__120_, s_r_90__119_, s_r_90__118_, s_r_90__117_, s_r_90__116_, s_r_90__115_, s_r_90__114_, s_r_90__113_, s_r_90__112_, s_r_90__111_, s_r_90__110_, s_r_90__109_, s_r_90__108_, s_r_90__107_, s_r_90__106_, s_r_90__105_, s_r_90__104_, s_r_90__103_, s_r_90__102_, s_r_90__101_, s_r_90__100_, s_r_90__99_, s_r_90__98_, s_r_90__97_, s_r_90__96_, s_r_90__95_, s_r_90__94_, s_r_90__93_, s_r_90__92_, s_r_90__91_, s_r_90__90_, s_r_90__89_, s_r_90__88_, s_r_90__87_, s_r_90__86_, s_r_90__85_, s_r_90__84_, s_r_90__83_, s_r_90__82_, s_r_90__81_, s_r_90__80_, s_r_90__79_, s_r_90__78_, s_r_90__77_, s_r_90__76_, s_r_90__75_, s_r_90__74_, s_r_90__73_, s_r_90__72_, s_r_90__71_, s_r_90__70_, s_r_90__69_, s_r_90__68_, s_r_90__67_, s_r_90__66_, s_r_90__65_, s_r_90__64_, s_r_90__63_, s_r_90__62_, s_r_90__61_, s_r_90__60_, s_r_90__59_, s_r_90__58_, s_r_90__57_, s_r_90__56_, s_r_90__55_, s_r_90__54_, s_r_90__53_, s_r_90__52_, s_r_90__51_, s_r_90__50_, s_r_90__49_, s_r_90__48_, s_r_90__47_, s_r_90__46_, s_r_90__45_, s_r_90__44_, s_r_90__43_, s_r_90__42_, s_r_90__41_, s_r_90__40_, s_r_90__39_, s_r_90__38_, s_r_90__37_, s_r_90__36_, s_r_90__35_, s_r_90__34_, s_r_90__33_, s_r_90__32_, s_r_90__31_, s_r_90__30_, s_r_90__29_, s_r_90__28_, s_r_90__27_, s_r_90__26_, s_r_90__25_, s_r_90__24_, s_r_90__23_, s_r_90__22_, s_r_90__21_, s_r_90__20_, s_r_90__19_, s_r_90__18_, s_r_90__17_, s_r_90__16_, s_r_90__15_, s_r_90__14_, s_r_90__13_, s_r_90__12_, s_r_90__11_, s_r_90__10_, s_r_90__9_, s_r_90__8_, s_r_90__7_, s_r_90__6_, s_r_90__5_, s_r_90__4_, s_r_90__3_, s_r_90__2_, s_r_90__1_, s_r_90__0_ }),
    .c_o(c_r[90]),
    .prod_accum_o({ prod_accum_90__91_, prod_accum_90__90_, prod_accum_90__89_, prod_accum_90__88_, prod_accum_90__87_, prod_accum_90__86_, prod_accum_90__85_, prod_accum_90__84_, prod_accum_90__83_, prod_accum_90__82_, prod_accum_90__81_, prod_accum_90__80_, prod_accum_90__79_, prod_accum_90__78_, prod_accum_90__77_, prod_accum_90__76_, prod_accum_90__75_, prod_accum_90__74_, prod_accum_90__73_, prod_accum_90__72_, prod_accum_90__71_, prod_accum_90__70_, prod_accum_90__69_, prod_accum_90__68_, prod_accum_90__67_, prod_accum_90__66_, prod_accum_90__65_, prod_accum_90__64_, prod_accum_90__63_, prod_accum_90__62_, prod_accum_90__61_, prod_accum_90__60_, prod_accum_90__59_, prod_accum_90__58_, prod_accum_90__57_, prod_accum_90__56_, prod_accum_90__55_, prod_accum_90__54_, prod_accum_90__53_, prod_accum_90__52_, prod_accum_90__51_, prod_accum_90__50_, prod_accum_90__49_, prod_accum_90__48_, prod_accum_90__47_, prod_accum_90__46_, prod_accum_90__45_, prod_accum_90__44_, prod_accum_90__43_, prod_accum_90__42_, prod_accum_90__41_, prod_accum_90__40_, prod_accum_90__39_, prod_accum_90__38_, prod_accum_90__37_, prod_accum_90__36_, prod_accum_90__35_, prod_accum_90__34_, prod_accum_90__33_, prod_accum_90__32_, prod_accum_90__31_, prod_accum_90__30_, prod_accum_90__29_, prod_accum_90__28_, prod_accum_90__27_, prod_accum_90__26_, prod_accum_90__25_, prod_accum_90__24_, prod_accum_90__23_, prod_accum_90__22_, prod_accum_90__21_, prod_accum_90__20_, prod_accum_90__19_, prod_accum_90__18_, prod_accum_90__17_, prod_accum_90__16_, prod_accum_90__15_, prod_accum_90__14_, prod_accum_90__13_, prod_accum_90__12_, prod_accum_90__11_, prod_accum_90__10_, prod_accum_90__9_, prod_accum_90__8_, prod_accum_90__7_, prod_accum_90__6_, prod_accum_90__5_, prod_accum_90__4_, prod_accum_90__3_, prod_accum_90__2_, prod_accum_90__1_, prod_accum_90__0_ })
  );


  bsg_mul_array_row_128_91_x
  genblk1_91__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[11647:11520]),
    .b_i(b_r[11647:11520]),
    .s_i({ s_r_90__127_, s_r_90__126_, s_r_90__125_, s_r_90__124_, s_r_90__123_, s_r_90__122_, s_r_90__121_, s_r_90__120_, s_r_90__119_, s_r_90__118_, s_r_90__117_, s_r_90__116_, s_r_90__115_, s_r_90__114_, s_r_90__113_, s_r_90__112_, s_r_90__111_, s_r_90__110_, s_r_90__109_, s_r_90__108_, s_r_90__107_, s_r_90__106_, s_r_90__105_, s_r_90__104_, s_r_90__103_, s_r_90__102_, s_r_90__101_, s_r_90__100_, s_r_90__99_, s_r_90__98_, s_r_90__97_, s_r_90__96_, s_r_90__95_, s_r_90__94_, s_r_90__93_, s_r_90__92_, s_r_90__91_, s_r_90__90_, s_r_90__89_, s_r_90__88_, s_r_90__87_, s_r_90__86_, s_r_90__85_, s_r_90__84_, s_r_90__83_, s_r_90__82_, s_r_90__81_, s_r_90__80_, s_r_90__79_, s_r_90__78_, s_r_90__77_, s_r_90__76_, s_r_90__75_, s_r_90__74_, s_r_90__73_, s_r_90__72_, s_r_90__71_, s_r_90__70_, s_r_90__69_, s_r_90__68_, s_r_90__67_, s_r_90__66_, s_r_90__65_, s_r_90__64_, s_r_90__63_, s_r_90__62_, s_r_90__61_, s_r_90__60_, s_r_90__59_, s_r_90__58_, s_r_90__57_, s_r_90__56_, s_r_90__55_, s_r_90__54_, s_r_90__53_, s_r_90__52_, s_r_90__51_, s_r_90__50_, s_r_90__49_, s_r_90__48_, s_r_90__47_, s_r_90__46_, s_r_90__45_, s_r_90__44_, s_r_90__43_, s_r_90__42_, s_r_90__41_, s_r_90__40_, s_r_90__39_, s_r_90__38_, s_r_90__37_, s_r_90__36_, s_r_90__35_, s_r_90__34_, s_r_90__33_, s_r_90__32_, s_r_90__31_, s_r_90__30_, s_r_90__29_, s_r_90__28_, s_r_90__27_, s_r_90__26_, s_r_90__25_, s_r_90__24_, s_r_90__23_, s_r_90__22_, s_r_90__21_, s_r_90__20_, s_r_90__19_, s_r_90__18_, s_r_90__17_, s_r_90__16_, s_r_90__15_, s_r_90__14_, s_r_90__13_, s_r_90__12_, s_r_90__11_, s_r_90__10_, s_r_90__9_, s_r_90__8_, s_r_90__7_, s_r_90__6_, s_r_90__5_, s_r_90__4_, s_r_90__3_, s_r_90__2_, s_r_90__1_, s_r_90__0_ }),
    .c_i(c_r[90]),
    .prod_accum_i({ prod_accum_90__91_, prod_accum_90__90_, prod_accum_90__89_, prod_accum_90__88_, prod_accum_90__87_, prod_accum_90__86_, prod_accum_90__85_, prod_accum_90__84_, prod_accum_90__83_, prod_accum_90__82_, prod_accum_90__81_, prod_accum_90__80_, prod_accum_90__79_, prod_accum_90__78_, prod_accum_90__77_, prod_accum_90__76_, prod_accum_90__75_, prod_accum_90__74_, prod_accum_90__73_, prod_accum_90__72_, prod_accum_90__71_, prod_accum_90__70_, prod_accum_90__69_, prod_accum_90__68_, prod_accum_90__67_, prod_accum_90__66_, prod_accum_90__65_, prod_accum_90__64_, prod_accum_90__63_, prod_accum_90__62_, prod_accum_90__61_, prod_accum_90__60_, prod_accum_90__59_, prod_accum_90__58_, prod_accum_90__57_, prod_accum_90__56_, prod_accum_90__55_, prod_accum_90__54_, prod_accum_90__53_, prod_accum_90__52_, prod_accum_90__51_, prod_accum_90__50_, prod_accum_90__49_, prod_accum_90__48_, prod_accum_90__47_, prod_accum_90__46_, prod_accum_90__45_, prod_accum_90__44_, prod_accum_90__43_, prod_accum_90__42_, prod_accum_90__41_, prod_accum_90__40_, prod_accum_90__39_, prod_accum_90__38_, prod_accum_90__37_, prod_accum_90__36_, prod_accum_90__35_, prod_accum_90__34_, prod_accum_90__33_, prod_accum_90__32_, prod_accum_90__31_, prod_accum_90__30_, prod_accum_90__29_, prod_accum_90__28_, prod_accum_90__27_, prod_accum_90__26_, prod_accum_90__25_, prod_accum_90__24_, prod_accum_90__23_, prod_accum_90__22_, prod_accum_90__21_, prod_accum_90__20_, prod_accum_90__19_, prod_accum_90__18_, prod_accum_90__17_, prod_accum_90__16_, prod_accum_90__15_, prod_accum_90__14_, prod_accum_90__13_, prod_accum_90__12_, prod_accum_90__11_, prod_accum_90__10_, prod_accum_90__9_, prod_accum_90__8_, prod_accum_90__7_, prod_accum_90__6_, prod_accum_90__5_, prod_accum_90__4_, prod_accum_90__3_, prod_accum_90__2_, prod_accum_90__1_, prod_accum_90__0_ }),
    .a_o(a_r[11775:11648]),
    .b_o(b_r[11775:11648]),
    .s_o({ s_r_91__127_, s_r_91__126_, s_r_91__125_, s_r_91__124_, s_r_91__123_, s_r_91__122_, s_r_91__121_, s_r_91__120_, s_r_91__119_, s_r_91__118_, s_r_91__117_, s_r_91__116_, s_r_91__115_, s_r_91__114_, s_r_91__113_, s_r_91__112_, s_r_91__111_, s_r_91__110_, s_r_91__109_, s_r_91__108_, s_r_91__107_, s_r_91__106_, s_r_91__105_, s_r_91__104_, s_r_91__103_, s_r_91__102_, s_r_91__101_, s_r_91__100_, s_r_91__99_, s_r_91__98_, s_r_91__97_, s_r_91__96_, s_r_91__95_, s_r_91__94_, s_r_91__93_, s_r_91__92_, s_r_91__91_, s_r_91__90_, s_r_91__89_, s_r_91__88_, s_r_91__87_, s_r_91__86_, s_r_91__85_, s_r_91__84_, s_r_91__83_, s_r_91__82_, s_r_91__81_, s_r_91__80_, s_r_91__79_, s_r_91__78_, s_r_91__77_, s_r_91__76_, s_r_91__75_, s_r_91__74_, s_r_91__73_, s_r_91__72_, s_r_91__71_, s_r_91__70_, s_r_91__69_, s_r_91__68_, s_r_91__67_, s_r_91__66_, s_r_91__65_, s_r_91__64_, s_r_91__63_, s_r_91__62_, s_r_91__61_, s_r_91__60_, s_r_91__59_, s_r_91__58_, s_r_91__57_, s_r_91__56_, s_r_91__55_, s_r_91__54_, s_r_91__53_, s_r_91__52_, s_r_91__51_, s_r_91__50_, s_r_91__49_, s_r_91__48_, s_r_91__47_, s_r_91__46_, s_r_91__45_, s_r_91__44_, s_r_91__43_, s_r_91__42_, s_r_91__41_, s_r_91__40_, s_r_91__39_, s_r_91__38_, s_r_91__37_, s_r_91__36_, s_r_91__35_, s_r_91__34_, s_r_91__33_, s_r_91__32_, s_r_91__31_, s_r_91__30_, s_r_91__29_, s_r_91__28_, s_r_91__27_, s_r_91__26_, s_r_91__25_, s_r_91__24_, s_r_91__23_, s_r_91__22_, s_r_91__21_, s_r_91__20_, s_r_91__19_, s_r_91__18_, s_r_91__17_, s_r_91__16_, s_r_91__15_, s_r_91__14_, s_r_91__13_, s_r_91__12_, s_r_91__11_, s_r_91__10_, s_r_91__9_, s_r_91__8_, s_r_91__7_, s_r_91__6_, s_r_91__5_, s_r_91__4_, s_r_91__3_, s_r_91__2_, s_r_91__1_, s_r_91__0_ }),
    .c_o(c_r[91]),
    .prod_accum_o({ prod_accum_91__92_, prod_accum_91__91_, prod_accum_91__90_, prod_accum_91__89_, prod_accum_91__88_, prod_accum_91__87_, prod_accum_91__86_, prod_accum_91__85_, prod_accum_91__84_, prod_accum_91__83_, prod_accum_91__82_, prod_accum_91__81_, prod_accum_91__80_, prod_accum_91__79_, prod_accum_91__78_, prod_accum_91__77_, prod_accum_91__76_, prod_accum_91__75_, prod_accum_91__74_, prod_accum_91__73_, prod_accum_91__72_, prod_accum_91__71_, prod_accum_91__70_, prod_accum_91__69_, prod_accum_91__68_, prod_accum_91__67_, prod_accum_91__66_, prod_accum_91__65_, prod_accum_91__64_, prod_accum_91__63_, prod_accum_91__62_, prod_accum_91__61_, prod_accum_91__60_, prod_accum_91__59_, prod_accum_91__58_, prod_accum_91__57_, prod_accum_91__56_, prod_accum_91__55_, prod_accum_91__54_, prod_accum_91__53_, prod_accum_91__52_, prod_accum_91__51_, prod_accum_91__50_, prod_accum_91__49_, prod_accum_91__48_, prod_accum_91__47_, prod_accum_91__46_, prod_accum_91__45_, prod_accum_91__44_, prod_accum_91__43_, prod_accum_91__42_, prod_accum_91__41_, prod_accum_91__40_, prod_accum_91__39_, prod_accum_91__38_, prod_accum_91__37_, prod_accum_91__36_, prod_accum_91__35_, prod_accum_91__34_, prod_accum_91__33_, prod_accum_91__32_, prod_accum_91__31_, prod_accum_91__30_, prod_accum_91__29_, prod_accum_91__28_, prod_accum_91__27_, prod_accum_91__26_, prod_accum_91__25_, prod_accum_91__24_, prod_accum_91__23_, prod_accum_91__22_, prod_accum_91__21_, prod_accum_91__20_, prod_accum_91__19_, prod_accum_91__18_, prod_accum_91__17_, prod_accum_91__16_, prod_accum_91__15_, prod_accum_91__14_, prod_accum_91__13_, prod_accum_91__12_, prod_accum_91__11_, prod_accum_91__10_, prod_accum_91__9_, prod_accum_91__8_, prod_accum_91__7_, prod_accum_91__6_, prod_accum_91__5_, prod_accum_91__4_, prod_accum_91__3_, prod_accum_91__2_, prod_accum_91__1_, prod_accum_91__0_ })
  );


  bsg_mul_array_row_128_92_x
  genblk1_92__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[11775:11648]),
    .b_i(b_r[11775:11648]),
    .s_i({ s_r_91__127_, s_r_91__126_, s_r_91__125_, s_r_91__124_, s_r_91__123_, s_r_91__122_, s_r_91__121_, s_r_91__120_, s_r_91__119_, s_r_91__118_, s_r_91__117_, s_r_91__116_, s_r_91__115_, s_r_91__114_, s_r_91__113_, s_r_91__112_, s_r_91__111_, s_r_91__110_, s_r_91__109_, s_r_91__108_, s_r_91__107_, s_r_91__106_, s_r_91__105_, s_r_91__104_, s_r_91__103_, s_r_91__102_, s_r_91__101_, s_r_91__100_, s_r_91__99_, s_r_91__98_, s_r_91__97_, s_r_91__96_, s_r_91__95_, s_r_91__94_, s_r_91__93_, s_r_91__92_, s_r_91__91_, s_r_91__90_, s_r_91__89_, s_r_91__88_, s_r_91__87_, s_r_91__86_, s_r_91__85_, s_r_91__84_, s_r_91__83_, s_r_91__82_, s_r_91__81_, s_r_91__80_, s_r_91__79_, s_r_91__78_, s_r_91__77_, s_r_91__76_, s_r_91__75_, s_r_91__74_, s_r_91__73_, s_r_91__72_, s_r_91__71_, s_r_91__70_, s_r_91__69_, s_r_91__68_, s_r_91__67_, s_r_91__66_, s_r_91__65_, s_r_91__64_, s_r_91__63_, s_r_91__62_, s_r_91__61_, s_r_91__60_, s_r_91__59_, s_r_91__58_, s_r_91__57_, s_r_91__56_, s_r_91__55_, s_r_91__54_, s_r_91__53_, s_r_91__52_, s_r_91__51_, s_r_91__50_, s_r_91__49_, s_r_91__48_, s_r_91__47_, s_r_91__46_, s_r_91__45_, s_r_91__44_, s_r_91__43_, s_r_91__42_, s_r_91__41_, s_r_91__40_, s_r_91__39_, s_r_91__38_, s_r_91__37_, s_r_91__36_, s_r_91__35_, s_r_91__34_, s_r_91__33_, s_r_91__32_, s_r_91__31_, s_r_91__30_, s_r_91__29_, s_r_91__28_, s_r_91__27_, s_r_91__26_, s_r_91__25_, s_r_91__24_, s_r_91__23_, s_r_91__22_, s_r_91__21_, s_r_91__20_, s_r_91__19_, s_r_91__18_, s_r_91__17_, s_r_91__16_, s_r_91__15_, s_r_91__14_, s_r_91__13_, s_r_91__12_, s_r_91__11_, s_r_91__10_, s_r_91__9_, s_r_91__8_, s_r_91__7_, s_r_91__6_, s_r_91__5_, s_r_91__4_, s_r_91__3_, s_r_91__2_, s_r_91__1_, s_r_91__0_ }),
    .c_i(c_r[91]),
    .prod_accum_i({ prod_accum_91__92_, prod_accum_91__91_, prod_accum_91__90_, prod_accum_91__89_, prod_accum_91__88_, prod_accum_91__87_, prod_accum_91__86_, prod_accum_91__85_, prod_accum_91__84_, prod_accum_91__83_, prod_accum_91__82_, prod_accum_91__81_, prod_accum_91__80_, prod_accum_91__79_, prod_accum_91__78_, prod_accum_91__77_, prod_accum_91__76_, prod_accum_91__75_, prod_accum_91__74_, prod_accum_91__73_, prod_accum_91__72_, prod_accum_91__71_, prod_accum_91__70_, prod_accum_91__69_, prod_accum_91__68_, prod_accum_91__67_, prod_accum_91__66_, prod_accum_91__65_, prod_accum_91__64_, prod_accum_91__63_, prod_accum_91__62_, prod_accum_91__61_, prod_accum_91__60_, prod_accum_91__59_, prod_accum_91__58_, prod_accum_91__57_, prod_accum_91__56_, prod_accum_91__55_, prod_accum_91__54_, prod_accum_91__53_, prod_accum_91__52_, prod_accum_91__51_, prod_accum_91__50_, prod_accum_91__49_, prod_accum_91__48_, prod_accum_91__47_, prod_accum_91__46_, prod_accum_91__45_, prod_accum_91__44_, prod_accum_91__43_, prod_accum_91__42_, prod_accum_91__41_, prod_accum_91__40_, prod_accum_91__39_, prod_accum_91__38_, prod_accum_91__37_, prod_accum_91__36_, prod_accum_91__35_, prod_accum_91__34_, prod_accum_91__33_, prod_accum_91__32_, prod_accum_91__31_, prod_accum_91__30_, prod_accum_91__29_, prod_accum_91__28_, prod_accum_91__27_, prod_accum_91__26_, prod_accum_91__25_, prod_accum_91__24_, prod_accum_91__23_, prod_accum_91__22_, prod_accum_91__21_, prod_accum_91__20_, prod_accum_91__19_, prod_accum_91__18_, prod_accum_91__17_, prod_accum_91__16_, prod_accum_91__15_, prod_accum_91__14_, prod_accum_91__13_, prod_accum_91__12_, prod_accum_91__11_, prod_accum_91__10_, prod_accum_91__9_, prod_accum_91__8_, prod_accum_91__7_, prod_accum_91__6_, prod_accum_91__5_, prod_accum_91__4_, prod_accum_91__3_, prod_accum_91__2_, prod_accum_91__1_, prod_accum_91__0_ }),
    .a_o(a_r[11903:11776]),
    .b_o(b_r[11903:11776]),
    .s_o({ s_r_92__127_, s_r_92__126_, s_r_92__125_, s_r_92__124_, s_r_92__123_, s_r_92__122_, s_r_92__121_, s_r_92__120_, s_r_92__119_, s_r_92__118_, s_r_92__117_, s_r_92__116_, s_r_92__115_, s_r_92__114_, s_r_92__113_, s_r_92__112_, s_r_92__111_, s_r_92__110_, s_r_92__109_, s_r_92__108_, s_r_92__107_, s_r_92__106_, s_r_92__105_, s_r_92__104_, s_r_92__103_, s_r_92__102_, s_r_92__101_, s_r_92__100_, s_r_92__99_, s_r_92__98_, s_r_92__97_, s_r_92__96_, s_r_92__95_, s_r_92__94_, s_r_92__93_, s_r_92__92_, s_r_92__91_, s_r_92__90_, s_r_92__89_, s_r_92__88_, s_r_92__87_, s_r_92__86_, s_r_92__85_, s_r_92__84_, s_r_92__83_, s_r_92__82_, s_r_92__81_, s_r_92__80_, s_r_92__79_, s_r_92__78_, s_r_92__77_, s_r_92__76_, s_r_92__75_, s_r_92__74_, s_r_92__73_, s_r_92__72_, s_r_92__71_, s_r_92__70_, s_r_92__69_, s_r_92__68_, s_r_92__67_, s_r_92__66_, s_r_92__65_, s_r_92__64_, s_r_92__63_, s_r_92__62_, s_r_92__61_, s_r_92__60_, s_r_92__59_, s_r_92__58_, s_r_92__57_, s_r_92__56_, s_r_92__55_, s_r_92__54_, s_r_92__53_, s_r_92__52_, s_r_92__51_, s_r_92__50_, s_r_92__49_, s_r_92__48_, s_r_92__47_, s_r_92__46_, s_r_92__45_, s_r_92__44_, s_r_92__43_, s_r_92__42_, s_r_92__41_, s_r_92__40_, s_r_92__39_, s_r_92__38_, s_r_92__37_, s_r_92__36_, s_r_92__35_, s_r_92__34_, s_r_92__33_, s_r_92__32_, s_r_92__31_, s_r_92__30_, s_r_92__29_, s_r_92__28_, s_r_92__27_, s_r_92__26_, s_r_92__25_, s_r_92__24_, s_r_92__23_, s_r_92__22_, s_r_92__21_, s_r_92__20_, s_r_92__19_, s_r_92__18_, s_r_92__17_, s_r_92__16_, s_r_92__15_, s_r_92__14_, s_r_92__13_, s_r_92__12_, s_r_92__11_, s_r_92__10_, s_r_92__9_, s_r_92__8_, s_r_92__7_, s_r_92__6_, s_r_92__5_, s_r_92__4_, s_r_92__3_, s_r_92__2_, s_r_92__1_, s_r_92__0_ }),
    .c_o(c_r[92]),
    .prod_accum_o({ prod_accum_92__93_, prod_accum_92__92_, prod_accum_92__91_, prod_accum_92__90_, prod_accum_92__89_, prod_accum_92__88_, prod_accum_92__87_, prod_accum_92__86_, prod_accum_92__85_, prod_accum_92__84_, prod_accum_92__83_, prod_accum_92__82_, prod_accum_92__81_, prod_accum_92__80_, prod_accum_92__79_, prod_accum_92__78_, prod_accum_92__77_, prod_accum_92__76_, prod_accum_92__75_, prod_accum_92__74_, prod_accum_92__73_, prod_accum_92__72_, prod_accum_92__71_, prod_accum_92__70_, prod_accum_92__69_, prod_accum_92__68_, prod_accum_92__67_, prod_accum_92__66_, prod_accum_92__65_, prod_accum_92__64_, prod_accum_92__63_, prod_accum_92__62_, prod_accum_92__61_, prod_accum_92__60_, prod_accum_92__59_, prod_accum_92__58_, prod_accum_92__57_, prod_accum_92__56_, prod_accum_92__55_, prod_accum_92__54_, prod_accum_92__53_, prod_accum_92__52_, prod_accum_92__51_, prod_accum_92__50_, prod_accum_92__49_, prod_accum_92__48_, prod_accum_92__47_, prod_accum_92__46_, prod_accum_92__45_, prod_accum_92__44_, prod_accum_92__43_, prod_accum_92__42_, prod_accum_92__41_, prod_accum_92__40_, prod_accum_92__39_, prod_accum_92__38_, prod_accum_92__37_, prod_accum_92__36_, prod_accum_92__35_, prod_accum_92__34_, prod_accum_92__33_, prod_accum_92__32_, prod_accum_92__31_, prod_accum_92__30_, prod_accum_92__29_, prod_accum_92__28_, prod_accum_92__27_, prod_accum_92__26_, prod_accum_92__25_, prod_accum_92__24_, prod_accum_92__23_, prod_accum_92__22_, prod_accum_92__21_, prod_accum_92__20_, prod_accum_92__19_, prod_accum_92__18_, prod_accum_92__17_, prod_accum_92__16_, prod_accum_92__15_, prod_accum_92__14_, prod_accum_92__13_, prod_accum_92__12_, prod_accum_92__11_, prod_accum_92__10_, prod_accum_92__9_, prod_accum_92__8_, prod_accum_92__7_, prod_accum_92__6_, prod_accum_92__5_, prod_accum_92__4_, prod_accum_92__3_, prod_accum_92__2_, prod_accum_92__1_, prod_accum_92__0_ })
  );


  bsg_mul_array_row_128_93_x
  genblk1_93__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[11903:11776]),
    .b_i(b_r[11903:11776]),
    .s_i({ s_r_92__127_, s_r_92__126_, s_r_92__125_, s_r_92__124_, s_r_92__123_, s_r_92__122_, s_r_92__121_, s_r_92__120_, s_r_92__119_, s_r_92__118_, s_r_92__117_, s_r_92__116_, s_r_92__115_, s_r_92__114_, s_r_92__113_, s_r_92__112_, s_r_92__111_, s_r_92__110_, s_r_92__109_, s_r_92__108_, s_r_92__107_, s_r_92__106_, s_r_92__105_, s_r_92__104_, s_r_92__103_, s_r_92__102_, s_r_92__101_, s_r_92__100_, s_r_92__99_, s_r_92__98_, s_r_92__97_, s_r_92__96_, s_r_92__95_, s_r_92__94_, s_r_92__93_, s_r_92__92_, s_r_92__91_, s_r_92__90_, s_r_92__89_, s_r_92__88_, s_r_92__87_, s_r_92__86_, s_r_92__85_, s_r_92__84_, s_r_92__83_, s_r_92__82_, s_r_92__81_, s_r_92__80_, s_r_92__79_, s_r_92__78_, s_r_92__77_, s_r_92__76_, s_r_92__75_, s_r_92__74_, s_r_92__73_, s_r_92__72_, s_r_92__71_, s_r_92__70_, s_r_92__69_, s_r_92__68_, s_r_92__67_, s_r_92__66_, s_r_92__65_, s_r_92__64_, s_r_92__63_, s_r_92__62_, s_r_92__61_, s_r_92__60_, s_r_92__59_, s_r_92__58_, s_r_92__57_, s_r_92__56_, s_r_92__55_, s_r_92__54_, s_r_92__53_, s_r_92__52_, s_r_92__51_, s_r_92__50_, s_r_92__49_, s_r_92__48_, s_r_92__47_, s_r_92__46_, s_r_92__45_, s_r_92__44_, s_r_92__43_, s_r_92__42_, s_r_92__41_, s_r_92__40_, s_r_92__39_, s_r_92__38_, s_r_92__37_, s_r_92__36_, s_r_92__35_, s_r_92__34_, s_r_92__33_, s_r_92__32_, s_r_92__31_, s_r_92__30_, s_r_92__29_, s_r_92__28_, s_r_92__27_, s_r_92__26_, s_r_92__25_, s_r_92__24_, s_r_92__23_, s_r_92__22_, s_r_92__21_, s_r_92__20_, s_r_92__19_, s_r_92__18_, s_r_92__17_, s_r_92__16_, s_r_92__15_, s_r_92__14_, s_r_92__13_, s_r_92__12_, s_r_92__11_, s_r_92__10_, s_r_92__9_, s_r_92__8_, s_r_92__7_, s_r_92__6_, s_r_92__5_, s_r_92__4_, s_r_92__3_, s_r_92__2_, s_r_92__1_, s_r_92__0_ }),
    .c_i(c_r[92]),
    .prod_accum_i({ prod_accum_92__93_, prod_accum_92__92_, prod_accum_92__91_, prod_accum_92__90_, prod_accum_92__89_, prod_accum_92__88_, prod_accum_92__87_, prod_accum_92__86_, prod_accum_92__85_, prod_accum_92__84_, prod_accum_92__83_, prod_accum_92__82_, prod_accum_92__81_, prod_accum_92__80_, prod_accum_92__79_, prod_accum_92__78_, prod_accum_92__77_, prod_accum_92__76_, prod_accum_92__75_, prod_accum_92__74_, prod_accum_92__73_, prod_accum_92__72_, prod_accum_92__71_, prod_accum_92__70_, prod_accum_92__69_, prod_accum_92__68_, prod_accum_92__67_, prod_accum_92__66_, prod_accum_92__65_, prod_accum_92__64_, prod_accum_92__63_, prod_accum_92__62_, prod_accum_92__61_, prod_accum_92__60_, prod_accum_92__59_, prod_accum_92__58_, prod_accum_92__57_, prod_accum_92__56_, prod_accum_92__55_, prod_accum_92__54_, prod_accum_92__53_, prod_accum_92__52_, prod_accum_92__51_, prod_accum_92__50_, prod_accum_92__49_, prod_accum_92__48_, prod_accum_92__47_, prod_accum_92__46_, prod_accum_92__45_, prod_accum_92__44_, prod_accum_92__43_, prod_accum_92__42_, prod_accum_92__41_, prod_accum_92__40_, prod_accum_92__39_, prod_accum_92__38_, prod_accum_92__37_, prod_accum_92__36_, prod_accum_92__35_, prod_accum_92__34_, prod_accum_92__33_, prod_accum_92__32_, prod_accum_92__31_, prod_accum_92__30_, prod_accum_92__29_, prod_accum_92__28_, prod_accum_92__27_, prod_accum_92__26_, prod_accum_92__25_, prod_accum_92__24_, prod_accum_92__23_, prod_accum_92__22_, prod_accum_92__21_, prod_accum_92__20_, prod_accum_92__19_, prod_accum_92__18_, prod_accum_92__17_, prod_accum_92__16_, prod_accum_92__15_, prod_accum_92__14_, prod_accum_92__13_, prod_accum_92__12_, prod_accum_92__11_, prod_accum_92__10_, prod_accum_92__9_, prod_accum_92__8_, prod_accum_92__7_, prod_accum_92__6_, prod_accum_92__5_, prod_accum_92__4_, prod_accum_92__3_, prod_accum_92__2_, prod_accum_92__1_, prod_accum_92__0_ }),
    .a_o(a_r[12031:11904]),
    .b_o(b_r[12031:11904]),
    .s_o({ s_r_93__127_, s_r_93__126_, s_r_93__125_, s_r_93__124_, s_r_93__123_, s_r_93__122_, s_r_93__121_, s_r_93__120_, s_r_93__119_, s_r_93__118_, s_r_93__117_, s_r_93__116_, s_r_93__115_, s_r_93__114_, s_r_93__113_, s_r_93__112_, s_r_93__111_, s_r_93__110_, s_r_93__109_, s_r_93__108_, s_r_93__107_, s_r_93__106_, s_r_93__105_, s_r_93__104_, s_r_93__103_, s_r_93__102_, s_r_93__101_, s_r_93__100_, s_r_93__99_, s_r_93__98_, s_r_93__97_, s_r_93__96_, s_r_93__95_, s_r_93__94_, s_r_93__93_, s_r_93__92_, s_r_93__91_, s_r_93__90_, s_r_93__89_, s_r_93__88_, s_r_93__87_, s_r_93__86_, s_r_93__85_, s_r_93__84_, s_r_93__83_, s_r_93__82_, s_r_93__81_, s_r_93__80_, s_r_93__79_, s_r_93__78_, s_r_93__77_, s_r_93__76_, s_r_93__75_, s_r_93__74_, s_r_93__73_, s_r_93__72_, s_r_93__71_, s_r_93__70_, s_r_93__69_, s_r_93__68_, s_r_93__67_, s_r_93__66_, s_r_93__65_, s_r_93__64_, s_r_93__63_, s_r_93__62_, s_r_93__61_, s_r_93__60_, s_r_93__59_, s_r_93__58_, s_r_93__57_, s_r_93__56_, s_r_93__55_, s_r_93__54_, s_r_93__53_, s_r_93__52_, s_r_93__51_, s_r_93__50_, s_r_93__49_, s_r_93__48_, s_r_93__47_, s_r_93__46_, s_r_93__45_, s_r_93__44_, s_r_93__43_, s_r_93__42_, s_r_93__41_, s_r_93__40_, s_r_93__39_, s_r_93__38_, s_r_93__37_, s_r_93__36_, s_r_93__35_, s_r_93__34_, s_r_93__33_, s_r_93__32_, s_r_93__31_, s_r_93__30_, s_r_93__29_, s_r_93__28_, s_r_93__27_, s_r_93__26_, s_r_93__25_, s_r_93__24_, s_r_93__23_, s_r_93__22_, s_r_93__21_, s_r_93__20_, s_r_93__19_, s_r_93__18_, s_r_93__17_, s_r_93__16_, s_r_93__15_, s_r_93__14_, s_r_93__13_, s_r_93__12_, s_r_93__11_, s_r_93__10_, s_r_93__9_, s_r_93__8_, s_r_93__7_, s_r_93__6_, s_r_93__5_, s_r_93__4_, s_r_93__3_, s_r_93__2_, s_r_93__1_, s_r_93__0_ }),
    .c_o(c_r[93]),
    .prod_accum_o({ prod_accum_93__94_, prod_accum_93__93_, prod_accum_93__92_, prod_accum_93__91_, prod_accum_93__90_, prod_accum_93__89_, prod_accum_93__88_, prod_accum_93__87_, prod_accum_93__86_, prod_accum_93__85_, prod_accum_93__84_, prod_accum_93__83_, prod_accum_93__82_, prod_accum_93__81_, prod_accum_93__80_, prod_accum_93__79_, prod_accum_93__78_, prod_accum_93__77_, prod_accum_93__76_, prod_accum_93__75_, prod_accum_93__74_, prod_accum_93__73_, prod_accum_93__72_, prod_accum_93__71_, prod_accum_93__70_, prod_accum_93__69_, prod_accum_93__68_, prod_accum_93__67_, prod_accum_93__66_, prod_accum_93__65_, prod_accum_93__64_, prod_accum_93__63_, prod_accum_93__62_, prod_accum_93__61_, prod_accum_93__60_, prod_accum_93__59_, prod_accum_93__58_, prod_accum_93__57_, prod_accum_93__56_, prod_accum_93__55_, prod_accum_93__54_, prod_accum_93__53_, prod_accum_93__52_, prod_accum_93__51_, prod_accum_93__50_, prod_accum_93__49_, prod_accum_93__48_, prod_accum_93__47_, prod_accum_93__46_, prod_accum_93__45_, prod_accum_93__44_, prod_accum_93__43_, prod_accum_93__42_, prod_accum_93__41_, prod_accum_93__40_, prod_accum_93__39_, prod_accum_93__38_, prod_accum_93__37_, prod_accum_93__36_, prod_accum_93__35_, prod_accum_93__34_, prod_accum_93__33_, prod_accum_93__32_, prod_accum_93__31_, prod_accum_93__30_, prod_accum_93__29_, prod_accum_93__28_, prod_accum_93__27_, prod_accum_93__26_, prod_accum_93__25_, prod_accum_93__24_, prod_accum_93__23_, prod_accum_93__22_, prod_accum_93__21_, prod_accum_93__20_, prod_accum_93__19_, prod_accum_93__18_, prod_accum_93__17_, prod_accum_93__16_, prod_accum_93__15_, prod_accum_93__14_, prod_accum_93__13_, prod_accum_93__12_, prod_accum_93__11_, prod_accum_93__10_, prod_accum_93__9_, prod_accum_93__8_, prod_accum_93__7_, prod_accum_93__6_, prod_accum_93__5_, prod_accum_93__4_, prod_accum_93__3_, prod_accum_93__2_, prod_accum_93__1_, prod_accum_93__0_ })
  );


  bsg_mul_array_row_128_94_x
  genblk1_94__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[12031:11904]),
    .b_i(b_r[12031:11904]),
    .s_i({ s_r_93__127_, s_r_93__126_, s_r_93__125_, s_r_93__124_, s_r_93__123_, s_r_93__122_, s_r_93__121_, s_r_93__120_, s_r_93__119_, s_r_93__118_, s_r_93__117_, s_r_93__116_, s_r_93__115_, s_r_93__114_, s_r_93__113_, s_r_93__112_, s_r_93__111_, s_r_93__110_, s_r_93__109_, s_r_93__108_, s_r_93__107_, s_r_93__106_, s_r_93__105_, s_r_93__104_, s_r_93__103_, s_r_93__102_, s_r_93__101_, s_r_93__100_, s_r_93__99_, s_r_93__98_, s_r_93__97_, s_r_93__96_, s_r_93__95_, s_r_93__94_, s_r_93__93_, s_r_93__92_, s_r_93__91_, s_r_93__90_, s_r_93__89_, s_r_93__88_, s_r_93__87_, s_r_93__86_, s_r_93__85_, s_r_93__84_, s_r_93__83_, s_r_93__82_, s_r_93__81_, s_r_93__80_, s_r_93__79_, s_r_93__78_, s_r_93__77_, s_r_93__76_, s_r_93__75_, s_r_93__74_, s_r_93__73_, s_r_93__72_, s_r_93__71_, s_r_93__70_, s_r_93__69_, s_r_93__68_, s_r_93__67_, s_r_93__66_, s_r_93__65_, s_r_93__64_, s_r_93__63_, s_r_93__62_, s_r_93__61_, s_r_93__60_, s_r_93__59_, s_r_93__58_, s_r_93__57_, s_r_93__56_, s_r_93__55_, s_r_93__54_, s_r_93__53_, s_r_93__52_, s_r_93__51_, s_r_93__50_, s_r_93__49_, s_r_93__48_, s_r_93__47_, s_r_93__46_, s_r_93__45_, s_r_93__44_, s_r_93__43_, s_r_93__42_, s_r_93__41_, s_r_93__40_, s_r_93__39_, s_r_93__38_, s_r_93__37_, s_r_93__36_, s_r_93__35_, s_r_93__34_, s_r_93__33_, s_r_93__32_, s_r_93__31_, s_r_93__30_, s_r_93__29_, s_r_93__28_, s_r_93__27_, s_r_93__26_, s_r_93__25_, s_r_93__24_, s_r_93__23_, s_r_93__22_, s_r_93__21_, s_r_93__20_, s_r_93__19_, s_r_93__18_, s_r_93__17_, s_r_93__16_, s_r_93__15_, s_r_93__14_, s_r_93__13_, s_r_93__12_, s_r_93__11_, s_r_93__10_, s_r_93__9_, s_r_93__8_, s_r_93__7_, s_r_93__6_, s_r_93__5_, s_r_93__4_, s_r_93__3_, s_r_93__2_, s_r_93__1_, s_r_93__0_ }),
    .c_i(c_r[93]),
    .prod_accum_i({ prod_accum_93__94_, prod_accum_93__93_, prod_accum_93__92_, prod_accum_93__91_, prod_accum_93__90_, prod_accum_93__89_, prod_accum_93__88_, prod_accum_93__87_, prod_accum_93__86_, prod_accum_93__85_, prod_accum_93__84_, prod_accum_93__83_, prod_accum_93__82_, prod_accum_93__81_, prod_accum_93__80_, prod_accum_93__79_, prod_accum_93__78_, prod_accum_93__77_, prod_accum_93__76_, prod_accum_93__75_, prod_accum_93__74_, prod_accum_93__73_, prod_accum_93__72_, prod_accum_93__71_, prod_accum_93__70_, prod_accum_93__69_, prod_accum_93__68_, prod_accum_93__67_, prod_accum_93__66_, prod_accum_93__65_, prod_accum_93__64_, prod_accum_93__63_, prod_accum_93__62_, prod_accum_93__61_, prod_accum_93__60_, prod_accum_93__59_, prod_accum_93__58_, prod_accum_93__57_, prod_accum_93__56_, prod_accum_93__55_, prod_accum_93__54_, prod_accum_93__53_, prod_accum_93__52_, prod_accum_93__51_, prod_accum_93__50_, prod_accum_93__49_, prod_accum_93__48_, prod_accum_93__47_, prod_accum_93__46_, prod_accum_93__45_, prod_accum_93__44_, prod_accum_93__43_, prod_accum_93__42_, prod_accum_93__41_, prod_accum_93__40_, prod_accum_93__39_, prod_accum_93__38_, prod_accum_93__37_, prod_accum_93__36_, prod_accum_93__35_, prod_accum_93__34_, prod_accum_93__33_, prod_accum_93__32_, prod_accum_93__31_, prod_accum_93__30_, prod_accum_93__29_, prod_accum_93__28_, prod_accum_93__27_, prod_accum_93__26_, prod_accum_93__25_, prod_accum_93__24_, prod_accum_93__23_, prod_accum_93__22_, prod_accum_93__21_, prod_accum_93__20_, prod_accum_93__19_, prod_accum_93__18_, prod_accum_93__17_, prod_accum_93__16_, prod_accum_93__15_, prod_accum_93__14_, prod_accum_93__13_, prod_accum_93__12_, prod_accum_93__11_, prod_accum_93__10_, prod_accum_93__9_, prod_accum_93__8_, prod_accum_93__7_, prod_accum_93__6_, prod_accum_93__5_, prod_accum_93__4_, prod_accum_93__3_, prod_accum_93__2_, prod_accum_93__1_, prod_accum_93__0_ }),
    .a_o(a_r[12159:12032]),
    .b_o(b_r[12159:12032]),
    .s_o({ s_r_94__127_, s_r_94__126_, s_r_94__125_, s_r_94__124_, s_r_94__123_, s_r_94__122_, s_r_94__121_, s_r_94__120_, s_r_94__119_, s_r_94__118_, s_r_94__117_, s_r_94__116_, s_r_94__115_, s_r_94__114_, s_r_94__113_, s_r_94__112_, s_r_94__111_, s_r_94__110_, s_r_94__109_, s_r_94__108_, s_r_94__107_, s_r_94__106_, s_r_94__105_, s_r_94__104_, s_r_94__103_, s_r_94__102_, s_r_94__101_, s_r_94__100_, s_r_94__99_, s_r_94__98_, s_r_94__97_, s_r_94__96_, s_r_94__95_, s_r_94__94_, s_r_94__93_, s_r_94__92_, s_r_94__91_, s_r_94__90_, s_r_94__89_, s_r_94__88_, s_r_94__87_, s_r_94__86_, s_r_94__85_, s_r_94__84_, s_r_94__83_, s_r_94__82_, s_r_94__81_, s_r_94__80_, s_r_94__79_, s_r_94__78_, s_r_94__77_, s_r_94__76_, s_r_94__75_, s_r_94__74_, s_r_94__73_, s_r_94__72_, s_r_94__71_, s_r_94__70_, s_r_94__69_, s_r_94__68_, s_r_94__67_, s_r_94__66_, s_r_94__65_, s_r_94__64_, s_r_94__63_, s_r_94__62_, s_r_94__61_, s_r_94__60_, s_r_94__59_, s_r_94__58_, s_r_94__57_, s_r_94__56_, s_r_94__55_, s_r_94__54_, s_r_94__53_, s_r_94__52_, s_r_94__51_, s_r_94__50_, s_r_94__49_, s_r_94__48_, s_r_94__47_, s_r_94__46_, s_r_94__45_, s_r_94__44_, s_r_94__43_, s_r_94__42_, s_r_94__41_, s_r_94__40_, s_r_94__39_, s_r_94__38_, s_r_94__37_, s_r_94__36_, s_r_94__35_, s_r_94__34_, s_r_94__33_, s_r_94__32_, s_r_94__31_, s_r_94__30_, s_r_94__29_, s_r_94__28_, s_r_94__27_, s_r_94__26_, s_r_94__25_, s_r_94__24_, s_r_94__23_, s_r_94__22_, s_r_94__21_, s_r_94__20_, s_r_94__19_, s_r_94__18_, s_r_94__17_, s_r_94__16_, s_r_94__15_, s_r_94__14_, s_r_94__13_, s_r_94__12_, s_r_94__11_, s_r_94__10_, s_r_94__9_, s_r_94__8_, s_r_94__7_, s_r_94__6_, s_r_94__5_, s_r_94__4_, s_r_94__3_, s_r_94__2_, s_r_94__1_, s_r_94__0_ }),
    .c_o(c_r[94]),
    .prod_accum_o({ prod_accum_94__95_, prod_accum_94__94_, prod_accum_94__93_, prod_accum_94__92_, prod_accum_94__91_, prod_accum_94__90_, prod_accum_94__89_, prod_accum_94__88_, prod_accum_94__87_, prod_accum_94__86_, prod_accum_94__85_, prod_accum_94__84_, prod_accum_94__83_, prod_accum_94__82_, prod_accum_94__81_, prod_accum_94__80_, prod_accum_94__79_, prod_accum_94__78_, prod_accum_94__77_, prod_accum_94__76_, prod_accum_94__75_, prod_accum_94__74_, prod_accum_94__73_, prod_accum_94__72_, prod_accum_94__71_, prod_accum_94__70_, prod_accum_94__69_, prod_accum_94__68_, prod_accum_94__67_, prod_accum_94__66_, prod_accum_94__65_, prod_accum_94__64_, prod_accum_94__63_, prod_accum_94__62_, prod_accum_94__61_, prod_accum_94__60_, prod_accum_94__59_, prod_accum_94__58_, prod_accum_94__57_, prod_accum_94__56_, prod_accum_94__55_, prod_accum_94__54_, prod_accum_94__53_, prod_accum_94__52_, prod_accum_94__51_, prod_accum_94__50_, prod_accum_94__49_, prod_accum_94__48_, prod_accum_94__47_, prod_accum_94__46_, prod_accum_94__45_, prod_accum_94__44_, prod_accum_94__43_, prod_accum_94__42_, prod_accum_94__41_, prod_accum_94__40_, prod_accum_94__39_, prod_accum_94__38_, prod_accum_94__37_, prod_accum_94__36_, prod_accum_94__35_, prod_accum_94__34_, prod_accum_94__33_, prod_accum_94__32_, prod_accum_94__31_, prod_accum_94__30_, prod_accum_94__29_, prod_accum_94__28_, prod_accum_94__27_, prod_accum_94__26_, prod_accum_94__25_, prod_accum_94__24_, prod_accum_94__23_, prod_accum_94__22_, prod_accum_94__21_, prod_accum_94__20_, prod_accum_94__19_, prod_accum_94__18_, prod_accum_94__17_, prod_accum_94__16_, prod_accum_94__15_, prod_accum_94__14_, prod_accum_94__13_, prod_accum_94__12_, prod_accum_94__11_, prod_accum_94__10_, prod_accum_94__9_, prod_accum_94__8_, prod_accum_94__7_, prod_accum_94__6_, prod_accum_94__5_, prod_accum_94__4_, prod_accum_94__3_, prod_accum_94__2_, prod_accum_94__1_, prod_accum_94__0_ })
  );


  bsg_mul_array_row_128_95_x
  genblk1_95__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[12159:12032]),
    .b_i(b_r[12159:12032]),
    .s_i({ s_r_94__127_, s_r_94__126_, s_r_94__125_, s_r_94__124_, s_r_94__123_, s_r_94__122_, s_r_94__121_, s_r_94__120_, s_r_94__119_, s_r_94__118_, s_r_94__117_, s_r_94__116_, s_r_94__115_, s_r_94__114_, s_r_94__113_, s_r_94__112_, s_r_94__111_, s_r_94__110_, s_r_94__109_, s_r_94__108_, s_r_94__107_, s_r_94__106_, s_r_94__105_, s_r_94__104_, s_r_94__103_, s_r_94__102_, s_r_94__101_, s_r_94__100_, s_r_94__99_, s_r_94__98_, s_r_94__97_, s_r_94__96_, s_r_94__95_, s_r_94__94_, s_r_94__93_, s_r_94__92_, s_r_94__91_, s_r_94__90_, s_r_94__89_, s_r_94__88_, s_r_94__87_, s_r_94__86_, s_r_94__85_, s_r_94__84_, s_r_94__83_, s_r_94__82_, s_r_94__81_, s_r_94__80_, s_r_94__79_, s_r_94__78_, s_r_94__77_, s_r_94__76_, s_r_94__75_, s_r_94__74_, s_r_94__73_, s_r_94__72_, s_r_94__71_, s_r_94__70_, s_r_94__69_, s_r_94__68_, s_r_94__67_, s_r_94__66_, s_r_94__65_, s_r_94__64_, s_r_94__63_, s_r_94__62_, s_r_94__61_, s_r_94__60_, s_r_94__59_, s_r_94__58_, s_r_94__57_, s_r_94__56_, s_r_94__55_, s_r_94__54_, s_r_94__53_, s_r_94__52_, s_r_94__51_, s_r_94__50_, s_r_94__49_, s_r_94__48_, s_r_94__47_, s_r_94__46_, s_r_94__45_, s_r_94__44_, s_r_94__43_, s_r_94__42_, s_r_94__41_, s_r_94__40_, s_r_94__39_, s_r_94__38_, s_r_94__37_, s_r_94__36_, s_r_94__35_, s_r_94__34_, s_r_94__33_, s_r_94__32_, s_r_94__31_, s_r_94__30_, s_r_94__29_, s_r_94__28_, s_r_94__27_, s_r_94__26_, s_r_94__25_, s_r_94__24_, s_r_94__23_, s_r_94__22_, s_r_94__21_, s_r_94__20_, s_r_94__19_, s_r_94__18_, s_r_94__17_, s_r_94__16_, s_r_94__15_, s_r_94__14_, s_r_94__13_, s_r_94__12_, s_r_94__11_, s_r_94__10_, s_r_94__9_, s_r_94__8_, s_r_94__7_, s_r_94__6_, s_r_94__5_, s_r_94__4_, s_r_94__3_, s_r_94__2_, s_r_94__1_, s_r_94__0_ }),
    .c_i(c_r[94]),
    .prod_accum_i({ prod_accum_94__95_, prod_accum_94__94_, prod_accum_94__93_, prod_accum_94__92_, prod_accum_94__91_, prod_accum_94__90_, prod_accum_94__89_, prod_accum_94__88_, prod_accum_94__87_, prod_accum_94__86_, prod_accum_94__85_, prod_accum_94__84_, prod_accum_94__83_, prod_accum_94__82_, prod_accum_94__81_, prod_accum_94__80_, prod_accum_94__79_, prod_accum_94__78_, prod_accum_94__77_, prod_accum_94__76_, prod_accum_94__75_, prod_accum_94__74_, prod_accum_94__73_, prod_accum_94__72_, prod_accum_94__71_, prod_accum_94__70_, prod_accum_94__69_, prod_accum_94__68_, prod_accum_94__67_, prod_accum_94__66_, prod_accum_94__65_, prod_accum_94__64_, prod_accum_94__63_, prod_accum_94__62_, prod_accum_94__61_, prod_accum_94__60_, prod_accum_94__59_, prod_accum_94__58_, prod_accum_94__57_, prod_accum_94__56_, prod_accum_94__55_, prod_accum_94__54_, prod_accum_94__53_, prod_accum_94__52_, prod_accum_94__51_, prod_accum_94__50_, prod_accum_94__49_, prod_accum_94__48_, prod_accum_94__47_, prod_accum_94__46_, prod_accum_94__45_, prod_accum_94__44_, prod_accum_94__43_, prod_accum_94__42_, prod_accum_94__41_, prod_accum_94__40_, prod_accum_94__39_, prod_accum_94__38_, prod_accum_94__37_, prod_accum_94__36_, prod_accum_94__35_, prod_accum_94__34_, prod_accum_94__33_, prod_accum_94__32_, prod_accum_94__31_, prod_accum_94__30_, prod_accum_94__29_, prod_accum_94__28_, prod_accum_94__27_, prod_accum_94__26_, prod_accum_94__25_, prod_accum_94__24_, prod_accum_94__23_, prod_accum_94__22_, prod_accum_94__21_, prod_accum_94__20_, prod_accum_94__19_, prod_accum_94__18_, prod_accum_94__17_, prod_accum_94__16_, prod_accum_94__15_, prod_accum_94__14_, prod_accum_94__13_, prod_accum_94__12_, prod_accum_94__11_, prod_accum_94__10_, prod_accum_94__9_, prod_accum_94__8_, prod_accum_94__7_, prod_accum_94__6_, prod_accum_94__5_, prod_accum_94__4_, prod_accum_94__3_, prod_accum_94__2_, prod_accum_94__1_, prod_accum_94__0_ }),
    .a_o(a_r[12287:12160]),
    .b_o(b_r[12287:12160]),
    .s_o({ s_r_95__127_, s_r_95__126_, s_r_95__125_, s_r_95__124_, s_r_95__123_, s_r_95__122_, s_r_95__121_, s_r_95__120_, s_r_95__119_, s_r_95__118_, s_r_95__117_, s_r_95__116_, s_r_95__115_, s_r_95__114_, s_r_95__113_, s_r_95__112_, s_r_95__111_, s_r_95__110_, s_r_95__109_, s_r_95__108_, s_r_95__107_, s_r_95__106_, s_r_95__105_, s_r_95__104_, s_r_95__103_, s_r_95__102_, s_r_95__101_, s_r_95__100_, s_r_95__99_, s_r_95__98_, s_r_95__97_, s_r_95__96_, s_r_95__95_, s_r_95__94_, s_r_95__93_, s_r_95__92_, s_r_95__91_, s_r_95__90_, s_r_95__89_, s_r_95__88_, s_r_95__87_, s_r_95__86_, s_r_95__85_, s_r_95__84_, s_r_95__83_, s_r_95__82_, s_r_95__81_, s_r_95__80_, s_r_95__79_, s_r_95__78_, s_r_95__77_, s_r_95__76_, s_r_95__75_, s_r_95__74_, s_r_95__73_, s_r_95__72_, s_r_95__71_, s_r_95__70_, s_r_95__69_, s_r_95__68_, s_r_95__67_, s_r_95__66_, s_r_95__65_, s_r_95__64_, s_r_95__63_, s_r_95__62_, s_r_95__61_, s_r_95__60_, s_r_95__59_, s_r_95__58_, s_r_95__57_, s_r_95__56_, s_r_95__55_, s_r_95__54_, s_r_95__53_, s_r_95__52_, s_r_95__51_, s_r_95__50_, s_r_95__49_, s_r_95__48_, s_r_95__47_, s_r_95__46_, s_r_95__45_, s_r_95__44_, s_r_95__43_, s_r_95__42_, s_r_95__41_, s_r_95__40_, s_r_95__39_, s_r_95__38_, s_r_95__37_, s_r_95__36_, s_r_95__35_, s_r_95__34_, s_r_95__33_, s_r_95__32_, s_r_95__31_, s_r_95__30_, s_r_95__29_, s_r_95__28_, s_r_95__27_, s_r_95__26_, s_r_95__25_, s_r_95__24_, s_r_95__23_, s_r_95__22_, s_r_95__21_, s_r_95__20_, s_r_95__19_, s_r_95__18_, s_r_95__17_, s_r_95__16_, s_r_95__15_, s_r_95__14_, s_r_95__13_, s_r_95__12_, s_r_95__11_, s_r_95__10_, s_r_95__9_, s_r_95__8_, s_r_95__7_, s_r_95__6_, s_r_95__5_, s_r_95__4_, s_r_95__3_, s_r_95__2_, s_r_95__1_, s_r_95__0_ }),
    .c_o(c_r[95]),
    .prod_accum_o({ prod_accum_95__96_, prod_accum_95__95_, prod_accum_95__94_, prod_accum_95__93_, prod_accum_95__92_, prod_accum_95__91_, prod_accum_95__90_, prod_accum_95__89_, prod_accum_95__88_, prod_accum_95__87_, prod_accum_95__86_, prod_accum_95__85_, prod_accum_95__84_, prod_accum_95__83_, prod_accum_95__82_, prod_accum_95__81_, prod_accum_95__80_, prod_accum_95__79_, prod_accum_95__78_, prod_accum_95__77_, prod_accum_95__76_, prod_accum_95__75_, prod_accum_95__74_, prod_accum_95__73_, prod_accum_95__72_, prod_accum_95__71_, prod_accum_95__70_, prod_accum_95__69_, prod_accum_95__68_, prod_accum_95__67_, prod_accum_95__66_, prod_accum_95__65_, prod_accum_95__64_, prod_accum_95__63_, prod_accum_95__62_, prod_accum_95__61_, prod_accum_95__60_, prod_accum_95__59_, prod_accum_95__58_, prod_accum_95__57_, prod_accum_95__56_, prod_accum_95__55_, prod_accum_95__54_, prod_accum_95__53_, prod_accum_95__52_, prod_accum_95__51_, prod_accum_95__50_, prod_accum_95__49_, prod_accum_95__48_, prod_accum_95__47_, prod_accum_95__46_, prod_accum_95__45_, prod_accum_95__44_, prod_accum_95__43_, prod_accum_95__42_, prod_accum_95__41_, prod_accum_95__40_, prod_accum_95__39_, prod_accum_95__38_, prod_accum_95__37_, prod_accum_95__36_, prod_accum_95__35_, prod_accum_95__34_, prod_accum_95__33_, prod_accum_95__32_, prod_accum_95__31_, prod_accum_95__30_, prod_accum_95__29_, prod_accum_95__28_, prod_accum_95__27_, prod_accum_95__26_, prod_accum_95__25_, prod_accum_95__24_, prod_accum_95__23_, prod_accum_95__22_, prod_accum_95__21_, prod_accum_95__20_, prod_accum_95__19_, prod_accum_95__18_, prod_accum_95__17_, prod_accum_95__16_, prod_accum_95__15_, prod_accum_95__14_, prod_accum_95__13_, prod_accum_95__12_, prod_accum_95__11_, prod_accum_95__10_, prod_accum_95__9_, prod_accum_95__8_, prod_accum_95__7_, prod_accum_95__6_, prod_accum_95__5_, prod_accum_95__4_, prod_accum_95__3_, prod_accum_95__2_, prod_accum_95__1_, prod_accum_95__0_ })
  );


  bsg_mul_array_row_128_96_x
  genblk1_96__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[12287:12160]),
    .b_i(b_r[12287:12160]),
    .s_i({ s_r_95__127_, s_r_95__126_, s_r_95__125_, s_r_95__124_, s_r_95__123_, s_r_95__122_, s_r_95__121_, s_r_95__120_, s_r_95__119_, s_r_95__118_, s_r_95__117_, s_r_95__116_, s_r_95__115_, s_r_95__114_, s_r_95__113_, s_r_95__112_, s_r_95__111_, s_r_95__110_, s_r_95__109_, s_r_95__108_, s_r_95__107_, s_r_95__106_, s_r_95__105_, s_r_95__104_, s_r_95__103_, s_r_95__102_, s_r_95__101_, s_r_95__100_, s_r_95__99_, s_r_95__98_, s_r_95__97_, s_r_95__96_, s_r_95__95_, s_r_95__94_, s_r_95__93_, s_r_95__92_, s_r_95__91_, s_r_95__90_, s_r_95__89_, s_r_95__88_, s_r_95__87_, s_r_95__86_, s_r_95__85_, s_r_95__84_, s_r_95__83_, s_r_95__82_, s_r_95__81_, s_r_95__80_, s_r_95__79_, s_r_95__78_, s_r_95__77_, s_r_95__76_, s_r_95__75_, s_r_95__74_, s_r_95__73_, s_r_95__72_, s_r_95__71_, s_r_95__70_, s_r_95__69_, s_r_95__68_, s_r_95__67_, s_r_95__66_, s_r_95__65_, s_r_95__64_, s_r_95__63_, s_r_95__62_, s_r_95__61_, s_r_95__60_, s_r_95__59_, s_r_95__58_, s_r_95__57_, s_r_95__56_, s_r_95__55_, s_r_95__54_, s_r_95__53_, s_r_95__52_, s_r_95__51_, s_r_95__50_, s_r_95__49_, s_r_95__48_, s_r_95__47_, s_r_95__46_, s_r_95__45_, s_r_95__44_, s_r_95__43_, s_r_95__42_, s_r_95__41_, s_r_95__40_, s_r_95__39_, s_r_95__38_, s_r_95__37_, s_r_95__36_, s_r_95__35_, s_r_95__34_, s_r_95__33_, s_r_95__32_, s_r_95__31_, s_r_95__30_, s_r_95__29_, s_r_95__28_, s_r_95__27_, s_r_95__26_, s_r_95__25_, s_r_95__24_, s_r_95__23_, s_r_95__22_, s_r_95__21_, s_r_95__20_, s_r_95__19_, s_r_95__18_, s_r_95__17_, s_r_95__16_, s_r_95__15_, s_r_95__14_, s_r_95__13_, s_r_95__12_, s_r_95__11_, s_r_95__10_, s_r_95__9_, s_r_95__8_, s_r_95__7_, s_r_95__6_, s_r_95__5_, s_r_95__4_, s_r_95__3_, s_r_95__2_, s_r_95__1_, s_r_95__0_ }),
    .c_i(c_r[95]),
    .prod_accum_i({ prod_accum_95__96_, prod_accum_95__95_, prod_accum_95__94_, prod_accum_95__93_, prod_accum_95__92_, prod_accum_95__91_, prod_accum_95__90_, prod_accum_95__89_, prod_accum_95__88_, prod_accum_95__87_, prod_accum_95__86_, prod_accum_95__85_, prod_accum_95__84_, prod_accum_95__83_, prod_accum_95__82_, prod_accum_95__81_, prod_accum_95__80_, prod_accum_95__79_, prod_accum_95__78_, prod_accum_95__77_, prod_accum_95__76_, prod_accum_95__75_, prod_accum_95__74_, prod_accum_95__73_, prod_accum_95__72_, prod_accum_95__71_, prod_accum_95__70_, prod_accum_95__69_, prod_accum_95__68_, prod_accum_95__67_, prod_accum_95__66_, prod_accum_95__65_, prod_accum_95__64_, prod_accum_95__63_, prod_accum_95__62_, prod_accum_95__61_, prod_accum_95__60_, prod_accum_95__59_, prod_accum_95__58_, prod_accum_95__57_, prod_accum_95__56_, prod_accum_95__55_, prod_accum_95__54_, prod_accum_95__53_, prod_accum_95__52_, prod_accum_95__51_, prod_accum_95__50_, prod_accum_95__49_, prod_accum_95__48_, prod_accum_95__47_, prod_accum_95__46_, prod_accum_95__45_, prod_accum_95__44_, prod_accum_95__43_, prod_accum_95__42_, prod_accum_95__41_, prod_accum_95__40_, prod_accum_95__39_, prod_accum_95__38_, prod_accum_95__37_, prod_accum_95__36_, prod_accum_95__35_, prod_accum_95__34_, prod_accum_95__33_, prod_accum_95__32_, prod_accum_95__31_, prod_accum_95__30_, prod_accum_95__29_, prod_accum_95__28_, prod_accum_95__27_, prod_accum_95__26_, prod_accum_95__25_, prod_accum_95__24_, prod_accum_95__23_, prod_accum_95__22_, prod_accum_95__21_, prod_accum_95__20_, prod_accum_95__19_, prod_accum_95__18_, prod_accum_95__17_, prod_accum_95__16_, prod_accum_95__15_, prod_accum_95__14_, prod_accum_95__13_, prod_accum_95__12_, prod_accum_95__11_, prod_accum_95__10_, prod_accum_95__9_, prod_accum_95__8_, prod_accum_95__7_, prod_accum_95__6_, prod_accum_95__5_, prod_accum_95__4_, prod_accum_95__3_, prod_accum_95__2_, prod_accum_95__1_, prod_accum_95__0_ }),
    .a_o(a_r[12415:12288]),
    .b_o(b_r[12415:12288]),
    .s_o({ s_r_96__127_, s_r_96__126_, s_r_96__125_, s_r_96__124_, s_r_96__123_, s_r_96__122_, s_r_96__121_, s_r_96__120_, s_r_96__119_, s_r_96__118_, s_r_96__117_, s_r_96__116_, s_r_96__115_, s_r_96__114_, s_r_96__113_, s_r_96__112_, s_r_96__111_, s_r_96__110_, s_r_96__109_, s_r_96__108_, s_r_96__107_, s_r_96__106_, s_r_96__105_, s_r_96__104_, s_r_96__103_, s_r_96__102_, s_r_96__101_, s_r_96__100_, s_r_96__99_, s_r_96__98_, s_r_96__97_, s_r_96__96_, s_r_96__95_, s_r_96__94_, s_r_96__93_, s_r_96__92_, s_r_96__91_, s_r_96__90_, s_r_96__89_, s_r_96__88_, s_r_96__87_, s_r_96__86_, s_r_96__85_, s_r_96__84_, s_r_96__83_, s_r_96__82_, s_r_96__81_, s_r_96__80_, s_r_96__79_, s_r_96__78_, s_r_96__77_, s_r_96__76_, s_r_96__75_, s_r_96__74_, s_r_96__73_, s_r_96__72_, s_r_96__71_, s_r_96__70_, s_r_96__69_, s_r_96__68_, s_r_96__67_, s_r_96__66_, s_r_96__65_, s_r_96__64_, s_r_96__63_, s_r_96__62_, s_r_96__61_, s_r_96__60_, s_r_96__59_, s_r_96__58_, s_r_96__57_, s_r_96__56_, s_r_96__55_, s_r_96__54_, s_r_96__53_, s_r_96__52_, s_r_96__51_, s_r_96__50_, s_r_96__49_, s_r_96__48_, s_r_96__47_, s_r_96__46_, s_r_96__45_, s_r_96__44_, s_r_96__43_, s_r_96__42_, s_r_96__41_, s_r_96__40_, s_r_96__39_, s_r_96__38_, s_r_96__37_, s_r_96__36_, s_r_96__35_, s_r_96__34_, s_r_96__33_, s_r_96__32_, s_r_96__31_, s_r_96__30_, s_r_96__29_, s_r_96__28_, s_r_96__27_, s_r_96__26_, s_r_96__25_, s_r_96__24_, s_r_96__23_, s_r_96__22_, s_r_96__21_, s_r_96__20_, s_r_96__19_, s_r_96__18_, s_r_96__17_, s_r_96__16_, s_r_96__15_, s_r_96__14_, s_r_96__13_, s_r_96__12_, s_r_96__11_, s_r_96__10_, s_r_96__9_, s_r_96__8_, s_r_96__7_, s_r_96__6_, s_r_96__5_, s_r_96__4_, s_r_96__3_, s_r_96__2_, s_r_96__1_, s_r_96__0_ }),
    .c_o(c_r[96]),
    .prod_accum_o({ prod_accum_96__97_, prod_accum_96__96_, prod_accum_96__95_, prod_accum_96__94_, prod_accum_96__93_, prod_accum_96__92_, prod_accum_96__91_, prod_accum_96__90_, prod_accum_96__89_, prod_accum_96__88_, prod_accum_96__87_, prod_accum_96__86_, prod_accum_96__85_, prod_accum_96__84_, prod_accum_96__83_, prod_accum_96__82_, prod_accum_96__81_, prod_accum_96__80_, prod_accum_96__79_, prod_accum_96__78_, prod_accum_96__77_, prod_accum_96__76_, prod_accum_96__75_, prod_accum_96__74_, prod_accum_96__73_, prod_accum_96__72_, prod_accum_96__71_, prod_accum_96__70_, prod_accum_96__69_, prod_accum_96__68_, prod_accum_96__67_, prod_accum_96__66_, prod_accum_96__65_, prod_accum_96__64_, prod_accum_96__63_, prod_accum_96__62_, prod_accum_96__61_, prod_accum_96__60_, prod_accum_96__59_, prod_accum_96__58_, prod_accum_96__57_, prod_accum_96__56_, prod_accum_96__55_, prod_accum_96__54_, prod_accum_96__53_, prod_accum_96__52_, prod_accum_96__51_, prod_accum_96__50_, prod_accum_96__49_, prod_accum_96__48_, prod_accum_96__47_, prod_accum_96__46_, prod_accum_96__45_, prod_accum_96__44_, prod_accum_96__43_, prod_accum_96__42_, prod_accum_96__41_, prod_accum_96__40_, prod_accum_96__39_, prod_accum_96__38_, prod_accum_96__37_, prod_accum_96__36_, prod_accum_96__35_, prod_accum_96__34_, prod_accum_96__33_, prod_accum_96__32_, prod_accum_96__31_, prod_accum_96__30_, prod_accum_96__29_, prod_accum_96__28_, prod_accum_96__27_, prod_accum_96__26_, prod_accum_96__25_, prod_accum_96__24_, prod_accum_96__23_, prod_accum_96__22_, prod_accum_96__21_, prod_accum_96__20_, prod_accum_96__19_, prod_accum_96__18_, prod_accum_96__17_, prod_accum_96__16_, prod_accum_96__15_, prod_accum_96__14_, prod_accum_96__13_, prod_accum_96__12_, prod_accum_96__11_, prod_accum_96__10_, prod_accum_96__9_, prod_accum_96__8_, prod_accum_96__7_, prod_accum_96__6_, prod_accum_96__5_, prod_accum_96__4_, prod_accum_96__3_, prod_accum_96__2_, prod_accum_96__1_, prod_accum_96__0_ })
  );


  bsg_mul_array_row_128_97_x
  genblk1_97__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[12415:12288]),
    .b_i(b_r[12415:12288]),
    .s_i({ s_r_96__127_, s_r_96__126_, s_r_96__125_, s_r_96__124_, s_r_96__123_, s_r_96__122_, s_r_96__121_, s_r_96__120_, s_r_96__119_, s_r_96__118_, s_r_96__117_, s_r_96__116_, s_r_96__115_, s_r_96__114_, s_r_96__113_, s_r_96__112_, s_r_96__111_, s_r_96__110_, s_r_96__109_, s_r_96__108_, s_r_96__107_, s_r_96__106_, s_r_96__105_, s_r_96__104_, s_r_96__103_, s_r_96__102_, s_r_96__101_, s_r_96__100_, s_r_96__99_, s_r_96__98_, s_r_96__97_, s_r_96__96_, s_r_96__95_, s_r_96__94_, s_r_96__93_, s_r_96__92_, s_r_96__91_, s_r_96__90_, s_r_96__89_, s_r_96__88_, s_r_96__87_, s_r_96__86_, s_r_96__85_, s_r_96__84_, s_r_96__83_, s_r_96__82_, s_r_96__81_, s_r_96__80_, s_r_96__79_, s_r_96__78_, s_r_96__77_, s_r_96__76_, s_r_96__75_, s_r_96__74_, s_r_96__73_, s_r_96__72_, s_r_96__71_, s_r_96__70_, s_r_96__69_, s_r_96__68_, s_r_96__67_, s_r_96__66_, s_r_96__65_, s_r_96__64_, s_r_96__63_, s_r_96__62_, s_r_96__61_, s_r_96__60_, s_r_96__59_, s_r_96__58_, s_r_96__57_, s_r_96__56_, s_r_96__55_, s_r_96__54_, s_r_96__53_, s_r_96__52_, s_r_96__51_, s_r_96__50_, s_r_96__49_, s_r_96__48_, s_r_96__47_, s_r_96__46_, s_r_96__45_, s_r_96__44_, s_r_96__43_, s_r_96__42_, s_r_96__41_, s_r_96__40_, s_r_96__39_, s_r_96__38_, s_r_96__37_, s_r_96__36_, s_r_96__35_, s_r_96__34_, s_r_96__33_, s_r_96__32_, s_r_96__31_, s_r_96__30_, s_r_96__29_, s_r_96__28_, s_r_96__27_, s_r_96__26_, s_r_96__25_, s_r_96__24_, s_r_96__23_, s_r_96__22_, s_r_96__21_, s_r_96__20_, s_r_96__19_, s_r_96__18_, s_r_96__17_, s_r_96__16_, s_r_96__15_, s_r_96__14_, s_r_96__13_, s_r_96__12_, s_r_96__11_, s_r_96__10_, s_r_96__9_, s_r_96__8_, s_r_96__7_, s_r_96__6_, s_r_96__5_, s_r_96__4_, s_r_96__3_, s_r_96__2_, s_r_96__1_, s_r_96__0_ }),
    .c_i(c_r[96]),
    .prod_accum_i({ prod_accum_96__97_, prod_accum_96__96_, prod_accum_96__95_, prod_accum_96__94_, prod_accum_96__93_, prod_accum_96__92_, prod_accum_96__91_, prod_accum_96__90_, prod_accum_96__89_, prod_accum_96__88_, prod_accum_96__87_, prod_accum_96__86_, prod_accum_96__85_, prod_accum_96__84_, prod_accum_96__83_, prod_accum_96__82_, prod_accum_96__81_, prod_accum_96__80_, prod_accum_96__79_, prod_accum_96__78_, prod_accum_96__77_, prod_accum_96__76_, prod_accum_96__75_, prod_accum_96__74_, prod_accum_96__73_, prod_accum_96__72_, prod_accum_96__71_, prod_accum_96__70_, prod_accum_96__69_, prod_accum_96__68_, prod_accum_96__67_, prod_accum_96__66_, prod_accum_96__65_, prod_accum_96__64_, prod_accum_96__63_, prod_accum_96__62_, prod_accum_96__61_, prod_accum_96__60_, prod_accum_96__59_, prod_accum_96__58_, prod_accum_96__57_, prod_accum_96__56_, prod_accum_96__55_, prod_accum_96__54_, prod_accum_96__53_, prod_accum_96__52_, prod_accum_96__51_, prod_accum_96__50_, prod_accum_96__49_, prod_accum_96__48_, prod_accum_96__47_, prod_accum_96__46_, prod_accum_96__45_, prod_accum_96__44_, prod_accum_96__43_, prod_accum_96__42_, prod_accum_96__41_, prod_accum_96__40_, prod_accum_96__39_, prod_accum_96__38_, prod_accum_96__37_, prod_accum_96__36_, prod_accum_96__35_, prod_accum_96__34_, prod_accum_96__33_, prod_accum_96__32_, prod_accum_96__31_, prod_accum_96__30_, prod_accum_96__29_, prod_accum_96__28_, prod_accum_96__27_, prod_accum_96__26_, prod_accum_96__25_, prod_accum_96__24_, prod_accum_96__23_, prod_accum_96__22_, prod_accum_96__21_, prod_accum_96__20_, prod_accum_96__19_, prod_accum_96__18_, prod_accum_96__17_, prod_accum_96__16_, prod_accum_96__15_, prod_accum_96__14_, prod_accum_96__13_, prod_accum_96__12_, prod_accum_96__11_, prod_accum_96__10_, prod_accum_96__9_, prod_accum_96__8_, prod_accum_96__7_, prod_accum_96__6_, prod_accum_96__5_, prod_accum_96__4_, prod_accum_96__3_, prod_accum_96__2_, prod_accum_96__1_, prod_accum_96__0_ }),
    .a_o(a_r[12543:12416]),
    .b_o(b_r[12543:12416]),
    .s_o({ s_r_97__127_, s_r_97__126_, s_r_97__125_, s_r_97__124_, s_r_97__123_, s_r_97__122_, s_r_97__121_, s_r_97__120_, s_r_97__119_, s_r_97__118_, s_r_97__117_, s_r_97__116_, s_r_97__115_, s_r_97__114_, s_r_97__113_, s_r_97__112_, s_r_97__111_, s_r_97__110_, s_r_97__109_, s_r_97__108_, s_r_97__107_, s_r_97__106_, s_r_97__105_, s_r_97__104_, s_r_97__103_, s_r_97__102_, s_r_97__101_, s_r_97__100_, s_r_97__99_, s_r_97__98_, s_r_97__97_, s_r_97__96_, s_r_97__95_, s_r_97__94_, s_r_97__93_, s_r_97__92_, s_r_97__91_, s_r_97__90_, s_r_97__89_, s_r_97__88_, s_r_97__87_, s_r_97__86_, s_r_97__85_, s_r_97__84_, s_r_97__83_, s_r_97__82_, s_r_97__81_, s_r_97__80_, s_r_97__79_, s_r_97__78_, s_r_97__77_, s_r_97__76_, s_r_97__75_, s_r_97__74_, s_r_97__73_, s_r_97__72_, s_r_97__71_, s_r_97__70_, s_r_97__69_, s_r_97__68_, s_r_97__67_, s_r_97__66_, s_r_97__65_, s_r_97__64_, s_r_97__63_, s_r_97__62_, s_r_97__61_, s_r_97__60_, s_r_97__59_, s_r_97__58_, s_r_97__57_, s_r_97__56_, s_r_97__55_, s_r_97__54_, s_r_97__53_, s_r_97__52_, s_r_97__51_, s_r_97__50_, s_r_97__49_, s_r_97__48_, s_r_97__47_, s_r_97__46_, s_r_97__45_, s_r_97__44_, s_r_97__43_, s_r_97__42_, s_r_97__41_, s_r_97__40_, s_r_97__39_, s_r_97__38_, s_r_97__37_, s_r_97__36_, s_r_97__35_, s_r_97__34_, s_r_97__33_, s_r_97__32_, s_r_97__31_, s_r_97__30_, s_r_97__29_, s_r_97__28_, s_r_97__27_, s_r_97__26_, s_r_97__25_, s_r_97__24_, s_r_97__23_, s_r_97__22_, s_r_97__21_, s_r_97__20_, s_r_97__19_, s_r_97__18_, s_r_97__17_, s_r_97__16_, s_r_97__15_, s_r_97__14_, s_r_97__13_, s_r_97__12_, s_r_97__11_, s_r_97__10_, s_r_97__9_, s_r_97__8_, s_r_97__7_, s_r_97__6_, s_r_97__5_, s_r_97__4_, s_r_97__3_, s_r_97__2_, s_r_97__1_, s_r_97__0_ }),
    .c_o(c_r[97]),
    .prod_accum_o({ prod_accum_97__98_, prod_accum_97__97_, prod_accum_97__96_, prod_accum_97__95_, prod_accum_97__94_, prod_accum_97__93_, prod_accum_97__92_, prod_accum_97__91_, prod_accum_97__90_, prod_accum_97__89_, prod_accum_97__88_, prod_accum_97__87_, prod_accum_97__86_, prod_accum_97__85_, prod_accum_97__84_, prod_accum_97__83_, prod_accum_97__82_, prod_accum_97__81_, prod_accum_97__80_, prod_accum_97__79_, prod_accum_97__78_, prod_accum_97__77_, prod_accum_97__76_, prod_accum_97__75_, prod_accum_97__74_, prod_accum_97__73_, prod_accum_97__72_, prod_accum_97__71_, prod_accum_97__70_, prod_accum_97__69_, prod_accum_97__68_, prod_accum_97__67_, prod_accum_97__66_, prod_accum_97__65_, prod_accum_97__64_, prod_accum_97__63_, prod_accum_97__62_, prod_accum_97__61_, prod_accum_97__60_, prod_accum_97__59_, prod_accum_97__58_, prod_accum_97__57_, prod_accum_97__56_, prod_accum_97__55_, prod_accum_97__54_, prod_accum_97__53_, prod_accum_97__52_, prod_accum_97__51_, prod_accum_97__50_, prod_accum_97__49_, prod_accum_97__48_, prod_accum_97__47_, prod_accum_97__46_, prod_accum_97__45_, prod_accum_97__44_, prod_accum_97__43_, prod_accum_97__42_, prod_accum_97__41_, prod_accum_97__40_, prod_accum_97__39_, prod_accum_97__38_, prod_accum_97__37_, prod_accum_97__36_, prod_accum_97__35_, prod_accum_97__34_, prod_accum_97__33_, prod_accum_97__32_, prod_accum_97__31_, prod_accum_97__30_, prod_accum_97__29_, prod_accum_97__28_, prod_accum_97__27_, prod_accum_97__26_, prod_accum_97__25_, prod_accum_97__24_, prod_accum_97__23_, prod_accum_97__22_, prod_accum_97__21_, prod_accum_97__20_, prod_accum_97__19_, prod_accum_97__18_, prod_accum_97__17_, prod_accum_97__16_, prod_accum_97__15_, prod_accum_97__14_, prod_accum_97__13_, prod_accum_97__12_, prod_accum_97__11_, prod_accum_97__10_, prod_accum_97__9_, prod_accum_97__8_, prod_accum_97__7_, prod_accum_97__6_, prod_accum_97__5_, prod_accum_97__4_, prod_accum_97__3_, prod_accum_97__2_, prod_accum_97__1_, prod_accum_97__0_ })
  );


  bsg_mul_array_row_128_98_x
  genblk1_98__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[12543:12416]),
    .b_i(b_r[12543:12416]),
    .s_i({ s_r_97__127_, s_r_97__126_, s_r_97__125_, s_r_97__124_, s_r_97__123_, s_r_97__122_, s_r_97__121_, s_r_97__120_, s_r_97__119_, s_r_97__118_, s_r_97__117_, s_r_97__116_, s_r_97__115_, s_r_97__114_, s_r_97__113_, s_r_97__112_, s_r_97__111_, s_r_97__110_, s_r_97__109_, s_r_97__108_, s_r_97__107_, s_r_97__106_, s_r_97__105_, s_r_97__104_, s_r_97__103_, s_r_97__102_, s_r_97__101_, s_r_97__100_, s_r_97__99_, s_r_97__98_, s_r_97__97_, s_r_97__96_, s_r_97__95_, s_r_97__94_, s_r_97__93_, s_r_97__92_, s_r_97__91_, s_r_97__90_, s_r_97__89_, s_r_97__88_, s_r_97__87_, s_r_97__86_, s_r_97__85_, s_r_97__84_, s_r_97__83_, s_r_97__82_, s_r_97__81_, s_r_97__80_, s_r_97__79_, s_r_97__78_, s_r_97__77_, s_r_97__76_, s_r_97__75_, s_r_97__74_, s_r_97__73_, s_r_97__72_, s_r_97__71_, s_r_97__70_, s_r_97__69_, s_r_97__68_, s_r_97__67_, s_r_97__66_, s_r_97__65_, s_r_97__64_, s_r_97__63_, s_r_97__62_, s_r_97__61_, s_r_97__60_, s_r_97__59_, s_r_97__58_, s_r_97__57_, s_r_97__56_, s_r_97__55_, s_r_97__54_, s_r_97__53_, s_r_97__52_, s_r_97__51_, s_r_97__50_, s_r_97__49_, s_r_97__48_, s_r_97__47_, s_r_97__46_, s_r_97__45_, s_r_97__44_, s_r_97__43_, s_r_97__42_, s_r_97__41_, s_r_97__40_, s_r_97__39_, s_r_97__38_, s_r_97__37_, s_r_97__36_, s_r_97__35_, s_r_97__34_, s_r_97__33_, s_r_97__32_, s_r_97__31_, s_r_97__30_, s_r_97__29_, s_r_97__28_, s_r_97__27_, s_r_97__26_, s_r_97__25_, s_r_97__24_, s_r_97__23_, s_r_97__22_, s_r_97__21_, s_r_97__20_, s_r_97__19_, s_r_97__18_, s_r_97__17_, s_r_97__16_, s_r_97__15_, s_r_97__14_, s_r_97__13_, s_r_97__12_, s_r_97__11_, s_r_97__10_, s_r_97__9_, s_r_97__8_, s_r_97__7_, s_r_97__6_, s_r_97__5_, s_r_97__4_, s_r_97__3_, s_r_97__2_, s_r_97__1_, s_r_97__0_ }),
    .c_i(c_r[97]),
    .prod_accum_i({ prod_accum_97__98_, prod_accum_97__97_, prod_accum_97__96_, prod_accum_97__95_, prod_accum_97__94_, prod_accum_97__93_, prod_accum_97__92_, prod_accum_97__91_, prod_accum_97__90_, prod_accum_97__89_, prod_accum_97__88_, prod_accum_97__87_, prod_accum_97__86_, prod_accum_97__85_, prod_accum_97__84_, prod_accum_97__83_, prod_accum_97__82_, prod_accum_97__81_, prod_accum_97__80_, prod_accum_97__79_, prod_accum_97__78_, prod_accum_97__77_, prod_accum_97__76_, prod_accum_97__75_, prod_accum_97__74_, prod_accum_97__73_, prod_accum_97__72_, prod_accum_97__71_, prod_accum_97__70_, prod_accum_97__69_, prod_accum_97__68_, prod_accum_97__67_, prod_accum_97__66_, prod_accum_97__65_, prod_accum_97__64_, prod_accum_97__63_, prod_accum_97__62_, prod_accum_97__61_, prod_accum_97__60_, prod_accum_97__59_, prod_accum_97__58_, prod_accum_97__57_, prod_accum_97__56_, prod_accum_97__55_, prod_accum_97__54_, prod_accum_97__53_, prod_accum_97__52_, prod_accum_97__51_, prod_accum_97__50_, prod_accum_97__49_, prod_accum_97__48_, prod_accum_97__47_, prod_accum_97__46_, prod_accum_97__45_, prod_accum_97__44_, prod_accum_97__43_, prod_accum_97__42_, prod_accum_97__41_, prod_accum_97__40_, prod_accum_97__39_, prod_accum_97__38_, prod_accum_97__37_, prod_accum_97__36_, prod_accum_97__35_, prod_accum_97__34_, prod_accum_97__33_, prod_accum_97__32_, prod_accum_97__31_, prod_accum_97__30_, prod_accum_97__29_, prod_accum_97__28_, prod_accum_97__27_, prod_accum_97__26_, prod_accum_97__25_, prod_accum_97__24_, prod_accum_97__23_, prod_accum_97__22_, prod_accum_97__21_, prod_accum_97__20_, prod_accum_97__19_, prod_accum_97__18_, prod_accum_97__17_, prod_accum_97__16_, prod_accum_97__15_, prod_accum_97__14_, prod_accum_97__13_, prod_accum_97__12_, prod_accum_97__11_, prod_accum_97__10_, prod_accum_97__9_, prod_accum_97__8_, prod_accum_97__7_, prod_accum_97__6_, prod_accum_97__5_, prod_accum_97__4_, prod_accum_97__3_, prod_accum_97__2_, prod_accum_97__1_, prod_accum_97__0_ }),
    .a_o(a_r[12671:12544]),
    .b_o(b_r[12671:12544]),
    .s_o({ s_r_98__127_, s_r_98__126_, s_r_98__125_, s_r_98__124_, s_r_98__123_, s_r_98__122_, s_r_98__121_, s_r_98__120_, s_r_98__119_, s_r_98__118_, s_r_98__117_, s_r_98__116_, s_r_98__115_, s_r_98__114_, s_r_98__113_, s_r_98__112_, s_r_98__111_, s_r_98__110_, s_r_98__109_, s_r_98__108_, s_r_98__107_, s_r_98__106_, s_r_98__105_, s_r_98__104_, s_r_98__103_, s_r_98__102_, s_r_98__101_, s_r_98__100_, s_r_98__99_, s_r_98__98_, s_r_98__97_, s_r_98__96_, s_r_98__95_, s_r_98__94_, s_r_98__93_, s_r_98__92_, s_r_98__91_, s_r_98__90_, s_r_98__89_, s_r_98__88_, s_r_98__87_, s_r_98__86_, s_r_98__85_, s_r_98__84_, s_r_98__83_, s_r_98__82_, s_r_98__81_, s_r_98__80_, s_r_98__79_, s_r_98__78_, s_r_98__77_, s_r_98__76_, s_r_98__75_, s_r_98__74_, s_r_98__73_, s_r_98__72_, s_r_98__71_, s_r_98__70_, s_r_98__69_, s_r_98__68_, s_r_98__67_, s_r_98__66_, s_r_98__65_, s_r_98__64_, s_r_98__63_, s_r_98__62_, s_r_98__61_, s_r_98__60_, s_r_98__59_, s_r_98__58_, s_r_98__57_, s_r_98__56_, s_r_98__55_, s_r_98__54_, s_r_98__53_, s_r_98__52_, s_r_98__51_, s_r_98__50_, s_r_98__49_, s_r_98__48_, s_r_98__47_, s_r_98__46_, s_r_98__45_, s_r_98__44_, s_r_98__43_, s_r_98__42_, s_r_98__41_, s_r_98__40_, s_r_98__39_, s_r_98__38_, s_r_98__37_, s_r_98__36_, s_r_98__35_, s_r_98__34_, s_r_98__33_, s_r_98__32_, s_r_98__31_, s_r_98__30_, s_r_98__29_, s_r_98__28_, s_r_98__27_, s_r_98__26_, s_r_98__25_, s_r_98__24_, s_r_98__23_, s_r_98__22_, s_r_98__21_, s_r_98__20_, s_r_98__19_, s_r_98__18_, s_r_98__17_, s_r_98__16_, s_r_98__15_, s_r_98__14_, s_r_98__13_, s_r_98__12_, s_r_98__11_, s_r_98__10_, s_r_98__9_, s_r_98__8_, s_r_98__7_, s_r_98__6_, s_r_98__5_, s_r_98__4_, s_r_98__3_, s_r_98__2_, s_r_98__1_, s_r_98__0_ }),
    .c_o(c_r[98]),
    .prod_accum_o({ prod_accum_98__99_, prod_accum_98__98_, prod_accum_98__97_, prod_accum_98__96_, prod_accum_98__95_, prod_accum_98__94_, prod_accum_98__93_, prod_accum_98__92_, prod_accum_98__91_, prod_accum_98__90_, prod_accum_98__89_, prod_accum_98__88_, prod_accum_98__87_, prod_accum_98__86_, prod_accum_98__85_, prod_accum_98__84_, prod_accum_98__83_, prod_accum_98__82_, prod_accum_98__81_, prod_accum_98__80_, prod_accum_98__79_, prod_accum_98__78_, prod_accum_98__77_, prod_accum_98__76_, prod_accum_98__75_, prod_accum_98__74_, prod_accum_98__73_, prod_accum_98__72_, prod_accum_98__71_, prod_accum_98__70_, prod_accum_98__69_, prod_accum_98__68_, prod_accum_98__67_, prod_accum_98__66_, prod_accum_98__65_, prod_accum_98__64_, prod_accum_98__63_, prod_accum_98__62_, prod_accum_98__61_, prod_accum_98__60_, prod_accum_98__59_, prod_accum_98__58_, prod_accum_98__57_, prod_accum_98__56_, prod_accum_98__55_, prod_accum_98__54_, prod_accum_98__53_, prod_accum_98__52_, prod_accum_98__51_, prod_accum_98__50_, prod_accum_98__49_, prod_accum_98__48_, prod_accum_98__47_, prod_accum_98__46_, prod_accum_98__45_, prod_accum_98__44_, prod_accum_98__43_, prod_accum_98__42_, prod_accum_98__41_, prod_accum_98__40_, prod_accum_98__39_, prod_accum_98__38_, prod_accum_98__37_, prod_accum_98__36_, prod_accum_98__35_, prod_accum_98__34_, prod_accum_98__33_, prod_accum_98__32_, prod_accum_98__31_, prod_accum_98__30_, prod_accum_98__29_, prod_accum_98__28_, prod_accum_98__27_, prod_accum_98__26_, prod_accum_98__25_, prod_accum_98__24_, prod_accum_98__23_, prod_accum_98__22_, prod_accum_98__21_, prod_accum_98__20_, prod_accum_98__19_, prod_accum_98__18_, prod_accum_98__17_, prod_accum_98__16_, prod_accum_98__15_, prod_accum_98__14_, prod_accum_98__13_, prod_accum_98__12_, prod_accum_98__11_, prod_accum_98__10_, prod_accum_98__9_, prod_accum_98__8_, prod_accum_98__7_, prod_accum_98__6_, prod_accum_98__5_, prod_accum_98__4_, prod_accum_98__3_, prod_accum_98__2_, prod_accum_98__1_, prod_accum_98__0_ })
  );


  bsg_mul_array_row_128_99_x
  genblk1_99__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[12671:12544]),
    .b_i(b_r[12671:12544]),
    .s_i({ s_r_98__127_, s_r_98__126_, s_r_98__125_, s_r_98__124_, s_r_98__123_, s_r_98__122_, s_r_98__121_, s_r_98__120_, s_r_98__119_, s_r_98__118_, s_r_98__117_, s_r_98__116_, s_r_98__115_, s_r_98__114_, s_r_98__113_, s_r_98__112_, s_r_98__111_, s_r_98__110_, s_r_98__109_, s_r_98__108_, s_r_98__107_, s_r_98__106_, s_r_98__105_, s_r_98__104_, s_r_98__103_, s_r_98__102_, s_r_98__101_, s_r_98__100_, s_r_98__99_, s_r_98__98_, s_r_98__97_, s_r_98__96_, s_r_98__95_, s_r_98__94_, s_r_98__93_, s_r_98__92_, s_r_98__91_, s_r_98__90_, s_r_98__89_, s_r_98__88_, s_r_98__87_, s_r_98__86_, s_r_98__85_, s_r_98__84_, s_r_98__83_, s_r_98__82_, s_r_98__81_, s_r_98__80_, s_r_98__79_, s_r_98__78_, s_r_98__77_, s_r_98__76_, s_r_98__75_, s_r_98__74_, s_r_98__73_, s_r_98__72_, s_r_98__71_, s_r_98__70_, s_r_98__69_, s_r_98__68_, s_r_98__67_, s_r_98__66_, s_r_98__65_, s_r_98__64_, s_r_98__63_, s_r_98__62_, s_r_98__61_, s_r_98__60_, s_r_98__59_, s_r_98__58_, s_r_98__57_, s_r_98__56_, s_r_98__55_, s_r_98__54_, s_r_98__53_, s_r_98__52_, s_r_98__51_, s_r_98__50_, s_r_98__49_, s_r_98__48_, s_r_98__47_, s_r_98__46_, s_r_98__45_, s_r_98__44_, s_r_98__43_, s_r_98__42_, s_r_98__41_, s_r_98__40_, s_r_98__39_, s_r_98__38_, s_r_98__37_, s_r_98__36_, s_r_98__35_, s_r_98__34_, s_r_98__33_, s_r_98__32_, s_r_98__31_, s_r_98__30_, s_r_98__29_, s_r_98__28_, s_r_98__27_, s_r_98__26_, s_r_98__25_, s_r_98__24_, s_r_98__23_, s_r_98__22_, s_r_98__21_, s_r_98__20_, s_r_98__19_, s_r_98__18_, s_r_98__17_, s_r_98__16_, s_r_98__15_, s_r_98__14_, s_r_98__13_, s_r_98__12_, s_r_98__11_, s_r_98__10_, s_r_98__9_, s_r_98__8_, s_r_98__7_, s_r_98__6_, s_r_98__5_, s_r_98__4_, s_r_98__3_, s_r_98__2_, s_r_98__1_, s_r_98__0_ }),
    .c_i(c_r[98]),
    .prod_accum_i({ prod_accum_98__99_, prod_accum_98__98_, prod_accum_98__97_, prod_accum_98__96_, prod_accum_98__95_, prod_accum_98__94_, prod_accum_98__93_, prod_accum_98__92_, prod_accum_98__91_, prod_accum_98__90_, prod_accum_98__89_, prod_accum_98__88_, prod_accum_98__87_, prod_accum_98__86_, prod_accum_98__85_, prod_accum_98__84_, prod_accum_98__83_, prod_accum_98__82_, prod_accum_98__81_, prod_accum_98__80_, prod_accum_98__79_, prod_accum_98__78_, prod_accum_98__77_, prod_accum_98__76_, prod_accum_98__75_, prod_accum_98__74_, prod_accum_98__73_, prod_accum_98__72_, prod_accum_98__71_, prod_accum_98__70_, prod_accum_98__69_, prod_accum_98__68_, prod_accum_98__67_, prod_accum_98__66_, prod_accum_98__65_, prod_accum_98__64_, prod_accum_98__63_, prod_accum_98__62_, prod_accum_98__61_, prod_accum_98__60_, prod_accum_98__59_, prod_accum_98__58_, prod_accum_98__57_, prod_accum_98__56_, prod_accum_98__55_, prod_accum_98__54_, prod_accum_98__53_, prod_accum_98__52_, prod_accum_98__51_, prod_accum_98__50_, prod_accum_98__49_, prod_accum_98__48_, prod_accum_98__47_, prod_accum_98__46_, prod_accum_98__45_, prod_accum_98__44_, prod_accum_98__43_, prod_accum_98__42_, prod_accum_98__41_, prod_accum_98__40_, prod_accum_98__39_, prod_accum_98__38_, prod_accum_98__37_, prod_accum_98__36_, prod_accum_98__35_, prod_accum_98__34_, prod_accum_98__33_, prod_accum_98__32_, prod_accum_98__31_, prod_accum_98__30_, prod_accum_98__29_, prod_accum_98__28_, prod_accum_98__27_, prod_accum_98__26_, prod_accum_98__25_, prod_accum_98__24_, prod_accum_98__23_, prod_accum_98__22_, prod_accum_98__21_, prod_accum_98__20_, prod_accum_98__19_, prod_accum_98__18_, prod_accum_98__17_, prod_accum_98__16_, prod_accum_98__15_, prod_accum_98__14_, prod_accum_98__13_, prod_accum_98__12_, prod_accum_98__11_, prod_accum_98__10_, prod_accum_98__9_, prod_accum_98__8_, prod_accum_98__7_, prod_accum_98__6_, prod_accum_98__5_, prod_accum_98__4_, prod_accum_98__3_, prod_accum_98__2_, prod_accum_98__1_, prod_accum_98__0_ }),
    .a_o(a_r[12799:12672]),
    .b_o(b_r[12799:12672]),
    .s_o({ s_r_99__127_, s_r_99__126_, s_r_99__125_, s_r_99__124_, s_r_99__123_, s_r_99__122_, s_r_99__121_, s_r_99__120_, s_r_99__119_, s_r_99__118_, s_r_99__117_, s_r_99__116_, s_r_99__115_, s_r_99__114_, s_r_99__113_, s_r_99__112_, s_r_99__111_, s_r_99__110_, s_r_99__109_, s_r_99__108_, s_r_99__107_, s_r_99__106_, s_r_99__105_, s_r_99__104_, s_r_99__103_, s_r_99__102_, s_r_99__101_, s_r_99__100_, s_r_99__99_, s_r_99__98_, s_r_99__97_, s_r_99__96_, s_r_99__95_, s_r_99__94_, s_r_99__93_, s_r_99__92_, s_r_99__91_, s_r_99__90_, s_r_99__89_, s_r_99__88_, s_r_99__87_, s_r_99__86_, s_r_99__85_, s_r_99__84_, s_r_99__83_, s_r_99__82_, s_r_99__81_, s_r_99__80_, s_r_99__79_, s_r_99__78_, s_r_99__77_, s_r_99__76_, s_r_99__75_, s_r_99__74_, s_r_99__73_, s_r_99__72_, s_r_99__71_, s_r_99__70_, s_r_99__69_, s_r_99__68_, s_r_99__67_, s_r_99__66_, s_r_99__65_, s_r_99__64_, s_r_99__63_, s_r_99__62_, s_r_99__61_, s_r_99__60_, s_r_99__59_, s_r_99__58_, s_r_99__57_, s_r_99__56_, s_r_99__55_, s_r_99__54_, s_r_99__53_, s_r_99__52_, s_r_99__51_, s_r_99__50_, s_r_99__49_, s_r_99__48_, s_r_99__47_, s_r_99__46_, s_r_99__45_, s_r_99__44_, s_r_99__43_, s_r_99__42_, s_r_99__41_, s_r_99__40_, s_r_99__39_, s_r_99__38_, s_r_99__37_, s_r_99__36_, s_r_99__35_, s_r_99__34_, s_r_99__33_, s_r_99__32_, s_r_99__31_, s_r_99__30_, s_r_99__29_, s_r_99__28_, s_r_99__27_, s_r_99__26_, s_r_99__25_, s_r_99__24_, s_r_99__23_, s_r_99__22_, s_r_99__21_, s_r_99__20_, s_r_99__19_, s_r_99__18_, s_r_99__17_, s_r_99__16_, s_r_99__15_, s_r_99__14_, s_r_99__13_, s_r_99__12_, s_r_99__11_, s_r_99__10_, s_r_99__9_, s_r_99__8_, s_r_99__7_, s_r_99__6_, s_r_99__5_, s_r_99__4_, s_r_99__3_, s_r_99__2_, s_r_99__1_, s_r_99__0_ }),
    .c_o(c_r[99]),
    .prod_accum_o({ prod_accum_99__100_, prod_accum_99__99_, prod_accum_99__98_, prod_accum_99__97_, prod_accum_99__96_, prod_accum_99__95_, prod_accum_99__94_, prod_accum_99__93_, prod_accum_99__92_, prod_accum_99__91_, prod_accum_99__90_, prod_accum_99__89_, prod_accum_99__88_, prod_accum_99__87_, prod_accum_99__86_, prod_accum_99__85_, prod_accum_99__84_, prod_accum_99__83_, prod_accum_99__82_, prod_accum_99__81_, prod_accum_99__80_, prod_accum_99__79_, prod_accum_99__78_, prod_accum_99__77_, prod_accum_99__76_, prod_accum_99__75_, prod_accum_99__74_, prod_accum_99__73_, prod_accum_99__72_, prod_accum_99__71_, prod_accum_99__70_, prod_accum_99__69_, prod_accum_99__68_, prod_accum_99__67_, prod_accum_99__66_, prod_accum_99__65_, prod_accum_99__64_, prod_accum_99__63_, prod_accum_99__62_, prod_accum_99__61_, prod_accum_99__60_, prod_accum_99__59_, prod_accum_99__58_, prod_accum_99__57_, prod_accum_99__56_, prod_accum_99__55_, prod_accum_99__54_, prod_accum_99__53_, prod_accum_99__52_, prod_accum_99__51_, prod_accum_99__50_, prod_accum_99__49_, prod_accum_99__48_, prod_accum_99__47_, prod_accum_99__46_, prod_accum_99__45_, prod_accum_99__44_, prod_accum_99__43_, prod_accum_99__42_, prod_accum_99__41_, prod_accum_99__40_, prod_accum_99__39_, prod_accum_99__38_, prod_accum_99__37_, prod_accum_99__36_, prod_accum_99__35_, prod_accum_99__34_, prod_accum_99__33_, prod_accum_99__32_, prod_accum_99__31_, prod_accum_99__30_, prod_accum_99__29_, prod_accum_99__28_, prod_accum_99__27_, prod_accum_99__26_, prod_accum_99__25_, prod_accum_99__24_, prod_accum_99__23_, prod_accum_99__22_, prod_accum_99__21_, prod_accum_99__20_, prod_accum_99__19_, prod_accum_99__18_, prod_accum_99__17_, prod_accum_99__16_, prod_accum_99__15_, prod_accum_99__14_, prod_accum_99__13_, prod_accum_99__12_, prod_accum_99__11_, prod_accum_99__10_, prod_accum_99__9_, prod_accum_99__8_, prod_accum_99__7_, prod_accum_99__6_, prod_accum_99__5_, prod_accum_99__4_, prod_accum_99__3_, prod_accum_99__2_, prod_accum_99__1_, prod_accum_99__0_ })
  );


  bsg_mul_array_row_128_100_x
  genblk1_100__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[12799:12672]),
    .b_i(b_r[12799:12672]),
    .s_i({ s_r_99__127_, s_r_99__126_, s_r_99__125_, s_r_99__124_, s_r_99__123_, s_r_99__122_, s_r_99__121_, s_r_99__120_, s_r_99__119_, s_r_99__118_, s_r_99__117_, s_r_99__116_, s_r_99__115_, s_r_99__114_, s_r_99__113_, s_r_99__112_, s_r_99__111_, s_r_99__110_, s_r_99__109_, s_r_99__108_, s_r_99__107_, s_r_99__106_, s_r_99__105_, s_r_99__104_, s_r_99__103_, s_r_99__102_, s_r_99__101_, s_r_99__100_, s_r_99__99_, s_r_99__98_, s_r_99__97_, s_r_99__96_, s_r_99__95_, s_r_99__94_, s_r_99__93_, s_r_99__92_, s_r_99__91_, s_r_99__90_, s_r_99__89_, s_r_99__88_, s_r_99__87_, s_r_99__86_, s_r_99__85_, s_r_99__84_, s_r_99__83_, s_r_99__82_, s_r_99__81_, s_r_99__80_, s_r_99__79_, s_r_99__78_, s_r_99__77_, s_r_99__76_, s_r_99__75_, s_r_99__74_, s_r_99__73_, s_r_99__72_, s_r_99__71_, s_r_99__70_, s_r_99__69_, s_r_99__68_, s_r_99__67_, s_r_99__66_, s_r_99__65_, s_r_99__64_, s_r_99__63_, s_r_99__62_, s_r_99__61_, s_r_99__60_, s_r_99__59_, s_r_99__58_, s_r_99__57_, s_r_99__56_, s_r_99__55_, s_r_99__54_, s_r_99__53_, s_r_99__52_, s_r_99__51_, s_r_99__50_, s_r_99__49_, s_r_99__48_, s_r_99__47_, s_r_99__46_, s_r_99__45_, s_r_99__44_, s_r_99__43_, s_r_99__42_, s_r_99__41_, s_r_99__40_, s_r_99__39_, s_r_99__38_, s_r_99__37_, s_r_99__36_, s_r_99__35_, s_r_99__34_, s_r_99__33_, s_r_99__32_, s_r_99__31_, s_r_99__30_, s_r_99__29_, s_r_99__28_, s_r_99__27_, s_r_99__26_, s_r_99__25_, s_r_99__24_, s_r_99__23_, s_r_99__22_, s_r_99__21_, s_r_99__20_, s_r_99__19_, s_r_99__18_, s_r_99__17_, s_r_99__16_, s_r_99__15_, s_r_99__14_, s_r_99__13_, s_r_99__12_, s_r_99__11_, s_r_99__10_, s_r_99__9_, s_r_99__8_, s_r_99__7_, s_r_99__6_, s_r_99__5_, s_r_99__4_, s_r_99__3_, s_r_99__2_, s_r_99__1_, s_r_99__0_ }),
    .c_i(c_r[99]),
    .prod_accum_i({ prod_accum_99__100_, prod_accum_99__99_, prod_accum_99__98_, prod_accum_99__97_, prod_accum_99__96_, prod_accum_99__95_, prod_accum_99__94_, prod_accum_99__93_, prod_accum_99__92_, prod_accum_99__91_, prod_accum_99__90_, prod_accum_99__89_, prod_accum_99__88_, prod_accum_99__87_, prod_accum_99__86_, prod_accum_99__85_, prod_accum_99__84_, prod_accum_99__83_, prod_accum_99__82_, prod_accum_99__81_, prod_accum_99__80_, prod_accum_99__79_, prod_accum_99__78_, prod_accum_99__77_, prod_accum_99__76_, prod_accum_99__75_, prod_accum_99__74_, prod_accum_99__73_, prod_accum_99__72_, prod_accum_99__71_, prod_accum_99__70_, prod_accum_99__69_, prod_accum_99__68_, prod_accum_99__67_, prod_accum_99__66_, prod_accum_99__65_, prod_accum_99__64_, prod_accum_99__63_, prod_accum_99__62_, prod_accum_99__61_, prod_accum_99__60_, prod_accum_99__59_, prod_accum_99__58_, prod_accum_99__57_, prod_accum_99__56_, prod_accum_99__55_, prod_accum_99__54_, prod_accum_99__53_, prod_accum_99__52_, prod_accum_99__51_, prod_accum_99__50_, prod_accum_99__49_, prod_accum_99__48_, prod_accum_99__47_, prod_accum_99__46_, prod_accum_99__45_, prod_accum_99__44_, prod_accum_99__43_, prod_accum_99__42_, prod_accum_99__41_, prod_accum_99__40_, prod_accum_99__39_, prod_accum_99__38_, prod_accum_99__37_, prod_accum_99__36_, prod_accum_99__35_, prod_accum_99__34_, prod_accum_99__33_, prod_accum_99__32_, prod_accum_99__31_, prod_accum_99__30_, prod_accum_99__29_, prod_accum_99__28_, prod_accum_99__27_, prod_accum_99__26_, prod_accum_99__25_, prod_accum_99__24_, prod_accum_99__23_, prod_accum_99__22_, prod_accum_99__21_, prod_accum_99__20_, prod_accum_99__19_, prod_accum_99__18_, prod_accum_99__17_, prod_accum_99__16_, prod_accum_99__15_, prod_accum_99__14_, prod_accum_99__13_, prod_accum_99__12_, prod_accum_99__11_, prod_accum_99__10_, prod_accum_99__9_, prod_accum_99__8_, prod_accum_99__7_, prod_accum_99__6_, prod_accum_99__5_, prod_accum_99__4_, prod_accum_99__3_, prod_accum_99__2_, prod_accum_99__1_, prod_accum_99__0_ }),
    .a_o(a_r[12927:12800]),
    .b_o(b_r[12927:12800]),
    .s_o({ s_r_100__127_, s_r_100__126_, s_r_100__125_, s_r_100__124_, s_r_100__123_, s_r_100__122_, s_r_100__121_, s_r_100__120_, s_r_100__119_, s_r_100__118_, s_r_100__117_, s_r_100__116_, s_r_100__115_, s_r_100__114_, s_r_100__113_, s_r_100__112_, s_r_100__111_, s_r_100__110_, s_r_100__109_, s_r_100__108_, s_r_100__107_, s_r_100__106_, s_r_100__105_, s_r_100__104_, s_r_100__103_, s_r_100__102_, s_r_100__101_, s_r_100__100_, s_r_100__99_, s_r_100__98_, s_r_100__97_, s_r_100__96_, s_r_100__95_, s_r_100__94_, s_r_100__93_, s_r_100__92_, s_r_100__91_, s_r_100__90_, s_r_100__89_, s_r_100__88_, s_r_100__87_, s_r_100__86_, s_r_100__85_, s_r_100__84_, s_r_100__83_, s_r_100__82_, s_r_100__81_, s_r_100__80_, s_r_100__79_, s_r_100__78_, s_r_100__77_, s_r_100__76_, s_r_100__75_, s_r_100__74_, s_r_100__73_, s_r_100__72_, s_r_100__71_, s_r_100__70_, s_r_100__69_, s_r_100__68_, s_r_100__67_, s_r_100__66_, s_r_100__65_, s_r_100__64_, s_r_100__63_, s_r_100__62_, s_r_100__61_, s_r_100__60_, s_r_100__59_, s_r_100__58_, s_r_100__57_, s_r_100__56_, s_r_100__55_, s_r_100__54_, s_r_100__53_, s_r_100__52_, s_r_100__51_, s_r_100__50_, s_r_100__49_, s_r_100__48_, s_r_100__47_, s_r_100__46_, s_r_100__45_, s_r_100__44_, s_r_100__43_, s_r_100__42_, s_r_100__41_, s_r_100__40_, s_r_100__39_, s_r_100__38_, s_r_100__37_, s_r_100__36_, s_r_100__35_, s_r_100__34_, s_r_100__33_, s_r_100__32_, s_r_100__31_, s_r_100__30_, s_r_100__29_, s_r_100__28_, s_r_100__27_, s_r_100__26_, s_r_100__25_, s_r_100__24_, s_r_100__23_, s_r_100__22_, s_r_100__21_, s_r_100__20_, s_r_100__19_, s_r_100__18_, s_r_100__17_, s_r_100__16_, s_r_100__15_, s_r_100__14_, s_r_100__13_, s_r_100__12_, s_r_100__11_, s_r_100__10_, s_r_100__9_, s_r_100__8_, s_r_100__7_, s_r_100__6_, s_r_100__5_, s_r_100__4_, s_r_100__3_, s_r_100__2_, s_r_100__1_, s_r_100__0_ }),
    .c_o(c_r[100]),
    .prod_accum_o({ prod_accum_100__101_, prod_accum_100__100_, prod_accum_100__99_, prod_accum_100__98_, prod_accum_100__97_, prod_accum_100__96_, prod_accum_100__95_, prod_accum_100__94_, prod_accum_100__93_, prod_accum_100__92_, prod_accum_100__91_, prod_accum_100__90_, prod_accum_100__89_, prod_accum_100__88_, prod_accum_100__87_, prod_accum_100__86_, prod_accum_100__85_, prod_accum_100__84_, prod_accum_100__83_, prod_accum_100__82_, prod_accum_100__81_, prod_accum_100__80_, prod_accum_100__79_, prod_accum_100__78_, prod_accum_100__77_, prod_accum_100__76_, prod_accum_100__75_, prod_accum_100__74_, prod_accum_100__73_, prod_accum_100__72_, prod_accum_100__71_, prod_accum_100__70_, prod_accum_100__69_, prod_accum_100__68_, prod_accum_100__67_, prod_accum_100__66_, prod_accum_100__65_, prod_accum_100__64_, prod_accum_100__63_, prod_accum_100__62_, prod_accum_100__61_, prod_accum_100__60_, prod_accum_100__59_, prod_accum_100__58_, prod_accum_100__57_, prod_accum_100__56_, prod_accum_100__55_, prod_accum_100__54_, prod_accum_100__53_, prod_accum_100__52_, prod_accum_100__51_, prod_accum_100__50_, prod_accum_100__49_, prod_accum_100__48_, prod_accum_100__47_, prod_accum_100__46_, prod_accum_100__45_, prod_accum_100__44_, prod_accum_100__43_, prod_accum_100__42_, prod_accum_100__41_, prod_accum_100__40_, prod_accum_100__39_, prod_accum_100__38_, prod_accum_100__37_, prod_accum_100__36_, prod_accum_100__35_, prod_accum_100__34_, prod_accum_100__33_, prod_accum_100__32_, prod_accum_100__31_, prod_accum_100__30_, prod_accum_100__29_, prod_accum_100__28_, prod_accum_100__27_, prod_accum_100__26_, prod_accum_100__25_, prod_accum_100__24_, prod_accum_100__23_, prod_accum_100__22_, prod_accum_100__21_, prod_accum_100__20_, prod_accum_100__19_, prod_accum_100__18_, prod_accum_100__17_, prod_accum_100__16_, prod_accum_100__15_, prod_accum_100__14_, prod_accum_100__13_, prod_accum_100__12_, prod_accum_100__11_, prod_accum_100__10_, prod_accum_100__9_, prod_accum_100__8_, prod_accum_100__7_, prod_accum_100__6_, prod_accum_100__5_, prod_accum_100__4_, prod_accum_100__3_, prod_accum_100__2_, prod_accum_100__1_, prod_accum_100__0_ })
  );


  bsg_mul_array_row_128_101_x
  genblk1_101__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[12927:12800]),
    .b_i(b_r[12927:12800]),
    .s_i({ s_r_100__127_, s_r_100__126_, s_r_100__125_, s_r_100__124_, s_r_100__123_, s_r_100__122_, s_r_100__121_, s_r_100__120_, s_r_100__119_, s_r_100__118_, s_r_100__117_, s_r_100__116_, s_r_100__115_, s_r_100__114_, s_r_100__113_, s_r_100__112_, s_r_100__111_, s_r_100__110_, s_r_100__109_, s_r_100__108_, s_r_100__107_, s_r_100__106_, s_r_100__105_, s_r_100__104_, s_r_100__103_, s_r_100__102_, s_r_100__101_, s_r_100__100_, s_r_100__99_, s_r_100__98_, s_r_100__97_, s_r_100__96_, s_r_100__95_, s_r_100__94_, s_r_100__93_, s_r_100__92_, s_r_100__91_, s_r_100__90_, s_r_100__89_, s_r_100__88_, s_r_100__87_, s_r_100__86_, s_r_100__85_, s_r_100__84_, s_r_100__83_, s_r_100__82_, s_r_100__81_, s_r_100__80_, s_r_100__79_, s_r_100__78_, s_r_100__77_, s_r_100__76_, s_r_100__75_, s_r_100__74_, s_r_100__73_, s_r_100__72_, s_r_100__71_, s_r_100__70_, s_r_100__69_, s_r_100__68_, s_r_100__67_, s_r_100__66_, s_r_100__65_, s_r_100__64_, s_r_100__63_, s_r_100__62_, s_r_100__61_, s_r_100__60_, s_r_100__59_, s_r_100__58_, s_r_100__57_, s_r_100__56_, s_r_100__55_, s_r_100__54_, s_r_100__53_, s_r_100__52_, s_r_100__51_, s_r_100__50_, s_r_100__49_, s_r_100__48_, s_r_100__47_, s_r_100__46_, s_r_100__45_, s_r_100__44_, s_r_100__43_, s_r_100__42_, s_r_100__41_, s_r_100__40_, s_r_100__39_, s_r_100__38_, s_r_100__37_, s_r_100__36_, s_r_100__35_, s_r_100__34_, s_r_100__33_, s_r_100__32_, s_r_100__31_, s_r_100__30_, s_r_100__29_, s_r_100__28_, s_r_100__27_, s_r_100__26_, s_r_100__25_, s_r_100__24_, s_r_100__23_, s_r_100__22_, s_r_100__21_, s_r_100__20_, s_r_100__19_, s_r_100__18_, s_r_100__17_, s_r_100__16_, s_r_100__15_, s_r_100__14_, s_r_100__13_, s_r_100__12_, s_r_100__11_, s_r_100__10_, s_r_100__9_, s_r_100__8_, s_r_100__7_, s_r_100__6_, s_r_100__5_, s_r_100__4_, s_r_100__3_, s_r_100__2_, s_r_100__1_, s_r_100__0_ }),
    .c_i(c_r[100]),
    .prod_accum_i({ prod_accum_100__101_, prod_accum_100__100_, prod_accum_100__99_, prod_accum_100__98_, prod_accum_100__97_, prod_accum_100__96_, prod_accum_100__95_, prod_accum_100__94_, prod_accum_100__93_, prod_accum_100__92_, prod_accum_100__91_, prod_accum_100__90_, prod_accum_100__89_, prod_accum_100__88_, prod_accum_100__87_, prod_accum_100__86_, prod_accum_100__85_, prod_accum_100__84_, prod_accum_100__83_, prod_accum_100__82_, prod_accum_100__81_, prod_accum_100__80_, prod_accum_100__79_, prod_accum_100__78_, prod_accum_100__77_, prod_accum_100__76_, prod_accum_100__75_, prod_accum_100__74_, prod_accum_100__73_, prod_accum_100__72_, prod_accum_100__71_, prod_accum_100__70_, prod_accum_100__69_, prod_accum_100__68_, prod_accum_100__67_, prod_accum_100__66_, prod_accum_100__65_, prod_accum_100__64_, prod_accum_100__63_, prod_accum_100__62_, prod_accum_100__61_, prod_accum_100__60_, prod_accum_100__59_, prod_accum_100__58_, prod_accum_100__57_, prod_accum_100__56_, prod_accum_100__55_, prod_accum_100__54_, prod_accum_100__53_, prod_accum_100__52_, prod_accum_100__51_, prod_accum_100__50_, prod_accum_100__49_, prod_accum_100__48_, prod_accum_100__47_, prod_accum_100__46_, prod_accum_100__45_, prod_accum_100__44_, prod_accum_100__43_, prod_accum_100__42_, prod_accum_100__41_, prod_accum_100__40_, prod_accum_100__39_, prod_accum_100__38_, prod_accum_100__37_, prod_accum_100__36_, prod_accum_100__35_, prod_accum_100__34_, prod_accum_100__33_, prod_accum_100__32_, prod_accum_100__31_, prod_accum_100__30_, prod_accum_100__29_, prod_accum_100__28_, prod_accum_100__27_, prod_accum_100__26_, prod_accum_100__25_, prod_accum_100__24_, prod_accum_100__23_, prod_accum_100__22_, prod_accum_100__21_, prod_accum_100__20_, prod_accum_100__19_, prod_accum_100__18_, prod_accum_100__17_, prod_accum_100__16_, prod_accum_100__15_, prod_accum_100__14_, prod_accum_100__13_, prod_accum_100__12_, prod_accum_100__11_, prod_accum_100__10_, prod_accum_100__9_, prod_accum_100__8_, prod_accum_100__7_, prod_accum_100__6_, prod_accum_100__5_, prod_accum_100__4_, prod_accum_100__3_, prod_accum_100__2_, prod_accum_100__1_, prod_accum_100__0_ }),
    .a_o(a_r[13055:12928]),
    .b_o(b_r[13055:12928]),
    .s_o({ s_r_101__127_, s_r_101__126_, s_r_101__125_, s_r_101__124_, s_r_101__123_, s_r_101__122_, s_r_101__121_, s_r_101__120_, s_r_101__119_, s_r_101__118_, s_r_101__117_, s_r_101__116_, s_r_101__115_, s_r_101__114_, s_r_101__113_, s_r_101__112_, s_r_101__111_, s_r_101__110_, s_r_101__109_, s_r_101__108_, s_r_101__107_, s_r_101__106_, s_r_101__105_, s_r_101__104_, s_r_101__103_, s_r_101__102_, s_r_101__101_, s_r_101__100_, s_r_101__99_, s_r_101__98_, s_r_101__97_, s_r_101__96_, s_r_101__95_, s_r_101__94_, s_r_101__93_, s_r_101__92_, s_r_101__91_, s_r_101__90_, s_r_101__89_, s_r_101__88_, s_r_101__87_, s_r_101__86_, s_r_101__85_, s_r_101__84_, s_r_101__83_, s_r_101__82_, s_r_101__81_, s_r_101__80_, s_r_101__79_, s_r_101__78_, s_r_101__77_, s_r_101__76_, s_r_101__75_, s_r_101__74_, s_r_101__73_, s_r_101__72_, s_r_101__71_, s_r_101__70_, s_r_101__69_, s_r_101__68_, s_r_101__67_, s_r_101__66_, s_r_101__65_, s_r_101__64_, s_r_101__63_, s_r_101__62_, s_r_101__61_, s_r_101__60_, s_r_101__59_, s_r_101__58_, s_r_101__57_, s_r_101__56_, s_r_101__55_, s_r_101__54_, s_r_101__53_, s_r_101__52_, s_r_101__51_, s_r_101__50_, s_r_101__49_, s_r_101__48_, s_r_101__47_, s_r_101__46_, s_r_101__45_, s_r_101__44_, s_r_101__43_, s_r_101__42_, s_r_101__41_, s_r_101__40_, s_r_101__39_, s_r_101__38_, s_r_101__37_, s_r_101__36_, s_r_101__35_, s_r_101__34_, s_r_101__33_, s_r_101__32_, s_r_101__31_, s_r_101__30_, s_r_101__29_, s_r_101__28_, s_r_101__27_, s_r_101__26_, s_r_101__25_, s_r_101__24_, s_r_101__23_, s_r_101__22_, s_r_101__21_, s_r_101__20_, s_r_101__19_, s_r_101__18_, s_r_101__17_, s_r_101__16_, s_r_101__15_, s_r_101__14_, s_r_101__13_, s_r_101__12_, s_r_101__11_, s_r_101__10_, s_r_101__9_, s_r_101__8_, s_r_101__7_, s_r_101__6_, s_r_101__5_, s_r_101__4_, s_r_101__3_, s_r_101__2_, s_r_101__1_, s_r_101__0_ }),
    .c_o(c_r[101]),
    .prod_accum_o({ prod_accum_101__102_, prod_accum_101__101_, prod_accum_101__100_, prod_accum_101__99_, prod_accum_101__98_, prod_accum_101__97_, prod_accum_101__96_, prod_accum_101__95_, prod_accum_101__94_, prod_accum_101__93_, prod_accum_101__92_, prod_accum_101__91_, prod_accum_101__90_, prod_accum_101__89_, prod_accum_101__88_, prod_accum_101__87_, prod_accum_101__86_, prod_accum_101__85_, prod_accum_101__84_, prod_accum_101__83_, prod_accum_101__82_, prod_accum_101__81_, prod_accum_101__80_, prod_accum_101__79_, prod_accum_101__78_, prod_accum_101__77_, prod_accum_101__76_, prod_accum_101__75_, prod_accum_101__74_, prod_accum_101__73_, prod_accum_101__72_, prod_accum_101__71_, prod_accum_101__70_, prod_accum_101__69_, prod_accum_101__68_, prod_accum_101__67_, prod_accum_101__66_, prod_accum_101__65_, prod_accum_101__64_, prod_accum_101__63_, prod_accum_101__62_, prod_accum_101__61_, prod_accum_101__60_, prod_accum_101__59_, prod_accum_101__58_, prod_accum_101__57_, prod_accum_101__56_, prod_accum_101__55_, prod_accum_101__54_, prod_accum_101__53_, prod_accum_101__52_, prod_accum_101__51_, prod_accum_101__50_, prod_accum_101__49_, prod_accum_101__48_, prod_accum_101__47_, prod_accum_101__46_, prod_accum_101__45_, prod_accum_101__44_, prod_accum_101__43_, prod_accum_101__42_, prod_accum_101__41_, prod_accum_101__40_, prod_accum_101__39_, prod_accum_101__38_, prod_accum_101__37_, prod_accum_101__36_, prod_accum_101__35_, prod_accum_101__34_, prod_accum_101__33_, prod_accum_101__32_, prod_accum_101__31_, prod_accum_101__30_, prod_accum_101__29_, prod_accum_101__28_, prod_accum_101__27_, prod_accum_101__26_, prod_accum_101__25_, prod_accum_101__24_, prod_accum_101__23_, prod_accum_101__22_, prod_accum_101__21_, prod_accum_101__20_, prod_accum_101__19_, prod_accum_101__18_, prod_accum_101__17_, prod_accum_101__16_, prod_accum_101__15_, prod_accum_101__14_, prod_accum_101__13_, prod_accum_101__12_, prod_accum_101__11_, prod_accum_101__10_, prod_accum_101__9_, prod_accum_101__8_, prod_accum_101__7_, prod_accum_101__6_, prod_accum_101__5_, prod_accum_101__4_, prod_accum_101__3_, prod_accum_101__2_, prod_accum_101__1_, prod_accum_101__0_ })
  );


  bsg_mul_array_row_128_102_x
  genblk1_102__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[13055:12928]),
    .b_i(b_r[13055:12928]),
    .s_i({ s_r_101__127_, s_r_101__126_, s_r_101__125_, s_r_101__124_, s_r_101__123_, s_r_101__122_, s_r_101__121_, s_r_101__120_, s_r_101__119_, s_r_101__118_, s_r_101__117_, s_r_101__116_, s_r_101__115_, s_r_101__114_, s_r_101__113_, s_r_101__112_, s_r_101__111_, s_r_101__110_, s_r_101__109_, s_r_101__108_, s_r_101__107_, s_r_101__106_, s_r_101__105_, s_r_101__104_, s_r_101__103_, s_r_101__102_, s_r_101__101_, s_r_101__100_, s_r_101__99_, s_r_101__98_, s_r_101__97_, s_r_101__96_, s_r_101__95_, s_r_101__94_, s_r_101__93_, s_r_101__92_, s_r_101__91_, s_r_101__90_, s_r_101__89_, s_r_101__88_, s_r_101__87_, s_r_101__86_, s_r_101__85_, s_r_101__84_, s_r_101__83_, s_r_101__82_, s_r_101__81_, s_r_101__80_, s_r_101__79_, s_r_101__78_, s_r_101__77_, s_r_101__76_, s_r_101__75_, s_r_101__74_, s_r_101__73_, s_r_101__72_, s_r_101__71_, s_r_101__70_, s_r_101__69_, s_r_101__68_, s_r_101__67_, s_r_101__66_, s_r_101__65_, s_r_101__64_, s_r_101__63_, s_r_101__62_, s_r_101__61_, s_r_101__60_, s_r_101__59_, s_r_101__58_, s_r_101__57_, s_r_101__56_, s_r_101__55_, s_r_101__54_, s_r_101__53_, s_r_101__52_, s_r_101__51_, s_r_101__50_, s_r_101__49_, s_r_101__48_, s_r_101__47_, s_r_101__46_, s_r_101__45_, s_r_101__44_, s_r_101__43_, s_r_101__42_, s_r_101__41_, s_r_101__40_, s_r_101__39_, s_r_101__38_, s_r_101__37_, s_r_101__36_, s_r_101__35_, s_r_101__34_, s_r_101__33_, s_r_101__32_, s_r_101__31_, s_r_101__30_, s_r_101__29_, s_r_101__28_, s_r_101__27_, s_r_101__26_, s_r_101__25_, s_r_101__24_, s_r_101__23_, s_r_101__22_, s_r_101__21_, s_r_101__20_, s_r_101__19_, s_r_101__18_, s_r_101__17_, s_r_101__16_, s_r_101__15_, s_r_101__14_, s_r_101__13_, s_r_101__12_, s_r_101__11_, s_r_101__10_, s_r_101__9_, s_r_101__8_, s_r_101__7_, s_r_101__6_, s_r_101__5_, s_r_101__4_, s_r_101__3_, s_r_101__2_, s_r_101__1_, s_r_101__0_ }),
    .c_i(c_r[101]),
    .prod_accum_i({ prod_accum_101__102_, prod_accum_101__101_, prod_accum_101__100_, prod_accum_101__99_, prod_accum_101__98_, prod_accum_101__97_, prod_accum_101__96_, prod_accum_101__95_, prod_accum_101__94_, prod_accum_101__93_, prod_accum_101__92_, prod_accum_101__91_, prod_accum_101__90_, prod_accum_101__89_, prod_accum_101__88_, prod_accum_101__87_, prod_accum_101__86_, prod_accum_101__85_, prod_accum_101__84_, prod_accum_101__83_, prod_accum_101__82_, prod_accum_101__81_, prod_accum_101__80_, prod_accum_101__79_, prod_accum_101__78_, prod_accum_101__77_, prod_accum_101__76_, prod_accum_101__75_, prod_accum_101__74_, prod_accum_101__73_, prod_accum_101__72_, prod_accum_101__71_, prod_accum_101__70_, prod_accum_101__69_, prod_accum_101__68_, prod_accum_101__67_, prod_accum_101__66_, prod_accum_101__65_, prod_accum_101__64_, prod_accum_101__63_, prod_accum_101__62_, prod_accum_101__61_, prod_accum_101__60_, prod_accum_101__59_, prod_accum_101__58_, prod_accum_101__57_, prod_accum_101__56_, prod_accum_101__55_, prod_accum_101__54_, prod_accum_101__53_, prod_accum_101__52_, prod_accum_101__51_, prod_accum_101__50_, prod_accum_101__49_, prod_accum_101__48_, prod_accum_101__47_, prod_accum_101__46_, prod_accum_101__45_, prod_accum_101__44_, prod_accum_101__43_, prod_accum_101__42_, prod_accum_101__41_, prod_accum_101__40_, prod_accum_101__39_, prod_accum_101__38_, prod_accum_101__37_, prod_accum_101__36_, prod_accum_101__35_, prod_accum_101__34_, prod_accum_101__33_, prod_accum_101__32_, prod_accum_101__31_, prod_accum_101__30_, prod_accum_101__29_, prod_accum_101__28_, prod_accum_101__27_, prod_accum_101__26_, prod_accum_101__25_, prod_accum_101__24_, prod_accum_101__23_, prod_accum_101__22_, prod_accum_101__21_, prod_accum_101__20_, prod_accum_101__19_, prod_accum_101__18_, prod_accum_101__17_, prod_accum_101__16_, prod_accum_101__15_, prod_accum_101__14_, prod_accum_101__13_, prod_accum_101__12_, prod_accum_101__11_, prod_accum_101__10_, prod_accum_101__9_, prod_accum_101__8_, prod_accum_101__7_, prod_accum_101__6_, prod_accum_101__5_, prod_accum_101__4_, prod_accum_101__3_, prod_accum_101__2_, prod_accum_101__1_, prod_accum_101__0_ }),
    .a_o(a_r[13183:13056]),
    .b_o(b_r[13183:13056]),
    .s_o({ s_r_102__127_, s_r_102__126_, s_r_102__125_, s_r_102__124_, s_r_102__123_, s_r_102__122_, s_r_102__121_, s_r_102__120_, s_r_102__119_, s_r_102__118_, s_r_102__117_, s_r_102__116_, s_r_102__115_, s_r_102__114_, s_r_102__113_, s_r_102__112_, s_r_102__111_, s_r_102__110_, s_r_102__109_, s_r_102__108_, s_r_102__107_, s_r_102__106_, s_r_102__105_, s_r_102__104_, s_r_102__103_, s_r_102__102_, s_r_102__101_, s_r_102__100_, s_r_102__99_, s_r_102__98_, s_r_102__97_, s_r_102__96_, s_r_102__95_, s_r_102__94_, s_r_102__93_, s_r_102__92_, s_r_102__91_, s_r_102__90_, s_r_102__89_, s_r_102__88_, s_r_102__87_, s_r_102__86_, s_r_102__85_, s_r_102__84_, s_r_102__83_, s_r_102__82_, s_r_102__81_, s_r_102__80_, s_r_102__79_, s_r_102__78_, s_r_102__77_, s_r_102__76_, s_r_102__75_, s_r_102__74_, s_r_102__73_, s_r_102__72_, s_r_102__71_, s_r_102__70_, s_r_102__69_, s_r_102__68_, s_r_102__67_, s_r_102__66_, s_r_102__65_, s_r_102__64_, s_r_102__63_, s_r_102__62_, s_r_102__61_, s_r_102__60_, s_r_102__59_, s_r_102__58_, s_r_102__57_, s_r_102__56_, s_r_102__55_, s_r_102__54_, s_r_102__53_, s_r_102__52_, s_r_102__51_, s_r_102__50_, s_r_102__49_, s_r_102__48_, s_r_102__47_, s_r_102__46_, s_r_102__45_, s_r_102__44_, s_r_102__43_, s_r_102__42_, s_r_102__41_, s_r_102__40_, s_r_102__39_, s_r_102__38_, s_r_102__37_, s_r_102__36_, s_r_102__35_, s_r_102__34_, s_r_102__33_, s_r_102__32_, s_r_102__31_, s_r_102__30_, s_r_102__29_, s_r_102__28_, s_r_102__27_, s_r_102__26_, s_r_102__25_, s_r_102__24_, s_r_102__23_, s_r_102__22_, s_r_102__21_, s_r_102__20_, s_r_102__19_, s_r_102__18_, s_r_102__17_, s_r_102__16_, s_r_102__15_, s_r_102__14_, s_r_102__13_, s_r_102__12_, s_r_102__11_, s_r_102__10_, s_r_102__9_, s_r_102__8_, s_r_102__7_, s_r_102__6_, s_r_102__5_, s_r_102__4_, s_r_102__3_, s_r_102__2_, s_r_102__1_, s_r_102__0_ }),
    .c_o(c_r[102]),
    .prod_accum_o({ prod_accum_102__103_, prod_accum_102__102_, prod_accum_102__101_, prod_accum_102__100_, prod_accum_102__99_, prod_accum_102__98_, prod_accum_102__97_, prod_accum_102__96_, prod_accum_102__95_, prod_accum_102__94_, prod_accum_102__93_, prod_accum_102__92_, prod_accum_102__91_, prod_accum_102__90_, prod_accum_102__89_, prod_accum_102__88_, prod_accum_102__87_, prod_accum_102__86_, prod_accum_102__85_, prod_accum_102__84_, prod_accum_102__83_, prod_accum_102__82_, prod_accum_102__81_, prod_accum_102__80_, prod_accum_102__79_, prod_accum_102__78_, prod_accum_102__77_, prod_accum_102__76_, prod_accum_102__75_, prod_accum_102__74_, prod_accum_102__73_, prod_accum_102__72_, prod_accum_102__71_, prod_accum_102__70_, prod_accum_102__69_, prod_accum_102__68_, prod_accum_102__67_, prod_accum_102__66_, prod_accum_102__65_, prod_accum_102__64_, prod_accum_102__63_, prod_accum_102__62_, prod_accum_102__61_, prod_accum_102__60_, prod_accum_102__59_, prod_accum_102__58_, prod_accum_102__57_, prod_accum_102__56_, prod_accum_102__55_, prod_accum_102__54_, prod_accum_102__53_, prod_accum_102__52_, prod_accum_102__51_, prod_accum_102__50_, prod_accum_102__49_, prod_accum_102__48_, prod_accum_102__47_, prod_accum_102__46_, prod_accum_102__45_, prod_accum_102__44_, prod_accum_102__43_, prod_accum_102__42_, prod_accum_102__41_, prod_accum_102__40_, prod_accum_102__39_, prod_accum_102__38_, prod_accum_102__37_, prod_accum_102__36_, prod_accum_102__35_, prod_accum_102__34_, prod_accum_102__33_, prod_accum_102__32_, prod_accum_102__31_, prod_accum_102__30_, prod_accum_102__29_, prod_accum_102__28_, prod_accum_102__27_, prod_accum_102__26_, prod_accum_102__25_, prod_accum_102__24_, prod_accum_102__23_, prod_accum_102__22_, prod_accum_102__21_, prod_accum_102__20_, prod_accum_102__19_, prod_accum_102__18_, prod_accum_102__17_, prod_accum_102__16_, prod_accum_102__15_, prod_accum_102__14_, prod_accum_102__13_, prod_accum_102__12_, prod_accum_102__11_, prod_accum_102__10_, prod_accum_102__9_, prod_accum_102__8_, prod_accum_102__7_, prod_accum_102__6_, prod_accum_102__5_, prod_accum_102__4_, prod_accum_102__3_, prod_accum_102__2_, prod_accum_102__1_, prod_accum_102__0_ })
  );


  bsg_mul_array_row_128_103_x
  genblk1_103__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[13183:13056]),
    .b_i(b_r[13183:13056]),
    .s_i({ s_r_102__127_, s_r_102__126_, s_r_102__125_, s_r_102__124_, s_r_102__123_, s_r_102__122_, s_r_102__121_, s_r_102__120_, s_r_102__119_, s_r_102__118_, s_r_102__117_, s_r_102__116_, s_r_102__115_, s_r_102__114_, s_r_102__113_, s_r_102__112_, s_r_102__111_, s_r_102__110_, s_r_102__109_, s_r_102__108_, s_r_102__107_, s_r_102__106_, s_r_102__105_, s_r_102__104_, s_r_102__103_, s_r_102__102_, s_r_102__101_, s_r_102__100_, s_r_102__99_, s_r_102__98_, s_r_102__97_, s_r_102__96_, s_r_102__95_, s_r_102__94_, s_r_102__93_, s_r_102__92_, s_r_102__91_, s_r_102__90_, s_r_102__89_, s_r_102__88_, s_r_102__87_, s_r_102__86_, s_r_102__85_, s_r_102__84_, s_r_102__83_, s_r_102__82_, s_r_102__81_, s_r_102__80_, s_r_102__79_, s_r_102__78_, s_r_102__77_, s_r_102__76_, s_r_102__75_, s_r_102__74_, s_r_102__73_, s_r_102__72_, s_r_102__71_, s_r_102__70_, s_r_102__69_, s_r_102__68_, s_r_102__67_, s_r_102__66_, s_r_102__65_, s_r_102__64_, s_r_102__63_, s_r_102__62_, s_r_102__61_, s_r_102__60_, s_r_102__59_, s_r_102__58_, s_r_102__57_, s_r_102__56_, s_r_102__55_, s_r_102__54_, s_r_102__53_, s_r_102__52_, s_r_102__51_, s_r_102__50_, s_r_102__49_, s_r_102__48_, s_r_102__47_, s_r_102__46_, s_r_102__45_, s_r_102__44_, s_r_102__43_, s_r_102__42_, s_r_102__41_, s_r_102__40_, s_r_102__39_, s_r_102__38_, s_r_102__37_, s_r_102__36_, s_r_102__35_, s_r_102__34_, s_r_102__33_, s_r_102__32_, s_r_102__31_, s_r_102__30_, s_r_102__29_, s_r_102__28_, s_r_102__27_, s_r_102__26_, s_r_102__25_, s_r_102__24_, s_r_102__23_, s_r_102__22_, s_r_102__21_, s_r_102__20_, s_r_102__19_, s_r_102__18_, s_r_102__17_, s_r_102__16_, s_r_102__15_, s_r_102__14_, s_r_102__13_, s_r_102__12_, s_r_102__11_, s_r_102__10_, s_r_102__9_, s_r_102__8_, s_r_102__7_, s_r_102__6_, s_r_102__5_, s_r_102__4_, s_r_102__3_, s_r_102__2_, s_r_102__1_, s_r_102__0_ }),
    .c_i(c_r[102]),
    .prod_accum_i({ prod_accum_102__103_, prod_accum_102__102_, prod_accum_102__101_, prod_accum_102__100_, prod_accum_102__99_, prod_accum_102__98_, prod_accum_102__97_, prod_accum_102__96_, prod_accum_102__95_, prod_accum_102__94_, prod_accum_102__93_, prod_accum_102__92_, prod_accum_102__91_, prod_accum_102__90_, prod_accum_102__89_, prod_accum_102__88_, prod_accum_102__87_, prod_accum_102__86_, prod_accum_102__85_, prod_accum_102__84_, prod_accum_102__83_, prod_accum_102__82_, prod_accum_102__81_, prod_accum_102__80_, prod_accum_102__79_, prod_accum_102__78_, prod_accum_102__77_, prod_accum_102__76_, prod_accum_102__75_, prod_accum_102__74_, prod_accum_102__73_, prod_accum_102__72_, prod_accum_102__71_, prod_accum_102__70_, prod_accum_102__69_, prod_accum_102__68_, prod_accum_102__67_, prod_accum_102__66_, prod_accum_102__65_, prod_accum_102__64_, prod_accum_102__63_, prod_accum_102__62_, prod_accum_102__61_, prod_accum_102__60_, prod_accum_102__59_, prod_accum_102__58_, prod_accum_102__57_, prod_accum_102__56_, prod_accum_102__55_, prod_accum_102__54_, prod_accum_102__53_, prod_accum_102__52_, prod_accum_102__51_, prod_accum_102__50_, prod_accum_102__49_, prod_accum_102__48_, prod_accum_102__47_, prod_accum_102__46_, prod_accum_102__45_, prod_accum_102__44_, prod_accum_102__43_, prod_accum_102__42_, prod_accum_102__41_, prod_accum_102__40_, prod_accum_102__39_, prod_accum_102__38_, prod_accum_102__37_, prod_accum_102__36_, prod_accum_102__35_, prod_accum_102__34_, prod_accum_102__33_, prod_accum_102__32_, prod_accum_102__31_, prod_accum_102__30_, prod_accum_102__29_, prod_accum_102__28_, prod_accum_102__27_, prod_accum_102__26_, prod_accum_102__25_, prod_accum_102__24_, prod_accum_102__23_, prod_accum_102__22_, prod_accum_102__21_, prod_accum_102__20_, prod_accum_102__19_, prod_accum_102__18_, prod_accum_102__17_, prod_accum_102__16_, prod_accum_102__15_, prod_accum_102__14_, prod_accum_102__13_, prod_accum_102__12_, prod_accum_102__11_, prod_accum_102__10_, prod_accum_102__9_, prod_accum_102__8_, prod_accum_102__7_, prod_accum_102__6_, prod_accum_102__5_, prod_accum_102__4_, prod_accum_102__3_, prod_accum_102__2_, prod_accum_102__1_, prod_accum_102__0_ }),
    .a_o(a_r[13311:13184]),
    .b_o(b_r[13311:13184]),
    .s_o({ s_r_103__127_, s_r_103__126_, s_r_103__125_, s_r_103__124_, s_r_103__123_, s_r_103__122_, s_r_103__121_, s_r_103__120_, s_r_103__119_, s_r_103__118_, s_r_103__117_, s_r_103__116_, s_r_103__115_, s_r_103__114_, s_r_103__113_, s_r_103__112_, s_r_103__111_, s_r_103__110_, s_r_103__109_, s_r_103__108_, s_r_103__107_, s_r_103__106_, s_r_103__105_, s_r_103__104_, s_r_103__103_, s_r_103__102_, s_r_103__101_, s_r_103__100_, s_r_103__99_, s_r_103__98_, s_r_103__97_, s_r_103__96_, s_r_103__95_, s_r_103__94_, s_r_103__93_, s_r_103__92_, s_r_103__91_, s_r_103__90_, s_r_103__89_, s_r_103__88_, s_r_103__87_, s_r_103__86_, s_r_103__85_, s_r_103__84_, s_r_103__83_, s_r_103__82_, s_r_103__81_, s_r_103__80_, s_r_103__79_, s_r_103__78_, s_r_103__77_, s_r_103__76_, s_r_103__75_, s_r_103__74_, s_r_103__73_, s_r_103__72_, s_r_103__71_, s_r_103__70_, s_r_103__69_, s_r_103__68_, s_r_103__67_, s_r_103__66_, s_r_103__65_, s_r_103__64_, s_r_103__63_, s_r_103__62_, s_r_103__61_, s_r_103__60_, s_r_103__59_, s_r_103__58_, s_r_103__57_, s_r_103__56_, s_r_103__55_, s_r_103__54_, s_r_103__53_, s_r_103__52_, s_r_103__51_, s_r_103__50_, s_r_103__49_, s_r_103__48_, s_r_103__47_, s_r_103__46_, s_r_103__45_, s_r_103__44_, s_r_103__43_, s_r_103__42_, s_r_103__41_, s_r_103__40_, s_r_103__39_, s_r_103__38_, s_r_103__37_, s_r_103__36_, s_r_103__35_, s_r_103__34_, s_r_103__33_, s_r_103__32_, s_r_103__31_, s_r_103__30_, s_r_103__29_, s_r_103__28_, s_r_103__27_, s_r_103__26_, s_r_103__25_, s_r_103__24_, s_r_103__23_, s_r_103__22_, s_r_103__21_, s_r_103__20_, s_r_103__19_, s_r_103__18_, s_r_103__17_, s_r_103__16_, s_r_103__15_, s_r_103__14_, s_r_103__13_, s_r_103__12_, s_r_103__11_, s_r_103__10_, s_r_103__9_, s_r_103__8_, s_r_103__7_, s_r_103__6_, s_r_103__5_, s_r_103__4_, s_r_103__3_, s_r_103__2_, s_r_103__1_, s_r_103__0_ }),
    .c_o(c_r[103]),
    .prod_accum_o({ prod_accum_103__104_, prod_accum_103__103_, prod_accum_103__102_, prod_accum_103__101_, prod_accum_103__100_, prod_accum_103__99_, prod_accum_103__98_, prod_accum_103__97_, prod_accum_103__96_, prod_accum_103__95_, prod_accum_103__94_, prod_accum_103__93_, prod_accum_103__92_, prod_accum_103__91_, prod_accum_103__90_, prod_accum_103__89_, prod_accum_103__88_, prod_accum_103__87_, prod_accum_103__86_, prod_accum_103__85_, prod_accum_103__84_, prod_accum_103__83_, prod_accum_103__82_, prod_accum_103__81_, prod_accum_103__80_, prod_accum_103__79_, prod_accum_103__78_, prod_accum_103__77_, prod_accum_103__76_, prod_accum_103__75_, prod_accum_103__74_, prod_accum_103__73_, prod_accum_103__72_, prod_accum_103__71_, prod_accum_103__70_, prod_accum_103__69_, prod_accum_103__68_, prod_accum_103__67_, prod_accum_103__66_, prod_accum_103__65_, prod_accum_103__64_, prod_accum_103__63_, prod_accum_103__62_, prod_accum_103__61_, prod_accum_103__60_, prod_accum_103__59_, prod_accum_103__58_, prod_accum_103__57_, prod_accum_103__56_, prod_accum_103__55_, prod_accum_103__54_, prod_accum_103__53_, prod_accum_103__52_, prod_accum_103__51_, prod_accum_103__50_, prod_accum_103__49_, prod_accum_103__48_, prod_accum_103__47_, prod_accum_103__46_, prod_accum_103__45_, prod_accum_103__44_, prod_accum_103__43_, prod_accum_103__42_, prod_accum_103__41_, prod_accum_103__40_, prod_accum_103__39_, prod_accum_103__38_, prod_accum_103__37_, prod_accum_103__36_, prod_accum_103__35_, prod_accum_103__34_, prod_accum_103__33_, prod_accum_103__32_, prod_accum_103__31_, prod_accum_103__30_, prod_accum_103__29_, prod_accum_103__28_, prod_accum_103__27_, prod_accum_103__26_, prod_accum_103__25_, prod_accum_103__24_, prod_accum_103__23_, prod_accum_103__22_, prod_accum_103__21_, prod_accum_103__20_, prod_accum_103__19_, prod_accum_103__18_, prod_accum_103__17_, prod_accum_103__16_, prod_accum_103__15_, prod_accum_103__14_, prod_accum_103__13_, prod_accum_103__12_, prod_accum_103__11_, prod_accum_103__10_, prod_accum_103__9_, prod_accum_103__8_, prod_accum_103__7_, prod_accum_103__6_, prod_accum_103__5_, prod_accum_103__4_, prod_accum_103__3_, prod_accum_103__2_, prod_accum_103__1_, prod_accum_103__0_ })
  );


  bsg_mul_array_row_128_104_x
  genblk1_104__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[13311:13184]),
    .b_i(b_r[13311:13184]),
    .s_i({ s_r_103__127_, s_r_103__126_, s_r_103__125_, s_r_103__124_, s_r_103__123_, s_r_103__122_, s_r_103__121_, s_r_103__120_, s_r_103__119_, s_r_103__118_, s_r_103__117_, s_r_103__116_, s_r_103__115_, s_r_103__114_, s_r_103__113_, s_r_103__112_, s_r_103__111_, s_r_103__110_, s_r_103__109_, s_r_103__108_, s_r_103__107_, s_r_103__106_, s_r_103__105_, s_r_103__104_, s_r_103__103_, s_r_103__102_, s_r_103__101_, s_r_103__100_, s_r_103__99_, s_r_103__98_, s_r_103__97_, s_r_103__96_, s_r_103__95_, s_r_103__94_, s_r_103__93_, s_r_103__92_, s_r_103__91_, s_r_103__90_, s_r_103__89_, s_r_103__88_, s_r_103__87_, s_r_103__86_, s_r_103__85_, s_r_103__84_, s_r_103__83_, s_r_103__82_, s_r_103__81_, s_r_103__80_, s_r_103__79_, s_r_103__78_, s_r_103__77_, s_r_103__76_, s_r_103__75_, s_r_103__74_, s_r_103__73_, s_r_103__72_, s_r_103__71_, s_r_103__70_, s_r_103__69_, s_r_103__68_, s_r_103__67_, s_r_103__66_, s_r_103__65_, s_r_103__64_, s_r_103__63_, s_r_103__62_, s_r_103__61_, s_r_103__60_, s_r_103__59_, s_r_103__58_, s_r_103__57_, s_r_103__56_, s_r_103__55_, s_r_103__54_, s_r_103__53_, s_r_103__52_, s_r_103__51_, s_r_103__50_, s_r_103__49_, s_r_103__48_, s_r_103__47_, s_r_103__46_, s_r_103__45_, s_r_103__44_, s_r_103__43_, s_r_103__42_, s_r_103__41_, s_r_103__40_, s_r_103__39_, s_r_103__38_, s_r_103__37_, s_r_103__36_, s_r_103__35_, s_r_103__34_, s_r_103__33_, s_r_103__32_, s_r_103__31_, s_r_103__30_, s_r_103__29_, s_r_103__28_, s_r_103__27_, s_r_103__26_, s_r_103__25_, s_r_103__24_, s_r_103__23_, s_r_103__22_, s_r_103__21_, s_r_103__20_, s_r_103__19_, s_r_103__18_, s_r_103__17_, s_r_103__16_, s_r_103__15_, s_r_103__14_, s_r_103__13_, s_r_103__12_, s_r_103__11_, s_r_103__10_, s_r_103__9_, s_r_103__8_, s_r_103__7_, s_r_103__6_, s_r_103__5_, s_r_103__4_, s_r_103__3_, s_r_103__2_, s_r_103__1_, s_r_103__0_ }),
    .c_i(c_r[103]),
    .prod_accum_i({ prod_accum_103__104_, prod_accum_103__103_, prod_accum_103__102_, prod_accum_103__101_, prod_accum_103__100_, prod_accum_103__99_, prod_accum_103__98_, prod_accum_103__97_, prod_accum_103__96_, prod_accum_103__95_, prod_accum_103__94_, prod_accum_103__93_, prod_accum_103__92_, prod_accum_103__91_, prod_accum_103__90_, prod_accum_103__89_, prod_accum_103__88_, prod_accum_103__87_, prod_accum_103__86_, prod_accum_103__85_, prod_accum_103__84_, prod_accum_103__83_, prod_accum_103__82_, prod_accum_103__81_, prod_accum_103__80_, prod_accum_103__79_, prod_accum_103__78_, prod_accum_103__77_, prod_accum_103__76_, prod_accum_103__75_, prod_accum_103__74_, prod_accum_103__73_, prod_accum_103__72_, prod_accum_103__71_, prod_accum_103__70_, prod_accum_103__69_, prod_accum_103__68_, prod_accum_103__67_, prod_accum_103__66_, prod_accum_103__65_, prod_accum_103__64_, prod_accum_103__63_, prod_accum_103__62_, prod_accum_103__61_, prod_accum_103__60_, prod_accum_103__59_, prod_accum_103__58_, prod_accum_103__57_, prod_accum_103__56_, prod_accum_103__55_, prod_accum_103__54_, prod_accum_103__53_, prod_accum_103__52_, prod_accum_103__51_, prod_accum_103__50_, prod_accum_103__49_, prod_accum_103__48_, prod_accum_103__47_, prod_accum_103__46_, prod_accum_103__45_, prod_accum_103__44_, prod_accum_103__43_, prod_accum_103__42_, prod_accum_103__41_, prod_accum_103__40_, prod_accum_103__39_, prod_accum_103__38_, prod_accum_103__37_, prod_accum_103__36_, prod_accum_103__35_, prod_accum_103__34_, prod_accum_103__33_, prod_accum_103__32_, prod_accum_103__31_, prod_accum_103__30_, prod_accum_103__29_, prod_accum_103__28_, prod_accum_103__27_, prod_accum_103__26_, prod_accum_103__25_, prod_accum_103__24_, prod_accum_103__23_, prod_accum_103__22_, prod_accum_103__21_, prod_accum_103__20_, prod_accum_103__19_, prod_accum_103__18_, prod_accum_103__17_, prod_accum_103__16_, prod_accum_103__15_, prod_accum_103__14_, prod_accum_103__13_, prod_accum_103__12_, prod_accum_103__11_, prod_accum_103__10_, prod_accum_103__9_, prod_accum_103__8_, prod_accum_103__7_, prod_accum_103__6_, prod_accum_103__5_, prod_accum_103__4_, prod_accum_103__3_, prod_accum_103__2_, prod_accum_103__1_, prod_accum_103__0_ }),
    .a_o(a_r[13439:13312]),
    .b_o(b_r[13439:13312]),
    .s_o({ s_r_104__127_, s_r_104__126_, s_r_104__125_, s_r_104__124_, s_r_104__123_, s_r_104__122_, s_r_104__121_, s_r_104__120_, s_r_104__119_, s_r_104__118_, s_r_104__117_, s_r_104__116_, s_r_104__115_, s_r_104__114_, s_r_104__113_, s_r_104__112_, s_r_104__111_, s_r_104__110_, s_r_104__109_, s_r_104__108_, s_r_104__107_, s_r_104__106_, s_r_104__105_, s_r_104__104_, s_r_104__103_, s_r_104__102_, s_r_104__101_, s_r_104__100_, s_r_104__99_, s_r_104__98_, s_r_104__97_, s_r_104__96_, s_r_104__95_, s_r_104__94_, s_r_104__93_, s_r_104__92_, s_r_104__91_, s_r_104__90_, s_r_104__89_, s_r_104__88_, s_r_104__87_, s_r_104__86_, s_r_104__85_, s_r_104__84_, s_r_104__83_, s_r_104__82_, s_r_104__81_, s_r_104__80_, s_r_104__79_, s_r_104__78_, s_r_104__77_, s_r_104__76_, s_r_104__75_, s_r_104__74_, s_r_104__73_, s_r_104__72_, s_r_104__71_, s_r_104__70_, s_r_104__69_, s_r_104__68_, s_r_104__67_, s_r_104__66_, s_r_104__65_, s_r_104__64_, s_r_104__63_, s_r_104__62_, s_r_104__61_, s_r_104__60_, s_r_104__59_, s_r_104__58_, s_r_104__57_, s_r_104__56_, s_r_104__55_, s_r_104__54_, s_r_104__53_, s_r_104__52_, s_r_104__51_, s_r_104__50_, s_r_104__49_, s_r_104__48_, s_r_104__47_, s_r_104__46_, s_r_104__45_, s_r_104__44_, s_r_104__43_, s_r_104__42_, s_r_104__41_, s_r_104__40_, s_r_104__39_, s_r_104__38_, s_r_104__37_, s_r_104__36_, s_r_104__35_, s_r_104__34_, s_r_104__33_, s_r_104__32_, s_r_104__31_, s_r_104__30_, s_r_104__29_, s_r_104__28_, s_r_104__27_, s_r_104__26_, s_r_104__25_, s_r_104__24_, s_r_104__23_, s_r_104__22_, s_r_104__21_, s_r_104__20_, s_r_104__19_, s_r_104__18_, s_r_104__17_, s_r_104__16_, s_r_104__15_, s_r_104__14_, s_r_104__13_, s_r_104__12_, s_r_104__11_, s_r_104__10_, s_r_104__9_, s_r_104__8_, s_r_104__7_, s_r_104__6_, s_r_104__5_, s_r_104__4_, s_r_104__3_, s_r_104__2_, s_r_104__1_, s_r_104__0_ }),
    .c_o(c_r[104]),
    .prod_accum_o({ prod_accum_104__105_, prod_accum_104__104_, prod_accum_104__103_, prod_accum_104__102_, prod_accum_104__101_, prod_accum_104__100_, prod_accum_104__99_, prod_accum_104__98_, prod_accum_104__97_, prod_accum_104__96_, prod_accum_104__95_, prod_accum_104__94_, prod_accum_104__93_, prod_accum_104__92_, prod_accum_104__91_, prod_accum_104__90_, prod_accum_104__89_, prod_accum_104__88_, prod_accum_104__87_, prod_accum_104__86_, prod_accum_104__85_, prod_accum_104__84_, prod_accum_104__83_, prod_accum_104__82_, prod_accum_104__81_, prod_accum_104__80_, prod_accum_104__79_, prod_accum_104__78_, prod_accum_104__77_, prod_accum_104__76_, prod_accum_104__75_, prod_accum_104__74_, prod_accum_104__73_, prod_accum_104__72_, prod_accum_104__71_, prod_accum_104__70_, prod_accum_104__69_, prod_accum_104__68_, prod_accum_104__67_, prod_accum_104__66_, prod_accum_104__65_, prod_accum_104__64_, prod_accum_104__63_, prod_accum_104__62_, prod_accum_104__61_, prod_accum_104__60_, prod_accum_104__59_, prod_accum_104__58_, prod_accum_104__57_, prod_accum_104__56_, prod_accum_104__55_, prod_accum_104__54_, prod_accum_104__53_, prod_accum_104__52_, prod_accum_104__51_, prod_accum_104__50_, prod_accum_104__49_, prod_accum_104__48_, prod_accum_104__47_, prod_accum_104__46_, prod_accum_104__45_, prod_accum_104__44_, prod_accum_104__43_, prod_accum_104__42_, prod_accum_104__41_, prod_accum_104__40_, prod_accum_104__39_, prod_accum_104__38_, prod_accum_104__37_, prod_accum_104__36_, prod_accum_104__35_, prod_accum_104__34_, prod_accum_104__33_, prod_accum_104__32_, prod_accum_104__31_, prod_accum_104__30_, prod_accum_104__29_, prod_accum_104__28_, prod_accum_104__27_, prod_accum_104__26_, prod_accum_104__25_, prod_accum_104__24_, prod_accum_104__23_, prod_accum_104__22_, prod_accum_104__21_, prod_accum_104__20_, prod_accum_104__19_, prod_accum_104__18_, prod_accum_104__17_, prod_accum_104__16_, prod_accum_104__15_, prod_accum_104__14_, prod_accum_104__13_, prod_accum_104__12_, prod_accum_104__11_, prod_accum_104__10_, prod_accum_104__9_, prod_accum_104__8_, prod_accum_104__7_, prod_accum_104__6_, prod_accum_104__5_, prod_accum_104__4_, prod_accum_104__3_, prod_accum_104__2_, prod_accum_104__1_, prod_accum_104__0_ })
  );


  bsg_mul_array_row_128_105_x
  genblk1_105__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[13439:13312]),
    .b_i(b_r[13439:13312]),
    .s_i({ s_r_104__127_, s_r_104__126_, s_r_104__125_, s_r_104__124_, s_r_104__123_, s_r_104__122_, s_r_104__121_, s_r_104__120_, s_r_104__119_, s_r_104__118_, s_r_104__117_, s_r_104__116_, s_r_104__115_, s_r_104__114_, s_r_104__113_, s_r_104__112_, s_r_104__111_, s_r_104__110_, s_r_104__109_, s_r_104__108_, s_r_104__107_, s_r_104__106_, s_r_104__105_, s_r_104__104_, s_r_104__103_, s_r_104__102_, s_r_104__101_, s_r_104__100_, s_r_104__99_, s_r_104__98_, s_r_104__97_, s_r_104__96_, s_r_104__95_, s_r_104__94_, s_r_104__93_, s_r_104__92_, s_r_104__91_, s_r_104__90_, s_r_104__89_, s_r_104__88_, s_r_104__87_, s_r_104__86_, s_r_104__85_, s_r_104__84_, s_r_104__83_, s_r_104__82_, s_r_104__81_, s_r_104__80_, s_r_104__79_, s_r_104__78_, s_r_104__77_, s_r_104__76_, s_r_104__75_, s_r_104__74_, s_r_104__73_, s_r_104__72_, s_r_104__71_, s_r_104__70_, s_r_104__69_, s_r_104__68_, s_r_104__67_, s_r_104__66_, s_r_104__65_, s_r_104__64_, s_r_104__63_, s_r_104__62_, s_r_104__61_, s_r_104__60_, s_r_104__59_, s_r_104__58_, s_r_104__57_, s_r_104__56_, s_r_104__55_, s_r_104__54_, s_r_104__53_, s_r_104__52_, s_r_104__51_, s_r_104__50_, s_r_104__49_, s_r_104__48_, s_r_104__47_, s_r_104__46_, s_r_104__45_, s_r_104__44_, s_r_104__43_, s_r_104__42_, s_r_104__41_, s_r_104__40_, s_r_104__39_, s_r_104__38_, s_r_104__37_, s_r_104__36_, s_r_104__35_, s_r_104__34_, s_r_104__33_, s_r_104__32_, s_r_104__31_, s_r_104__30_, s_r_104__29_, s_r_104__28_, s_r_104__27_, s_r_104__26_, s_r_104__25_, s_r_104__24_, s_r_104__23_, s_r_104__22_, s_r_104__21_, s_r_104__20_, s_r_104__19_, s_r_104__18_, s_r_104__17_, s_r_104__16_, s_r_104__15_, s_r_104__14_, s_r_104__13_, s_r_104__12_, s_r_104__11_, s_r_104__10_, s_r_104__9_, s_r_104__8_, s_r_104__7_, s_r_104__6_, s_r_104__5_, s_r_104__4_, s_r_104__3_, s_r_104__2_, s_r_104__1_, s_r_104__0_ }),
    .c_i(c_r[104]),
    .prod_accum_i({ prod_accum_104__105_, prod_accum_104__104_, prod_accum_104__103_, prod_accum_104__102_, prod_accum_104__101_, prod_accum_104__100_, prod_accum_104__99_, prod_accum_104__98_, prod_accum_104__97_, prod_accum_104__96_, prod_accum_104__95_, prod_accum_104__94_, prod_accum_104__93_, prod_accum_104__92_, prod_accum_104__91_, prod_accum_104__90_, prod_accum_104__89_, prod_accum_104__88_, prod_accum_104__87_, prod_accum_104__86_, prod_accum_104__85_, prod_accum_104__84_, prod_accum_104__83_, prod_accum_104__82_, prod_accum_104__81_, prod_accum_104__80_, prod_accum_104__79_, prod_accum_104__78_, prod_accum_104__77_, prod_accum_104__76_, prod_accum_104__75_, prod_accum_104__74_, prod_accum_104__73_, prod_accum_104__72_, prod_accum_104__71_, prod_accum_104__70_, prod_accum_104__69_, prod_accum_104__68_, prod_accum_104__67_, prod_accum_104__66_, prod_accum_104__65_, prod_accum_104__64_, prod_accum_104__63_, prod_accum_104__62_, prod_accum_104__61_, prod_accum_104__60_, prod_accum_104__59_, prod_accum_104__58_, prod_accum_104__57_, prod_accum_104__56_, prod_accum_104__55_, prod_accum_104__54_, prod_accum_104__53_, prod_accum_104__52_, prod_accum_104__51_, prod_accum_104__50_, prod_accum_104__49_, prod_accum_104__48_, prod_accum_104__47_, prod_accum_104__46_, prod_accum_104__45_, prod_accum_104__44_, prod_accum_104__43_, prod_accum_104__42_, prod_accum_104__41_, prod_accum_104__40_, prod_accum_104__39_, prod_accum_104__38_, prod_accum_104__37_, prod_accum_104__36_, prod_accum_104__35_, prod_accum_104__34_, prod_accum_104__33_, prod_accum_104__32_, prod_accum_104__31_, prod_accum_104__30_, prod_accum_104__29_, prod_accum_104__28_, prod_accum_104__27_, prod_accum_104__26_, prod_accum_104__25_, prod_accum_104__24_, prod_accum_104__23_, prod_accum_104__22_, prod_accum_104__21_, prod_accum_104__20_, prod_accum_104__19_, prod_accum_104__18_, prod_accum_104__17_, prod_accum_104__16_, prod_accum_104__15_, prod_accum_104__14_, prod_accum_104__13_, prod_accum_104__12_, prod_accum_104__11_, prod_accum_104__10_, prod_accum_104__9_, prod_accum_104__8_, prod_accum_104__7_, prod_accum_104__6_, prod_accum_104__5_, prod_accum_104__4_, prod_accum_104__3_, prod_accum_104__2_, prod_accum_104__1_, prod_accum_104__0_ }),
    .a_o(a_r[13567:13440]),
    .b_o(b_r[13567:13440]),
    .s_o({ s_r_105__127_, s_r_105__126_, s_r_105__125_, s_r_105__124_, s_r_105__123_, s_r_105__122_, s_r_105__121_, s_r_105__120_, s_r_105__119_, s_r_105__118_, s_r_105__117_, s_r_105__116_, s_r_105__115_, s_r_105__114_, s_r_105__113_, s_r_105__112_, s_r_105__111_, s_r_105__110_, s_r_105__109_, s_r_105__108_, s_r_105__107_, s_r_105__106_, s_r_105__105_, s_r_105__104_, s_r_105__103_, s_r_105__102_, s_r_105__101_, s_r_105__100_, s_r_105__99_, s_r_105__98_, s_r_105__97_, s_r_105__96_, s_r_105__95_, s_r_105__94_, s_r_105__93_, s_r_105__92_, s_r_105__91_, s_r_105__90_, s_r_105__89_, s_r_105__88_, s_r_105__87_, s_r_105__86_, s_r_105__85_, s_r_105__84_, s_r_105__83_, s_r_105__82_, s_r_105__81_, s_r_105__80_, s_r_105__79_, s_r_105__78_, s_r_105__77_, s_r_105__76_, s_r_105__75_, s_r_105__74_, s_r_105__73_, s_r_105__72_, s_r_105__71_, s_r_105__70_, s_r_105__69_, s_r_105__68_, s_r_105__67_, s_r_105__66_, s_r_105__65_, s_r_105__64_, s_r_105__63_, s_r_105__62_, s_r_105__61_, s_r_105__60_, s_r_105__59_, s_r_105__58_, s_r_105__57_, s_r_105__56_, s_r_105__55_, s_r_105__54_, s_r_105__53_, s_r_105__52_, s_r_105__51_, s_r_105__50_, s_r_105__49_, s_r_105__48_, s_r_105__47_, s_r_105__46_, s_r_105__45_, s_r_105__44_, s_r_105__43_, s_r_105__42_, s_r_105__41_, s_r_105__40_, s_r_105__39_, s_r_105__38_, s_r_105__37_, s_r_105__36_, s_r_105__35_, s_r_105__34_, s_r_105__33_, s_r_105__32_, s_r_105__31_, s_r_105__30_, s_r_105__29_, s_r_105__28_, s_r_105__27_, s_r_105__26_, s_r_105__25_, s_r_105__24_, s_r_105__23_, s_r_105__22_, s_r_105__21_, s_r_105__20_, s_r_105__19_, s_r_105__18_, s_r_105__17_, s_r_105__16_, s_r_105__15_, s_r_105__14_, s_r_105__13_, s_r_105__12_, s_r_105__11_, s_r_105__10_, s_r_105__9_, s_r_105__8_, s_r_105__7_, s_r_105__6_, s_r_105__5_, s_r_105__4_, s_r_105__3_, s_r_105__2_, s_r_105__1_, s_r_105__0_ }),
    .c_o(c_r[105]),
    .prod_accum_o({ prod_accum_105__106_, prod_accum_105__105_, prod_accum_105__104_, prod_accum_105__103_, prod_accum_105__102_, prod_accum_105__101_, prod_accum_105__100_, prod_accum_105__99_, prod_accum_105__98_, prod_accum_105__97_, prod_accum_105__96_, prod_accum_105__95_, prod_accum_105__94_, prod_accum_105__93_, prod_accum_105__92_, prod_accum_105__91_, prod_accum_105__90_, prod_accum_105__89_, prod_accum_105__88_, prod_accum_105__87_, prod_accum_105__86_, prod_accum_105__85_, prod_accum_105__84_, prod_accum_105__83_, prod_accum_105__82_, prod_accum_105__81_, prod_accum_105__80_, prod_accum_105__79_, prod_accum_105__78_, prod_accum_105__77_, prod_accum_105__76_, prod_accum_105__75_, prod_accum_105__74_, prod_accum_105__73_, prod_accum_105__72_, prod_accum_105__71_, prod_accum_105__70_, prod_accum_105__69_, prod_accum_105__68_, prod_accum_105__67_, prod_accum_105__66_, prod_accum_105__65_, prod_accum_105__64_, prod_accum_105__63_, prod_accum_105__62_, prod_accum_105__61_, prod_accum_105__60_, prod_accum_105__59_, prod_accum_105__58_, prod_accum_105__57_, prod_accum_105__56_, prod_accum_105__55_, prod_accum_105__54_, prod_accum_105__53_, prod_accum_105__52_, prod_accum_105__51_, prod_accum_105__50_, prod_accum_105__49_, prod_accum_105__48_, prod_accum_105__47_, prod_accum_105__46_, prod_accum_105__45_, prod_accum_105__44_, prod_accum_105__43_, prod_accum_105__42_, prod_accum_105__41_, prod_accum_105__40_, prod_accum_105__39_, prod_accum_105__38_, prod_accum_105__37_, prod_accum_105__36_, prod_accum_105__35_, prod_accum_105__34_, prod_accum_105__33_, prod_accum_105__32_, prod_accum_105__31_, prod_accum_105__30_, prod_accum_105__29_, prod_accum_105__28_, prod_accum_105__27_, prod_accum_105__26_, prod_accum_105__25_, prod_accum_105__24_, prod_accum_105__23_, prod_accum_105__22_, prod_accum_105__21_, prod_accum_105__20_, prod_accum_105__19_, prod_accum_105__18_, prod_accum_105__17_, prod_accum_105__16_, prod_accum_105__15_, prod_accum_105__14_, prod_accum_105__13_, prod_accum_105__12_, prod_accum_105__11_, prod_accum_105__10_, prod_accum_105__9_, prod_accum_105__8_, prod_accum_105__7_, prod_accum_105__6_, prod_accum_105__5_, prod_accum_105__4_, prod_accum_105__3_, prod_accum_105__2_, prod_accum_105__1_, prod_accum_105__0_ })
  );


  bsg_mul_array_row_128_106_x
  genblk1_106__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[13567:13440]),
    .b_i(b_r[13567:13440]),
    .s_i({ s_r_105__127_, s_r_105__126_, s_r_105__125_, s_r_105__124_, s_r_105__123_, s_r_105__122_, s_r_105__121_, s_r_105__120_, s_r_105__119_, s_r_105__118_, s_r_105__117_, s_r_105__116_, s_r_105__115_, s_r_105__114_, s_r_105__113_, s_r_105__112_, s_r_105__111_, s_r_105__110_, s_r_105__109_, s_r_105__108_, s_r_105__107_, s_r_105__106_, s_r_105__105_, s_r_105__104_, s_r_105__103_, s_r_105__102_, s_r_105__101_, s_r_105__100_, s_r_105__99_, s_r_105__98_, s_r_105__97_, s_r_105__96_, s_r_105__95_, s_r_105__94_, s_r_105__93_, s_r_105__92_, s_r_105__91_, s_r_105__90_, s_r_105__89_, s_r_105__88_, s_r_105__87_, s_r_105__86_, s_r_105__85_, s_r_105__84_, s_r_105__83_, s_r_105__82_, s_r_105__81_, s_r_105__80_, s_r_105__79_, s_r_105__78_, s_r_105__77_, s_r_105__76_, s_r_105__75_, s_r_105__74_, s_r_105__73_, s_r_105__72_, s_r_105__71_, s_r_105__70_, s_r_105__69_, s_r_105__68_, s_r_105__67_, s_r_105__66_, s_r_105__65_, s_r_105__64_, s_r_105__63_, s_r_105__62_, s_r_105__61_, s_r_105__60_, s_r_105__59_, s_r_105__58_, s_r_105__57_, s_r_105__56_, s_r_105__55_, s_r_105__54_, s_r_105__53_, s_r_105__52_, s_r_105__51_, s_r_105__50_, s_r_105__49_, s_r_105__48_, s_r_105__47_, s_r_105__46_, s_r_105__45_, s_r_105__44_, s_r_105__43_, s_r_105__42_, s_r_105__41_, s_r_105__40_, s_r_105__39_, s_r_105__38_, s_r_105__37_, s_r_105__36_, s_r_105__35_, s_r_105__34_, s_r_105__33_, s_r_105__32_, s_r_105__31_, s_r_105__30_, s_r_105__29_, s_r_105__28_, s_r_105__27_, s_r_105__26_, s_r_105__25_, s_r_105__24_, s_r_105__23_, s_r_105__22_, s_r_105__21_, s_r_105__20_, s_r_105__19_, s_r_105__18_, s_r_105__17_, s_r_105__16_, s_r_105__15_, s_r_105__14_, s_r_105__13_, s_r_105__12_, s_r_105__11_, s_r_105__10_, s_r_105__9_, s_r_105__8_, s_r_105__7_, s_r_105__6_, s_r_105__5_, s_r_105__4_, s_r_105__3_, s_r_105__2_, s_r_105__1_, s_r_105__0_ }),
    .c_i(c_r[105]),
    .prod_accum_i({ prod_accum_105__106_, prod_accum_105__105_, prod_accum_105__104_, prod_accum_105__103_, prod_accum_105__102_, prod_accum_105__101_, prod_accum_105__100_, prod_accum_105__99_, prod_accum_105__98_, prod_accum_105__97_, prod_accum_105__96_, prod_accum_105__95_, prod_accum_105__94_, prod_accum_105__93_, prod_accum_105__92_, prod_accum_105__91_, prod_accum_105__90_, prod_accum_105__89_, prod_accum_105__88_, prod_accum_105__87_, prod_accum_105__86_, prod_accum_105__85_, prod_accum_105__84_, prod_accum_105__83_, prod_accum_105__82_, prod_accum_105__81_, prod_accum_105__80_, prod_accum_105__79_, prod_accum_105__78_, prod_accum_105__77_, prod_accum_105__76_, prod_accum_105__75_, prod_accum_105__74_, prod_accum_105__73_, prod_accum_105__72_, prod_accum_105__71_, prod_accum_105__70_, prod_accum_105__69_, prod_accum_105__68_, prod_accum_105__67_, prod_accum_105__66_, prod_accum_105__65_, prod_accum_105__64_, prod_accum_105__63_, prod_accum_105__62_, prod_accum_105__61_, prod_accum_105__60_, prod_accum_105__59_, prod_accum_105__58_, prod_accum_105__57_, prod_accum_105__56_, prod_accum_105__55_, prod_accum_105__54_, prod_accum_105__53_, prod_accum_105__52_, prod_accum_105__51_, prod_accum_105__50_, prod_accum_105__49_, prod_accum_105__48_, prod_accum_105__47_, prod_accum_105__46_, prod_accum_105__45_, prod_accum_105__44_, prod_accum_105__43_, prod_accum_105__42_, prod_accum_105__41_, prod_accum_105__40_, prod_accum_105__39_, prod_accum_105__38_, prod_accum_105__37_, prod_accum_105__36_, prod_accum_105__35_, prod_accum_105__34_, prod_accum_105__33_, prod_accum_105__32_, prod_accum_105__31_, prod_accum_105__30_, prod_accum_105__29_, prod_accum_105__28_, prod_accum_105__27_, prod_accum_105__26_, prod_accum_105__25_, prod_accum_105__24_, prod_accum_105__23_, prod_accum_105__22_, prod_accum_105__21_, prod_accum_105__20_, prod_accum_105__19_, prod_accum_105__18_, prod_accum_105__17_, prod_accum_105__16_, prod_accum_105__15_, prod_accum_105__14_, prod_accum_105__13_, prod_accum_105__12_, prod_accum_105__11_, prod_accum_105__10_, prod_accum_105__9_, prod_accum_105__8_, prod_accum_105__7_, prod_accum_105__6_, prod_accum_105__5_, prod_accum_105__4_, prod_accum_105__3_, prod_accum_105__2_, prod_accum_105__1_, prod_accum_105__0_ }),
    .a_o(a_r[13695:13568]),
    .b_o(b_r[13695:13568]),
    .s_o({ s_r_106__127_, s_r_106__126_, s_r_106__125_, s_r_106__124_, s_r_106__123_, s_r_106__122_, s_r_106__121_, s_r_106__120_, s_r_106__119_, s_r_106__118_, s_r_106__117_, s_r_106__116_, s_r_106__115_, s_r_106__114_, s_r_106__113_, s_r_106__112_, s_r_106__111_, s_r_106__110_, s_r_106__109_, s_r_106__108_, s_r_106__107_, s_r_106__106_, s_r_106__105_, s_r_106__104_, s_r_106__103_, s_r_106__102_, s_r_106__101_, s_r_106__100_, s_r_106__99_, s_r_106__98_, s_r_106__97_, s_r_106__96_, s_r_106__95_, s_r_106__94_, s_r_106__93_, s_r_106__92_, s_r_106__91_, s_r_106__90_, s_r_106__89_, s_r_106__88_, s_r_106__87_, s_r_106__86_, s_r_106__85_, s_r_106__84_, s_r_106__83_, s_r_106__82_, s_r_106__81_, s_r_106__80_, s_r_106__79_, s_r_106__78_, s_r_106__77_, s_r_106__76_, s_r_106__75_, s_r_106__74_, s_r_106__73_, s_r_106__72_, s_r_106__71_, s_r_106__70_, s_r_106__69_, s_r_106__68_, s_r_106__67_, s_r_106__66_, s_r_106__65_, s_r_106__64_, s_r_106__63_, s_r_106__62_, s_r_106__61_, s_r_106__60_, s_r_106__59_, s_r_106__58_, s_r_106__57_, s_r_106__56_, s_r_106__55_, s_r_106__54_, s_r_106__53_, s_r_106__52_, s_r_106__51_, s_r_106__50_, s_r_106__49_, s_r_106__48_, s_r_106__47_, s_r_106__46_, s_r_106__45_, s_r_106__44_, s_r_106__43_, s_r_106__42_, s_r_106__41_, s_r_106__40_, s_r_106__39_, s_r_106__38_, s_r_106__37_, s_r_106__36_, s_r_106__35_, s_r_106__34_, s_r_106__33_, s_r_106__32_, s_r_106__31_, s_r_106__30_, s_r_106__29_, s_r_106__28_, s_r_106__27_, s_r_106__26_, s_r_106__25_, s_r_106__24_, s_r_106__23_, s_r_106__22_, s_r_106__21_, s_r_106__20_, s_r_106__19_, s_r_106__18_, s_r_106__17_, s_r_106__16_, s_r_106__15_, s_r_106__14_, s_r_106__13_, s_r_106__12_, s_r_106__11_, s_r_106__10_, s_r_106__9_, s_r_106__8_, s_r_106__7_, s_r_106__6_, s_r_106__5_, s_r_106__4_, s_r_106__3_, s_r_106__2_, s_r_106__1_, s_r_106__0_ }),
    .c_o(c_r[106]),
    .prod_accum_o({ prod_accum_106__107_, prod_accum_106__106_, prod_accum_106__105_, prod_accum_106__104_, prod_accum_106__103_, prod_accum_106__102_, prod_accum_106__101_, prod_accum_106__100_, prod_accum_106__99_, prod_accum_106__98_, prod_accum_106__97_, prod_accum_106__96_, prod_accum_106__95_, prod_accum_106__94_, prod_accum_106__93_, prod_accum_106__92_, prod_accum_106__91_, prod_accum_106__90_, prod_accum_106__89_, prod_accum_106__88_, prod_accum_106__87_, prod_accum_106__86_, prod_accum_106__85_, prod_accum_106__84_, prod_accum_106__83_, prod_accum_106__82_, prod_accum_106__81_, prod_accum_106__80_, prod_accum_106__79_, prod_accum_106__78_, prod_accum_106__77_, prod_accum_106__76_, prod_accum_106__75_, prod_accum_106__74_, prod_accum_106__73_, prod_accum_106__72_, prod_accum_106__71_, prod_accum_106__70_, prod_accum_106__69_, prod_accum_106__68_, prod_accum_106__67_, prod_accum_106__66_, prod_accum_106__65_, prod_accum_106__64_, prod_accum_106__63_, prod_accum_106__62_, prod_accum_106__61_, prod_accum_106__60_, prod_accum_106__59_, prod_accum_106__58_, prod_accum_106__57_, prod_accum_106__56_, prod_accum_106__55_, prod_accum_106__54_, prod_accum_106__53_, prod_accum_106__52_, prod_accum_106__51_, prod_accum_106__50_, prod_accum_106__49_, prod_accum_106__48_, prod_accum_106__47_, prod_accum_106__46_, prod_accum_106__45_, prod_accum_106__44_, prod_accum_106__43_, prod_accum_106__42_, prod_accum_106__41_, prod_accum_106__40_, prod_accum_106__39_, prod_accum_106__38_, prod_accum_106__37_, prod_accum_106__36_, prod_accum_106__35_, prod_accum_106__34_, prod_accum_106__33_, prod_accum_106__32_, prod_accum_106__31_, prod_accum_106__30_, prod_accum_106__29_, prod_accum_106__28_, prod_accum_106__27_, prod_accum_106__26_, prod_accum_106__25_, prod_accum_106__24_, prod_accum_106__23_, prod_accum_106__22_, prod_accum_106__21_, prod_accum_106__20_, prod_accum_106__19_, prod_accum_106__18_, prod_accum_106__17_, prod_accum_106__16_, prod_accum_106__15_, prod_accum_106__14_, prod_accum_106__13_, prod_accum_106__12_, prod_accum_106__11_, prod_accum_106__10_, prod_accum_106__9_, prod_accum_106__8_, prod_accum_106__7_, prod_accum_106__6_, prod_accum_106__5_, prod_accum_106__4_, prod_accum_106__3_, prod_accum_106__2_, prod_accum_106__1_, prod_accum_106__0_ })
  );


  bsg_mul_array_row_128_107_x
  genblk1_107__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[13695:13568]),
    .b_i(b_r[13695:13568]),
    .s_i({ s_r_106__127_, s_r_106__126_, s_r_106__125_, s_r_106__124_, s_r_106__123_, s_r_106__122_, s_r_106__121_, s_r_106__120_, s_r_106__119_, s_r_106__118_, s_r_106__117_, s_r_106__116_, s_r_106__115_, s_r_106__114_, s_r_106__113_, s_r_106__112_, s_r_106__111_, s_r_106__110_, s_r_106__109_, s_r_106__108_, s_r_106__107_, s_r_106__106_, s_r_106__105_, s_r_106__104_, s_r_106__103_, s_r_106__102_, s_r_106__101_, s_r_106__100_, s_r_106__99_, s_r_106__98_, s_r_106__97_, s_r_106__96_, s_r_106__95_, s_r_106__94_, s_r_106__93_, s_r_106__92_, s_r_106__91_, s_r_106__90_, s_r_106__89_, s_r_106__88_, s_r_106__87_, s_r_106__86_, s_r_106__85_, s_r_106__84_, s_r_106__83_, s_r_106__82_, s_r_106__81_, s_r_106__80_, s_r_106__79_, s_r_106__78_, s_r_106__77_, s_r_106__76_, s_r_106__75_, s_r_106__74_, s_r_106__73_, s_r_106__72_, s_r_106__71_, s_r_106__70_, s_r_106__69_, s_r_106__68_, s_r_106__67_, s_r_106__66_, s_r_106__65_, s_r_106__64_, s_r_106__63_, s_r_106__62_, s_r_106__61_, s_r_106__60_, s_r_106__59_, s_r_106__58_, s_r_106__57_, s_r_106__56_, s_r_106__55_, s_r_106__54_, s_r_106__53_, s_r_106__52_, s_r_106__51_, s_r_106__50_, s_r_106__49_, s_r_106__48_, s_r_106__47_, s_r_106__46_, s_r_106__45_, s_r_106__44_, s_r_106__43_, s_r_106__42_, s_r_106__41_, s_r_106__40_, s_r_106__39_, s_r_106__38_, s_r_106__37_, s_r_106__36_, s_r_106__35_, s_r_106__34_, s_r_106__33_, s_r_106__32_, s_r_106__31_, s_r_106__30_, s_r_106__29_, s_r_106__28_, s_r_106__27_, s_r_106__26_, s_r_106__25_, s_r_106__24_, s_r_106__23_, s_r_106__22_, s_r_106__21_, s_r_106__20_, s_r_106__19_, s_r_106__18_, s_r_106__17_, s_r_106__16_, s_r_106__15_, s_r_106__14_, s_r_106__13_, s_r_106__12_, s_r_106__11_, s_r_106__10_, s_r_106__9_, s_r_106__8_, s_r_106__7_, s_r_106__6_, s_r_106__5_, s_r_106__4_, s_r_106__3_, s_r_106__2_, s_r_106__1_, s_r_106__0_ }),
    .c_i(c_r[106]),
    .prod_accum_i({ prod_accum_106__107_, prod_accum_106__106_, prod_accum_106__105_, prod_accum_106__104_, prod_accum_106__103_, prod_accum_106__102_, prod_accum_106__101_, prod_accum_106__100_, prod_accum_106__99_, prod_accum_106__98_, prod_accum_106__97_, prod_accum_106__96_, prod_accum_106__95_, prod_accum_106__94_, prod_accum_106__93_, prod_accum_106__92_, prod_accum_106__91_, prod_accum_106__90_, prod_accum_106__89_, prod_accum_106__88_, prod_accum_106__87_, prod_accum_106__86_, prod_accum_106__85_, prod_accum_106__84_, prod_accum_106__83_, prod_accum_106__82_, prod_accum_106__81_, prod_accum_106__80_, prod_accum_106__79_, prod_accum_106__78_, prod_accum_106__77_, prod_accum_106__76_, prod_accum_106__75_, prod_accum_106__74_, prod_accum_106__73_, prod_accum_106__72_, prod_accum_106__71_, prod_accum_106__70_, prod_accum_106__69_, prod_accum_106__68_, prod_accum_106__67_, prod_accum_106__66_, prod_accum_106__65_, prod_accum_106__64_, prod_accum_106__63_, prod_accum_106__62_, prod_accum_106__61_, prod_accum_106__60_, prod_accum_106__59_, prod_accum_106__58_, prod_accum_106__57_, prod_accum_106__56_, prod_accum_106__55_, prod_accum_106__54_, prod_accum_106__53_, prod_accum_106__52_, prod_accum_106__51_, prod_accum_106__50_, prod_accum_106__49_, prod_accum_106__48_, prod_accum_106__47_, prod_accum_106__46_, prod_accum_106__45_, prod_accum_106__44_, prod_accum_106__43_, prod_accum_106__42_, prod_accum_106__41_, prod_accum_106__40_, prod_accum_106__39_, prod_accum_106__38_, prod_accum_106__37_, prod_accum_106__36_, prod_accum_106__35_, prod_accum_106__34_, prod_accum_106__33_, prod_accum_106__32_, prod_accum_106__31_, prod_accum_106__30_, prod_accum_106__29_, prod_accum_106__28_, prod_accum_106__27_, prod_accum_106__26_, prod_accum_106__25_, prod_accum_106__24_, prod_accum_106__23_, prod_accum_106__22_, prod_accum_106__21_, prod_accum_106__20_, prod_accum_106__19_, prod_accum_106__18_, prod_accum_106__17_, prod_accum_106__16_, prod_accum_106__15_, prod_accum_106__14_, prod_accum_106__13_, prod_accum_106__12_, prod_accum_106__11_, prod_accum_106__10_, prod_accum_106__9_, prod_accum_106__8_, prod_accum_106__7_, prod_accum_106__6_, prod_accum_106__5_, prod_accum_106__4_, prod_accum_106__3_, prod_accum_106__2_, prod_accum_106__1_, prod_accum_106__0_ }),
    .a_o(a_r[13823:13696]),
    .b_o(b_r[13823:13696]),
    .s_o({ s_r_107__127_, s_r_107__126_, s_r_107__125_, s_r_107__124_, s_r_107__123_, s_r_107__122_, s_r_107__121_, s_r_107__120_, s_r_107__119_, s_r_107__118_, s_r_107__117_, s_r_107__116_, s_r_107__115_, s_r_107__114_, s_r_107__113_, s_r_107__112_, s_r_107__111_, s_r_107__110_, s_r_107__109_, s_r_107__108_, s_r_107__107_, s_r_107__106_, s_r_107__105_, s_r_107__104_, s_r_107__103_, s_r_107__102_, s_r_107__101_, s_r_107__100_, s_r_107__99_, s_r_107__98_, s_r_107__97_, s_r_107__96_, s_r_107__95_, s_r_107__94_, s_r_107__93_, s_r_107__92_, s_r_107__91_, s_r_107__90_, s_r_107__89_, s_r_107__88_, s_r_107__87_, s_r_107__86_, s_r_107__85_, s_r_107__84_, s_r_107__83_, s_r_107__82_, s_r_107__81_, s_r_107__80_, s_r_107__79_, s_r_107__78_, s_r_107__77_, s_r_107__76_, s_r_107__75_, s_r_107__74_, s_r_107__73_, s_r_107__72_, s_r_107__71_, s_r_107__70_, s_r_107__69_, s_r_107__68_, s_r_107__67_, s_r_107__66_, s_r_107__65_, s_r_107__64_, s_r_107__63_, s_r_107__62_, s_r_107__61_, s_r_107__60_, s_r_107__59_, s_r_107__58_, s_r_107__57_, s_r_107__56_, s_r_107__55_, s_r_107__54_, s_r_107__53_, s_r_107__52_, s_r_107__51_, s_r_107__50_, s_r_107__49_, s_r_107__48_, s_r_107__47_, s_r_107__46_, s_r_107__45_, s_r_107__44_, s_r_107__43_, s_r_107__42_, s_r_107__41_, s_r_107__40_, s_r_107__39_, s_r_107__38_, s_r_107__37_, s_r_107__36_, s_r_107__35_, s_r_107__34_, s_r_107__33_, s_r_107__32_, s_r_107__31_, s_r_107__30_, s_r_107__29_, s_r_107__28_, s_r_107__27_, s_r_107__26_, s_r_107__25_, s_r_107__24_, s_r_107__23_, s_r_107__22_, s_r_107__21_, s_r_107__20_, s_r_107__19_, s_r_107__18_, s_r_107__17_, s_r_107__16_, s_r_107__15_, s_r_107__14_, s_r_107__13_, s_r_107__12_, s_r_107__11_, s_r_107__10_, s_r_107__9_, s_r_107__8_, s_r_107__7_, s_r_107__6_, s_r_107__5_, s_r_107__4_, s_r_107__3_, s_r_107__2_, s_r_107__1_, s_r_107__0_ }),
    .c_o(c_r[107]),
    .prod_accum_o({ prod_accum_107__108_, prod_accum_107__107_, prod_accum_107__106_, prod_accum_107__105_, prod_accum_107__104_, prod_accum_107__103_, prod_accum_107__102_, prod_accum_107__101_, prod_accum_107__100_, prod_accum_107__99_, prod_accum_107__98_, prod_accum_107__97_, prod_accum_107__96_, prod_accum_107__95_, prod_accum_107__94_, prod_accum_107__93_, prod_accum_107__92_, prod_accum_107__91_, prod_accum_107__90_, prod_accum_107__89_, prod_accum_107__88_, prod_accum_107__87_, prod_accum_107__86_, prod_accum_107__85_, prod_accum_107__84_, prod_accum_107__83_, prod_accum_107__82_, prod_accum_107__81_, prod_accum_107__80_, prod_accum_107__79_, prod_accum_107__78_, prod_accum_107__77_, prod_accum_107__76_, prod_accum_107__75_, prod_accum_107__74_, prod_accum_107__73_, prod_accum_107__72_, prod_accum_107__71_, prod_accum_107__70_, prod_accum_107__69_, prod_accum_107__68_, prod_accum_107__67_, prod_accum_107__66_, prod_accum_107__65_, prod_accum_107__64_, prod_accum_107__63_, prod_accum_107__62_, prod_accum_107__61_, prod_accum_107__60_, prod_accum_107__59_, prod_accum_107__58_, prod_accum_107__57_, prod_accum_107__56_, prod_accum_107__55_, prod_accum_107__54_, prod_accum_107__53_, prod_accum_107__52_, prod_accum_107__51_, prod_accum_107__50_, prod_accum_107__49_, prod_accum_107__48_, prod_accum_107__47_, prod_accum_107__46_, prod_accum_107__45_, prod_accum_107__44_, prod_accum_107__43_, prod_accum_107__42_, prod_accum_107__41_, prod_accum_107__40_, prod_accum_107__39_, prod_accum_107__38_, prod_accum_107__37_, prod_accum_107__36_, prod_accum_107__35_, prod_accum_107__34_, prod_accum_107__33_, prod_accum_107__32_, prod_accum_107__31_, prod_accum_107__30_, prod_accum_107__29_, prod_accum_107__28_, prod_accum_107__27_, prod_accum_107__26_, prod_accum_107__25_, prod_accum_107__24_, prod_accum_107__23_, prod_accum_107__22_, prod_accum_107__21_, prod_accum_107__20_, prod_accum_107__19_, prod_accum_107__18_, prod_accum_107__17_, prod_accum_107__16_, prod_accum_107__15_, prod_accum_107__14_, prod_accum_107__13_, prod_accum_107__12_, prod_accum_107__11_, prod_accum_107__10_, prod_accum_107__9_, prod_accum_107__8_, prod_accum_107__7_, prod_accum_107__6_, prod_accum_107__5_, prod_accum_107__4_, prod_accum_107__3_, prod_accum_107__2_, prod_accum_107__1_, prod_accum_107__0_ })
  );


  bsg_mul_array_row_128_108_x
  genblk1_108__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[13823:13696]),
    .b_i(b_r[13823:13696]),
    .s_i({ s_r_107__127_, s_r_107__126_, s_r_107__125_, s_r_107__124_, s_r_107__123_, s_r_107__122_, s_r_107__121_, s_r_107__120_, s_r_107__119_, s_r_107__118_, s_r_107__117_, s_r_107__116_, s_r_107__115_, s_r_107__114_, s_r_107__113_, s_r_107__112_, s_r_107__111_, s_r_107__110_, s_r_107__109_, s_r_107__108_, s_r_107__107_, s_r_107__106_, s_r_107__105_, s_r_107__104_, s_r_107__103_, s_r_107__102_, s_r_107__101_, s_r_107__100_, s_r_107__99_, s_r_107__98_, s_r_107__97_, s_r_107__96_, s_r_107__95_, s_r_107__94_, s_r_107__93_, s_r_107__92_, s_r_107__91_, s_r_107__90_, s_r_107__89_, s_r_107__88_, s_r_107__87_, s_r_107__86_, s_r_107__85_, s_r_107__84_, s_r_107__83_, s_r_107__82_, s_r_107__81_, s_r_107__80_, s_r_107__79_, s_r_107__78_, s_r_107__77_, s_r_107__76_, s_r_107__75_, s_r_107__74_, s_r_107__73_, s_r_107__72_, s_r_107__71_, s_r_107__70_, s_r_107__69_, s_r_107__68_, s_r_107__67_, s_r_107__66_, s_r_107__65_, s_r_107__64_, s_r_107__63_, s_r_107__62_, s_r_107__61_, s_r_107__60_, s_r_107__59_, s_r_107__58_, s_r_107__57_, s_r_107__56_, s_r_107__55_, s_r_107__54_, s_r_107__53_, s_r_107__52_, s_r_107__51_, s_r_107__50_, s_r_107__49_, s_r_107__48_, s_r_107__47_, s_r_107__46_, s_r_107__45_, s_r_107__44_, s_r_107__43_, s_r_107__42_, s_r_107__41_, s_r_107__40_, s_r_107__39_, s_r_107__38_, s_r_107__37_, s_r_107__36_, s_r_107__35_, s_r_107__34_, s_r_107__33_, s_r_107__32_, s_r_107__31_, s_r_107__30_, s_r_107__29_, s_r_107__28_, s_r_107__27_, s_r_107__26_, s_r_107__25_, s_r_107__24_, s_r_107__23_, s_r_107__22_, s_r_107__21_, s_r_107__20_, s_r_107__19_, s_r_107__18_, s_r_107__17_, s_r_107__16_, s_r_107__15_, s_r_107__14_, s_r_107__13_, s_r_107__12_, s_r_107__11_, s_r_107__10_, s_r_107__9_, s_r_107__8_, s_r_107__7_, s_r_107__6_, s_r_107__5_, s_r_107__4_, s_r_107__3_, s_r_107__2_, s_r_107__1_, s_r_107__0_ }),
    .c_i(c_r[107]),
    .prod_accum_i({ prod_accum_107__108_, prod_accum_107__107_, prod_accum_107__106_, prod_accum_107__105_, prod_accum_107__104_, prod_accum_107__103_, prod_accum_107__102_, prod_accum_107__101_, prod_accum_107__100_, prod_accum_107__99_, prod_accum_107__98_, prod_accum_107__97_, prod_accum_107__96_, prod_accum_107__95_, prod_accum_107__94_, prod_accum_107__93_, prod_accum_107__92_, prod_accum_107__91_, prod_accum_107__90_, prod_accum_107__89_, prod_accum_107__88_, prod_accum_107__87_, prod_accum_107__86_, prod_accum_107__85_, prod_accum_107__84_, prod_accum_107__83_, prod_accum_107__82_, prod_accum_107__81_, prod_accum_107__80_, prod_accum_107__79_, prod_accum_107__78_, prod_accum_107__77_, prod_accum_107__76_, prod_accum_107__75_, prod_accum_107__74_, prod_accum_107__73_, prod_accum_107__72_, prod_accum_107__71_, prod_accum_107__70_, prod_accum_107__69_, prod_accum_107__68_, prod_accum_107__67_, prod_accum_107__66_, prod_accum_107__65_, prod_accum_107__64_, prod_accum_107__63_, prod_accum_107__62_, prod_accum_107__61_, prod_accum_107__60_, prod_accum_107__59_, prod_accum_107__58_, prod_accum_107__57_, prod_accum_107__56_, prod_accum_107__55_, prod_accum_107__54_, prod_accum_107__53_, prod_accum_107__52_, prod_accum_107__51_, prod_accum_107__50_, prod_accum_107__49_, prod_accum_107__48_, prod_accum_107__47_, prod_accum_107__46_, prod_accum_107__45_, prod_accum_107__44_, prod_accum_107__43_, prod_accum_107__42_, prod_accum_107__41_, prod_accum_107__40_, prod_accum_107__39_, prod_accum_107__38_, prod_accum_107__37_, prod_accum_107__36_, prod_accum_107__35_, prod_accum_107__34_, prod_accum_107__33_, prod_accum_107__32_, prod_accum_107__31_, prod_accum_107__30_, prod_accum_107__29_, prod_accum_107__28_, prod_accum_107__27_, prod_accum_107__26_, prod_accum_107__25_, prod_accum_107__24_, prod_accum_107__23_, prod_accum_107__22_, prod_accum_107__21_, prod_accum_107__20_, prod_accum_107__19_, prod_accum_107__18_, prod_accum_107__17_, prod_accum_107__16_, prod_accum_107__15_, prod_accum_107__14_, prod_accum_107__13_, prod_accum_107__12_, prod_accum_107__11_, prod_accum_107__10_, prod_accum_107__9_, prod_accum_107__8_, prod_accum_107__7_, prod_accum_107__6_, prod_accum_107__5_, prod_accum_107__4_, prod_accum_107__3_, prod_accum_107__2_, prod_accum_107__1_, prod_accum_107__0_ }),
    .a_o(a_r[13951:13824]),
    .b_o(b_r[13951:13824]),
    .s_o({ s_r_108__127_, s_r_108__126_, s_r_108__125_, s_r_108__124_, s_r_108__123_, s_r_108__122_, s_r_108__121_, s_r_108__120_, s_r_108__119_, s_r_108__118_, s_r_108__117_, s_r_108__116_, s_r_108__115_, s_r_108__114_, s_r_108__113_, s_r_108__112_, s_r_108__111_, s_r_108__110_, s_r_108__109_, s_r_108__108_, s_r_108__107_, s_r_108__106_, s_r_108__105_, s_r_108__104_, s_r_108__103_, s_r_108__102_, s_r_108__101_, s_r_108__100_, s_r_108__99_, s_r_108__98_, s_r_108__97_, s_r_108__96_, s_r_108__95_, s_r_108__94_, s_r_108__93_, s_r_108__92_, s_r_108__91_, s_r_108__90_, s_r_108__89_, s_r_108__88_, s_r_108__87_, s_r_108__86_, s_r_108__85_, s_r_108__84_, s_r_108__83_, s_r_108__82_, s_r_108__81_, s_r_108__80_, s_r_108__79_, s_r_108__78_, s_r_108__77_, s_r_108__76_, s_r_108__75_, s_r_108__74_, s_r_108__73_, s_r_108__72_, s_r_108__71_, s_r_108__70_, s_r_108__69_, s_r_108__68_, s_r_108__67_, s_r_108__66_, s_r_108__65_, s_r_108__64_, s_r_108__63_, s_r_108__62_, s_r_108__61_, s_r_108__60_, s_r_108__59_, s_r_108__58_, s_r_108__57_, s_r_108__56_, s_r_108__55_, s_r_108__54_, s_r_108__53_, s_r_108__52_, s_r_108__51_, s_r_108__50_, s_r_108__49_, s_r_108__48_, s_r_108__47_, s_r_108__46_, s_r_108__45_, s_r_108__44_, s_r_108__43_, s_r_108__42_, s_r_108__41_, s_r_108__40_, s_r_108__39_, s_r_108__38_, s_r_108__37_, s_r_108__36_, s_r_108__35_, s_r_108__34_, s_r_108__33_, s_r_108__32_, s_r_108__31_, s_r_108__30_, s_r_108__29_, s_r_108__28_, s_r_108__27_, s_r_108__26_, s_r_108__25_, s_r_108__24_, s_r_108__23_, s_r_108__22_, s_r_108__21_, s_r_108__20_, s_r_108__19_, s_r_108__18_, s_r_108__17_, s_r_108__16_, s_r_108__15_, s_r_108__14_, s_r_108__13_, s_r_108__12_, s_r_108__11_, s_r_108__10_, s_r_108__9_, s_r_108__8_, s_r_108__7_, s_r_108__6_, s_r_108__5_, s_r_108__4_, s_r_108__3_, s_r_108__2_, s_r_108__1_, s_r_108__0_ }),
    .c_o(c_r[108]),
    .prod_accum_o({ prod_accum_108__109_, prod_accum_108__108_, prod_accum_108__107_, prod_accum_108__106_, prod_accum_108__105_, prod_accum_108__104_, prod_accum_108__103_, prod_accum_108__102_, prod_accum_108__101_, prod_accum_108__100_, prod_accum_108__99_, prod_accum_108__98_, prod_accum_108__97_, prod_accum_108__96_, prod_accum_108__95_, prod_accum_108__94_, prod_accum_108__93_, prod_accum_108__92_, prod_accum_108__91_, prod_accum_108__90_, prod_accum_108__89_, prod_accum_108__88_, prod_accum_108__87_, prod_accum_108__86_, prod_accum_108__85_, prod_accum_108__84_, prod_accum_108__83_, prod_accum_108__82_, prod_accum_108__81_, prod_accum_108__80_, prod_accum_108__79_, prod_accum_108__78_, prod_accum_108__77_, prod_accum_108__76_, prod_accum_108__75_, prod_accum_108__74_, prod_accum_108__73_, prod_accum_108__72_, prod_accum_108__71_, prod_accum_108__70_, prod_accum_108__69_, prod_accum_108__68_, prod_accum_108__67_, prod_accum_108__66_, prod_accum_108__65_, prod_accum_108__64_, prod_accum_108__63_, prod_accum_108__62_, prod_accum_108__61_, prod_accum_108__60_, prod_accum_108__59_, prod_accum_108__58_, prod_accum_108__57_, prod_accum_108__56_, prod_accum_108__55_, prod_accum_108__54_, prod_accum_108__53_, prod_accum_108__52_, prod_accum_108__51_, prod_accum_108__50_, prod_accum_108__49_, prod_accum_108__48_, prod_accum_108__47_, prod_accum_108__46_, prod_accum_108__45_, prod_accum_108__44_, prod_accum_108__43_, prod_accum_108__42_, prod_accum_108__41_, prod_accum_108__40_, prod_accum_108__39_, prod_accum_108__38_, prod_accum_108__37_, prod_accum_108__36_, prod_accum_108__35_, prod_accum_108__34_, prod_accum_108__33_, prod_accum_108__32_, prod_accum_108__31_, prod_accum_108__30_, prod_accum_108__29_, prod_accum_108__28_, prod_accum_108__27_, prod_accum_108__26_, prod_accum_108__25_, prod_accum_108__24_, prod_accum_108__23_, prod_accum_108__22_, prod_accum_108__21_, prod_accum_108__20_, prod_accum_108__19_, prod_accum_108__18_, prod_accum_108__17_, prod_accum_108__16_, prod_accum_108__15_, prod_accum_108__14_, prod_accum_108__13_, prod_accum_108__12_, prod_accum_108__11_, prod_accum_108__10_, prod_accum_108__9_, prod_accum_108__8_, prod_accum_108__7_, prod_accum_108__6_, prod_accum_108__5_, prod_accum_108__4_, prod_accum_108__3_, prod_accum_108__2_, prod_accum_108__1_, prod_accum_108__0_ })
  );


  bsg_mul_array_row_128_109_x
  genblk1_109__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[13951:13824]),
    .b_i(b_r[13951:13824]),
    .s_i({ s_r_108__127_, s_r_108__126_, s_r_108__125_, s_r_108__124_, s_r_108__123_, s_r_108__122_, s_r_108__121_, s_r_108__120_, s_r_108__119_, s_r_108__118_, s_r_108__117_, s_r_108__116_, s_r_108__115_, s_r_108__114_, s_r_108__113_, s_r_108__112_, s_r_108__111_, s_r_108__110_, s_r_108__109_, s_r_108__108_, s_r_108__107_, s_r_108__106_, s_r_108__105_, s_r_108__104_, s_r_108__103_, s_r_108__102_, s_r_108__101_, s_r_108__100_, s_r_108__99_, s_r_108__98_, s_r_108__97_, s_r_108__96_, s_r_108__95_, s_r_108__94_, s_r_108__93_, s_r_108__92_, s_r_108__91_, s_r_108__90_, s_r_108__89_, s_r_108__88_, s_r_108__87_, s_r_108__86_, s_r_108__85_, s_r_108__84_, s_r_108__83_, s_r_108__82_, s_r_108__81_, s_r_108__80_, s_r_108__79_, s_r_108__78_, s_r_108__77_, s_r_108__76_, s_r_108__75_, s_r_108__74_, s_r_108__73_, s_r_108__72_, s_r_108__71_, s_r_108__70_, s_r_108__69_, s_r_108__68_, s_r_108__67_, s_r_108__66_, s_r_108__65_, s_r_108__64_, s_r_108__63_, s_r_108__62_, s_r_108__61_, s_r_108__60_, s_r_108__59_, s_r_108__58_, s_r_108__57_, s_r_108__56_, s_r_108__55_, s_r_108__54_, s_r_108__53_, s_r_108__52_, s_r_108__51_, s_r_108__50_, s_r_108__49_, s_r_108__48_, s_r_108__47_, s_r_108__46_, s_r_108__45_, s_r_108__44_, s_r_108__43_, s_r_108__42_, s_r_108__41_, s_r_108__40_, s_r_108__39_, s_r_108__38_, s_r_108__37_, s_r_108__36_, s_r_108__35_, s_r_108__34_, s_r_108__33_, s_r_108__32_, s_r_108__31_, s_r_108__30_, s_r_108__29_, s_r_108__28_, s_r_108__27_, s_r_108__26_, s_r_108__25_, s_r_108__24_, s_r_108__23_, s_r_108__22_, s_r_108__21_, s_r_108__20_, s_r_108__19_, s_r_108__18_, s_r_108__17_, s_r_108__16_, s_r_108__15_, s_r_108__14_, s_r_108__13_, s_r_108__12_, s_r_108__11_, s_r_108__10_, s_r_108__9_, s_r_108__8_, s_r_108__7_, s_r_108__6_, s_r_108__5_, s_r_108__4_, s_r_108__3_, s_r_108__2_, s_r_108__1_, s_r_108__0_ }),
    .c_i(c_r[108]),
    .prod_accum_i({ prod_accum_108__109_, prod_accum_108__108_, prod_accum_108__107_, prod_accum_108__106_, prod_accum_108__105_, prod_accum_108__104_, prod_accum_108__103_, prod_accum_108__102_, prod_accum_108__101_, prod_accum_108__100_, prod_accum_108__99_, prod_accum_108__98_, prod_accum_108__97_, prod_accum_108__96_, prod_accum_108__95_, prod_accum_108__94_, prod_accum_108__93_, prod_accum_108__92_, prod_accum_108__91_, prod_accum_108__90_, prod_accum_108__89_, prod_accum_108__88_, prod_accum_108__87_, prod_accum_108__86_, prod_accum_108__85_, prod_accum_108__84_, prod_accum_108__83_, prod_accum_108__82_, prod_accum_108__81_, prod_accum_108__80_, prod_accum_108__79_, prod_accum_108__78_, prod_accum_108__77_, prod_accum_108__76_, prod_accum_108__75_, prod_accum_108__74_, prod_accum_108__73_, prod_accum_108__72_, prod_accum_108__71_, prod_accum_108__70_, prod_accum_108__69_, prod_accum_108__68_, prod_accum_108__67_, prod_accum_108__66_, prod_accum_108__65_, prod_accum_108__64_, prod_accum_108__63_, prod_accum_108__62_, prod_accum_108__61_, prod_accum_108__60_, prod_accum_108__59_, prod_accum_108__58_, prod_accum_108__57_, prod_accum_108__56_, prod_accum_108__55_, prod_accum_108__54_, prod_accum_108__53_, prod_accum_108__52_, prod_accum_108__51_, prod_accum_108__50_, prod_accum_108__49_, prod_accum_108__48_, prod_accum_108__47_, prod_accum_108__46_, prod_accum_108__45_, prod_accum_108__44_, prod_accum_108__43_, prod_accum_108__42_, prod_accum_108__41_, prod_accum_108__40_, prod_accum_108__39_, prod_accum_108__38_, prod_accum_108__37_, prod_accum_108__36_, prod_accum_108__35_, prod_accum_108__34_, prod_accum_108__33_, prod_accum_108__32_, prod_accum_108__31_, prod_accum_108__30_, prod_accum_108__29_, prod_accum_108__28_, prod_accum_108__27_, prod_accum_108__26_, prod_accum_108__25_, prod_accum_108__24_, prod_accum_108__23_, prod_accum_108__22_, prod_accum_108__21_, prod_accum_108__20_, prod_accum_108__19_, prod_accum_108__18_, prod_accum_108__17_, prod_accum_108__16_, prod_accum_108__15_, prod_accum_108__14_, prod_accum_108__13_, prod_accum_108__12_, prod_accum_108__11_, prod_accum_108__10_, prod_accum_108__9_, prod_accum_108__8_, prod_accum_108__7_, prod_accum_108__6_, prod_accum_108__5_, prod_accum_108__4_, prod_accum_108__3_, prod_accum_108__2_, prod_accum_108__1_, prod_accum_108__0_ }),
    .a_o(a_r[14079:13952]),
    .b_o(b_r[14079:13952]),
    .s_o({ s_r_109__127_, s_r_109__126_, s_r_109__125_, s_r_109__124_, s_r_109__123_, s_r_109__122_, s_r_109__121_, s_r_109__120_, s_r_109__119_, s_r_109__118_, s_r_109__117_, s_r_109__116_, s_r_109__115_, s_r_109__114_, s_r_109__113_, s_r_109__112_, s_r_109__111_, s_r_109__110_, s_r_109__109_, s_r_109__108_, s_r_109__107_, s_r_109__106_, s_r_109__105_, s_r_109__104_, s_r_109__103_, s_r_109__102_, s_r_109__101_, s_r_109__100_, s_r_109__99_, s_r_109__98_, s_r_109__97_, s_r_109__96_, s_r_109__95_, s_r_109__94_, s_r_109__93_, s_r_109__92_, s_r_109__91_, s_r_109__90_, s_r_109__89_, s_r_109__88_, s_r_109__87_, s_r_109__86_, s_r_109__85_, s_r_109__84_, s_r_109__83_, s_r_109__82_, s_r_109__81_, s_r_109__80_, s_r_109__79_, s_r_109__78_, s_r_109__77_, s_r_109__76_, s_r_109__75_, s_r_109__74_, s_r_109__73_, s_r_109__72_, s_r_109__71_, s_r_109__70_, s_r_109__69_, s_r_109__68_, s_r_109__67_, s_r_109__66_, s_r_109__65_, s_r_109__64_, s_r_109__63_, s_r_109__62_, s_r_109__61_, s_r_109__60_, s_r_109__59_, s_r_109__58_, s_r_109__57_, s_r_109__56_, s_r_109__55_, s_r_109__54_, s_r_109__53_, s_r_109__52_, s_r_109__51_, s_r_109__50_, s_r_109__49_, s_r_109__48_, s_r_109__47_, s_r_109__46_, s_r_109__45_, s_r_109__44_, s_r_109__43_, s_r_109__42_, s_r_109__41_, s_r_109__40_, s_r_109__39_, s_r_109__38_, s_r_109__37_, s_r_109__36_, s_r_109__35_, s_r_109__34_, s_r_109__33_, s_r_109__32_, s_r_109__31_, s_r_109__30_, s_r_109__29_, s_r_109__28_, s_r_109__27_, s_r_109__26_, s_r_109__25_, s_r_109__24_, s_r_109__23_, s_r_109__22_, s_r_109__21_, s_r_109__20_, s_r_109__19_, s_r_109__18_, s_r_109__17_, s_r_109__16_, s_r_109__15_, s_r_109__14_, s_r_109__13_, s_r_109__12_, s_r_109__11_, s_r_109__10_, s_r_109__9_, s_r_109__8_, s_r_109__7_, s_r_109__6_, s_r_109__5_, s_r_109__4_, s_r_109__3_, s_r_109__2_, s_r_109__1_, s_r_109__0_ }),
    .c_o(c_r[109]),
    .prod_accum_o({ prod_accum_109__110_, prod_accum_109__109_, prod_accum_109__108_, prod_accum_109__107_, prod_accum_109__106_, prod_accum_109__105_, prod_accum_109__104_, prod_accum_109__103_, prod_accum_109__102_, prod_accum_109__101_, prod_accum_109__100_, prod_accum_109__99_, prod_accum_109__98_, prod_accum_109__97_, prod_accum_109__96_, prod_accum_109__95_, prod_accum_109__94_, prod_accum_109__93_, prod_accum_109__92_, prod_accum_109__91_, prod_accum_109__90_, prod_accum_109__89_, prod_accum_109__88_, prod_accum_109__87_, prod_accum_109__86_, prod_accum_109__85_, prod_accum_109__84_, prod_accum_109__83_, prod_accum_109__82_, prod_accum_109__81_, prod_accum_109__80_, prod_accum_109__79_, prod_accum_109__78_, prod_accum_109__77_, prod_accum_109__76_, prod_accum_109__75_, prod_accum_109__74_, prod_accum_109__73_, prod_accum_109__72_, prod_accum_109__71_, prod_accum_109__70_, prod_accum_109__69_, prod_accum_109__68_, prod_accum_109__67_, prod_accum_109__66_, prod_accum_109__65_, prod_accum_109__64_, prod_accum_109__63_, prod_accum_109__62_, prod_accum_109__61_, prod_accum_109__60_, prod_accum_109__59_, prod_accum_109__58_, prod_accum_109__57_, prod_accum_109__56_, prod_accum_109__55_, prod_accum_109__54_, prod_accum_109__53_, prod_accum_109__52_, prod_accum_109__51_, prod_accum_109__50_, prod_accum_109__49_, prod_accum_109__48_, prod_accum_109__47_, prod_accum_109__46_, prod_accum_109__45_, prod_accum_109__44_, prod_accum_109__43_, prod_accum_109__42_, prod_accum_109__41_, prod_accum_109__40_, prod_accum_109__39_, prod_accum_109__38_, prod_accum_109__37_, prod_accum_109__36_, prod_accum_109__35_, prod_accum_109__34_, prod_accum_109__33_, prod_accum_109__32_, prod_accum_109__31_, prod_accum_109__30_, prod_accum_109__29_, prod_accum_109__28_, prod_accum_109__27_, prod_accum_109__26_, prod_accum_109__25_, prod_accum_109__24_, prod_accum_109__23_, prod_accum_109__22_, prod_accum_109__21_, prod_accum_109__20_, prod_accum_109__19_, prod_accum_109__18_, prod_accum_109__17_, prod_accum_109__16_, prod_accum_109__15_, prod_accum_109__14_, prod_accum_109__13_, prod_accum_109__12_, prod_accum_109__11_, prod_accum_109__10_, prod_accum_109__9_, prod_accum_109__8_, prod_accum_109__7_, prod_accum_109__6_, prod_accum_109__5_, prod_accum_109__4_, prod_accum_109__3_, prod_accum_109__2_, prod_accum_109__1_, prod_accum_109__0_ })
  );


  bsg_mul_array_row_128_110_x
  genblk1_110__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[14079:13952]),
    .b_i(b_r[14079:13952]),
    .s_i({ s_r_109__127_, s_r_109__126_, s_r_109__125_, s_r_109__124_, s_r_109__123_, s_r_109__122_, s_r_109__121_, s_r_109__120_, s_r_109__119_, s_r_109__118_, s_r_109__117_, s_r_109__116_, s_r_109__115_, s_r_109__114_, s_r_109__113_, s_r_109__112_, s_r_109__111_, s_r_109__110_, s_r_109__109_, s_r_109__108_, s_r_109__107_, s_r_109__106_, s_r_109__105_, s_r_109__104_, s_r_109__103_, s_r_109__102_, s_r_109__101_, s_r_109__100_, s_r_109__99_, s_r_109__98_, s_r_109__97_, s_r_109__96_, s_r_109__95_, s_r_109__94_, s_r_109__93_, s_r_109__92_, s_r_109__91_, s_r_109__90_, s_r_109__89_, s_r_109__88_, s_r_109__87_, s_r_109__86_, s_r_109__85_, s_r_109__84_, s_r_109__83_, s_r_109__82_, s_r_109__81_, s_r_109__80_, s_r_109__79_, s_r_109__78_, s_r_109__77_, s_r_109__76_, s_r_109__75_, s_r_109__74_, s_r_109__73_, s_r_109__72_, s_r_109__71_, s_r_109__70_, s_r_109__69_, s_r_109__68_, s_r_109__67_, s_r_109__66_, s_r_109__65_, s_r_109__64_, s_r_109__63_, s_r_109__62_, s_r_109__61_, s_r_109__60_, s_r_109__59_, s_r_109__58_, s_r_109__57_, s_r_109__56_, s_r_109__55_, s_r_109__54_, s_r_109__53_, s_r_109__52_, s_r_109__51_, s_r_109__50_, s_r_109__49_, s_r_109__48_, s_r_109__47_, s_r_109__46_, s_r_109__45_, s_r_109__44_, s_r_109__43_, s_r_109__42_, s_r_109__41_, s_r_109__40_, s_r_109__39_, s_r_109__38_, s_r_109__37_, s_r_109__36_, s_r_109__35_, s_r_109__34_, s_r_109__33_, s_r_109__32_, s_r_109__31_, s_r_109__30_, s_r_109__29_, s_r_109__28_, s_r_109__27_, s_r_109__26_, s_r_109__25_, s_r_109__24_, s_r_109__23_, s_r_109__22_, s_r_109__21_, s_r_109__20_, s_r_109__19_, s_r_109__18_, s_r_109__17_, s_r_109__16_, s_r_109__15_, s_r_109__14_, s_r_109__13_, s_r_109__12_, s_r_109__11_, s_r_109__10_, s_r_109__9_, s_r_109__8_, s_r_109__7_, s_r_109__6_, s_r_109__5_, s_r_109__4_, s_r_109__3_, s_r_109__2_, s_r_109__1_, s_r_109__0_ }),
    .c_i(c_r[109]),
    .prod_accum_i({ prod_accum_109__110_, prod_accum_109__109_, prod_accum_109__108_, prod_accum_109__107_, prod_accum_109__106_, prod_accum_109__105_, prod_accum_109__104_, prod_accum_109__103_, prod_accum_109__102_, prod_accum_109__101_, prod_accum_109__100_, prod_accum_109__99_, prod_accum_109__98_, prod_accum_109__97_, prod_accum_109__96_, prod_accum_109__95_, prod_accum_109__94_, prod_accum_109__93_, prod_accum_109__92_, prod_accum_109__91_, prod_accum_109__90_, prod_accum_109__89_, prod_accum_109__88_, prod_accum_109__87_, prod_accum_109__86_, prod_accum_109__85_, prod_accum_109__84_, prod_accum_109__83_, prod_accum_109__82_, prod_accum_109__81_, prod_accum_109__80_, prod_accum_109__79_, prod_accum_109__78_, prod_accum_109__77_, prod_accum_109__76_, prod_accum_109__75_, prod_accum_109__74_, prod_accum_109__73_, prod_accum_109__72_, prod_accum_109__71_, prod_accum_109__70_, prod_accum_109__69_, prod_accum_109__68_, prod_accum_109__67_, prod_accum_109__66_, prod_accum_109__65_, prod_accum_109__64_, prod_accum_109__63_, prod_accum_109__62_, prod_accum_109__61_, prod_accum_109__60_, prod_accum_109__59_, prod_accum_109__58_, prod_accum_109__57_, prod_accum_109__56_, prod_accum_109__55_, prod_accum_109__54_, prod_accum_109__53_, prod_accum_109__52_, prod_accum_109__51_, prod_accum_109__50_, prod_accum_109__49_, prod_accum_109__48_, prod_accum_109__47_, prod_accum_109__46_, prod_accum_109__45_, prod_accum_109__44_, prod_accum_109__43_, prod_accum_109__42_, prod_accum_109__41_, prod_accum_109__40_, prod_accum_109__39_, prod_accum_109__38_, prod_accum_109__37_, prod_accum_109__36_, prod_accum_109__35_, prod_accum_109__34_, prod_accum_109__33_, prod_accum_109__32_, prod_accum_109__31_, prod_accum_109__30_, prod_accum_109__29_, prod_accum_109__28_, prod_accum_109__27_, prod_accum_109__26_, prod_accum_109__25_, prod_accum_109__24_, prod_accum_109__23_, prod_accum_109__22_, prod_accum_109__21_, prod_accum_109__20_, prod_accum_109__19_, prod_accum_109__18_, prod_accum_109__17_, prod_accum_109__16_, prod_accum_109__15_, prod_accum_109__14_, prod_accum_109__13_, prod_accum_109__12_, prod_accum_109__11_, prod_accum_109__10_, prod_accum_109__9_, prod_accum_109__8_, prod_accum_109__7_, prod_accum_109__6_, prod_accum_109__5_, prod_accum_109__4_, prod_accum_109__3_, prod_accum_109__2_, prod_accum_109__1_, prod_accum_109__0_ }),
    .a_o(a_r[14207:14080]),
    .b_o(b_r[14207:14080]),
    .s_o({ s_r_110__127_, s_r_110__126_, s_r_110__125_, s_r_110__124_, s_r_110__123_, s_r_110__122_, s_r_110__121_, s_r_110__120_, s_r_110__119_, s_r_110__118_, s_r_110__117_, s_r_110__116_, s_r_110__115_, s_r_110__114_, s_r_110__113_, s_r_110__112_, s_r_110__111_, s_r_110__110_, s_r_110__109_, s_r_110__108_, s_r_110__107_, s_r_110__106_, s_r_110__105_, s_r_110__104_, s_r_110__103_, s_r_110__102_, s_r_110__101_, s_r_110__100_, s_r_110__99_, s_r_110__98_, s_r_110__97_, s_r_110__96_, s_r_110__95_, s_r_110__94_, s_r_110__93_, s_r_110__92_, s_r_110__91_, s_r_110__90_, s_r_110__89_, s_r_110__88_, s_r_110__87_, s_r_110__86_, s_r_110__85_, s_r_110__84_, s_r_110__83_, s_r_110__82_, s_r_110__81_, s_r_110__80_, s_r_110__79_, s_r_110__78_, s_r_110__77_, s_r_110__76_, s_r_110__75_, s_r_110__74_, s_r_110__73_, s_r_110__72_, s_r_110__71_, s_r_110__70_, s_r_110__69_, s_r_110__68_, s_r_110__67_, s_r_110__66_, s_r_110__65_, s_r_110__64_, s_r_110__63_, s_r_110__62_, s_r_110__61_, s_r_110__60_, s_r_110__59_, s_r_110__58_, s_r_110__57_, s_r_110__56_, s_r_110__55_, s_r_110__54_, s_r_110__53_, s_r_110__52_, s_r_110__51_, s_r_110__50_, s_r_110__49_, s_r_110__48_, s_r_110__47_, s_r_110__46_, s_r_110__45_, s_r_110__44_, s_r_110__43_, s_r_110__42_, s_r_110__41_, s_r_110__40_, s_r_110__39_, s_r_110__38_, s_r_110__37_, s_r_110__36_, s_r_110__35_, s_r_110__34_, s_r_110__33_, s_r_110__32_, s_r_110__31_, s_r_110__30_, s_r_110__29_, s_r_110__28_, s_r_110__27_, s_r_110__26_, s_r_110__25_, s_r_110__24_, s_r_110__23_, s_r_110__22_, s_r_110__21_, s_r_110__20_, s_r_110__19_, s_r_110__18_, s_r_110__17_, s_r_110__16_, s_r_110__15_, s_r_110__14_, s_r_110__13_, s_r_110__12_, s_r_110__11_, s_r_110__10_, s_r_110__9_, s_r_110__8_, s_r_110__7_, s_r_110__6_, s_r_110__5_, s_r_110__4_, s_r_110__3_, s_r_110__2_, s_r_110__1_, s_r_110__0_ }),
    .c_o(c_r[110]),
    .prod_accum_o({ prod_accum_110__111_, prod_accum_110__110_, prod_accum_110__109_, prod_accum_110__108_, prod_accum_110__107_, prod_accum_110__106_, prod_accum_110__105_, prod_accum_110__104_, prod_accum_110__103_, prod_accum_110__102_, prod_accum_110__101_, prod_accum_110__100_, prod_accum_110__99_, prod_accum_110__98_, prod_accum_110__97_, prod_accum_110__96_, prod_accum_110__95_, prod_accum_110__94_, prod_accum_110__93_, prod_accum_110__92_, prod_accum_110__91_, prod_accum_110__90_, prod_accum_110__89_, prod_accum_110__88_, prod_accum_110__87_, prod_accum_110__86_, prod_accum_110__85_, prod_accum_110__84_, prod_accum_110__83_, prod_accum_110__82_, prod_accum_110__81_, prod_accum_110__80_, prod_accum_110__79_, prod_accum_110__78_, prod_accum_110__77_, prod_accum_110__76_, prod_accum_110__75_, prod_accum_110__74_, prod_accum_110__73_, prod_accum_110__72_, prod_accum_110__71_, prod_accum_110__70_, prod_accum_110__69_, prod_accum_110__68_, prod_accum_110__67_, prod_accum_110__66_, prod_accum_110__65_, prod_accum_110__64_, prod_accum_110__63_, prod_accum_110__62_, prod_accum_110__61_, prod_accum_110__60_, prod_accum_110__59_, prod_accum_110__58_, prod_accum_110__57_, prod_accum_110__56_, prod_accum_110__55_, prod_accum_110__54_, prod_accum_110__53_, prod_accum_110__52_, prod_accum_110__51_, prod_accum_110__50_, prod_accum_110__49_, prod_accum_110__48_, prod_accum_110__47_, prod_accum_110__46_, prod_accum_110__45_, prod_accum_110__44_, prod_accum_110__43_, prod_accum_110__42_, prod_accum_110__41_, prod_accum_110__40_, prod_accum_110__39_, prod_accum_110__38_, prod_accum_110__37_, prod_accum_110__36_, prod_accum_110__35_, prod_accum_110__34_, prod_accum_110__33_, prod_accum_110__32_, prod_accum_110__31_, prod_accum_110__30_, prod_accum_110__29_, prod_accum_110__28_, prod_accum_110__27_, prod_accum_110__26_, prod_accum_110__25_, prod_accum_110__24_, prod_accum_110__23_, prod_accum_110__22_, prod_accum_110__21_, prod_accum_110__20_, prod_accum_110__19_, prod_accum_110__18_, prod_accum_110__17_, prod_accum_110__16_, prod_accum_110__15_, prod_accum_110__14_, prod_accum_110__13_, prod_accum_110__12_, prod_accum_110__11_, prod_accum_110__10_, prod_accum_110__9_, prod_accum_110__8_, prod_accum_110__7_, prod_accum_110__6_, prod_accum_110__5_, prod_accum_110__4_, prod_accum_110__3_, prod_accum_110__2_, prod_accum_110__1_, prod_accum_110__0_ })
  );


  bsg_mul_array_row_128_111_x
  genblk1_111__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[14207:14080]),
    .b_i(b_r[14207:14080]),
    .s_i({ s_r_110__127_, s_r_110__126_, s_r_110__125_, s_r_110__124_, s_r_110__123_, s_r_110__122_, s_r_110__121_, s_r_110__120_, s_r_110__119_, s_r_110__118_, s_r_110__117_, s_r_110__116_, s_r_110__115_, s_r_110__114_, s_r_110__113_, s_r_110__112_, s_r_110__111_, s_r_110__110_, s_r_110__109_, s_r_110__108_, s_r_110__107_, s_r_110__106_, s_r_110__105_, s_r_110__104_, s_r_110__103_, s_r_110__102_, s_r_110__101_, s_r_110__100_, s_r_110__99_, s_r_110__98_, s_r_110__97_, s_r_110__96_, s_r_110__95_, s_r_110__94_, s_r_110__93_, s_r_110__92_, s_r_110__91_, s_r_110__90_, s_r_110__89_, s_r_110__88_, s_r_110__87_, s_r_110__86_, s_r_110__85_, s_r_110__84_, s_r_110__83_, s_r_110__82_, s_r_110__81_, s_r_110__80_, s_r_110__79_, s_r_110__78_, s_r_110__77_, s_r_110__76_, s_r_110__75_, s_r_110__74_, s_r_110__73_, s_r_110__72_, s_r_110__71_, s_r_110__70_, s_r_110__69_, s_r_110__68_, s_r_110__67_, s_r_110__66_, s_r_110__65_, s_r_110__64_, s_r_110__63_, s_r_110__62_, s_r_110__61_, s_r_110__60_, s_r_110__59_, s_r_110__58_, s_r_110__57_, s_r_110__56_, s_r_110__55_, s_r_110__54_, s_r_110__53_, s_r_110__52_, s_r_110__51_, s_r_110__50_, s_r_110__49_, s_r_110__48_, s_r_110__47_, s_r_110__46_, s_r_110__45_, s_r_110__44_, s_r_110__43_, s_r_110__42_, s_r_110__41_, s_r_110__40_, s_r_110__39_, s_r_110__38_, s_r_110__37_, s_r_110__36_, s_r_110__35_, s_r_110__34_, s_r_110__33_, s_r_110__32_, s_r_110__31_, s_r_110__30_, s_r_110__29_, s_r_110__28_, s_r_110__27_, s_r_110__26_, s_r_110__25_, s_r_110__24_, s_r_110__23_, s_r_110__22_, s_r_110__21_, s_r_110__20_, s_r_110__19_, s_r_110__18_, s_r_110__17_, s_r_110__16_, s_r_110__15_, s_r_110__14_, s_r_110__13_, s_r_110__12_, s_r_110__11_, s_r_110__10_, s_r_110__9_, s_r_110__8_, s_r_110__7_, s_r_110__6_, s_r_110__5_, s_r_110__4_, s_r_110__3_, s_r_110__2_, s_r_110__1_, s_r_110__0_ }),
    .c_i(c_r[110]),
    .prod_accum_i({ prod_accum_110__111_, prod_accum_110__110_, prod_accum_110__109_, prod_accum_110__108_, prod_accum_110__107_, prod_accum_110__106_, prod_accum_110__105_, prod_accum_110__104_, prod_accum_110__103_, prod_accum_110__102_, prod_accum_110__101_, prod_accum_110__100_, prod_accum_110__99_, prod_accum_110__98_, prod_accum_110__97_, prod_accum_110__96_, prod_accum_110__95_, prod_accum_110__94_, prod_accum_110__93_, prod_accum_110__92_, prod_accum_110__91_, prod_accum_110__90_, prod_accum_110__89_, prod_accum_110__88_, prod_accum_110__87_, prod_accum_110__86_, prod_accum_110__85_, prod_accum_110__84_, prod_accum_110__83_, prod_accum_110__82_, prod_accum_110__81_, prod_accum_110__80_, prod_accum_110__79_, prod_accum_110__78_, prod_accum_110__77_, prod_accum_110__76_, prod_accum_110__75_, prod_accum_110__74_, prod_accum_110__73_, prod_accum_110__72_, prod_accum_110__71_, prod_accum_110__70_, prod_accum_110__69_, prod_accum_110__68_, prod_accum_110__67_, prod_accum_110__66_, prod_accum_110__65_, prod_accum_110__64_, prod_accum_110__63_, prod_accum_110__62_, prod_accum_110__61_, prod_accum_110__60_, prod_accum_110__59_, prod_accum_110__58_, prod_accum_110__57_, prod_accum_110__56_, prod_accum_110__55_, prod_accum_110__54_, prod_accum_110__53_, prod_accum_110__52_, prod_accum_110__51_, prod_accum_110__50_, prod_accum_110__49_, prod_accum_110__48_, prod_accum_110__47_, prod_accum_110__46_, prod_accum_110__45_, prod_accum_110__44_, prod_accum_110__43_, prod_accum_110__42_, prod_accum_110__41_, prod_accum_110__40_, prod_accum_110__39_, prod_accum_110__38_, prod_accum_110__37_, prod_accum_110__36_, prod_accum_110__35_, prod_accum_110__34_, prod_accum_110__33_, prod_accum_110__32_, prod_accum_110__31_, prod_accum_110__30_, prod_accum_110__29_, prod_accum_110__28_, prod_accum_110__27_, prod_accum_110__26_, prod_accum_110__25_, prod_accum_110__24_, prod_accum_110__23_, prod_accum_110__22_, prod_accum_110__21_, prod_accum_110__20_, prod_accum_110__19_, prod_accum_110__18_, prod_accum_110__17_, prod_accum_110__16_, prod_accum_110__15_, prod_accum_110__14_, prod_accum_110__13_, prod_accum_110__12_, prod_accum_110__11_, prod_accum_110__10_, prod_accum_110__9_, prod_accum_110__8_, prod_accum_110__7_, prod_accum_110__6_, prod_accum_110__5_, prod_accum_110__4_, prod_accum_110__3_, prod_accum_110__2_, prod_accum_110__1_, prod_accum_110__0_ }),
    .a_o(a_r[14335:14208]),
    .b_o(b_r[14335:14208]),
    .s_o({ s_r_111__127_, s_r_111__126_, s_r_111__125_, s_r_111__124_, s_r_111__123_, s_r_111__122_, s_r_111__121_, s_r_111__120_, s_r_111__119_, s_r_111__118_, s_r_111__117_, s_r_111__116_, s_r_111__115_, s_r_111__114_, s_r_111__113_, s_r_111__112_, s_r_111__111_, s_r_111__110_, s_r_111__109_, s_r_111__108_, s_r_111__107_, s_r_111__106_, s_r_111__105_, s_r_111__104_, s_r_111__103_, s_r_111__102_, s_r_111__101_, s_r_111__100_, s_r_111__99_, s_r_111__98_, s_r_111__97_, s_r_111__96_, s_r_111__95_, s_r_111__94_, s_r_111__93_, s_r_111__92_, s_r_111__91_, s_r_111__90_, s_r_111__89_, s_r_111__88_, s_r_111__87_, s_r_111__86_, s_r_111__85_, s_r_111__84_, s_r_111__83_, s_r_111__82_, s_r_111__81_, s_r_111__80_, s_r_111__79_, s_r_111__78_, s_r_111__77_, s_r_111__76_, s_r_111__75_, s_r_111__74_, s_r_111__73_, s_r_111__72_, s_r_111__71_, s_r_111__70_, s_r_111__69_, s_r_111__68_, s_r_111__67_, s_r_111__66_, s_r_111__65_, s_r_111__64_, s_r_111__63_, s_r_111__62_, s_r_111__61_, s_r_111__60_, s_r_111__59_, s_r_111__58_, s_r_111__57_, s_r_111__56_, s_r_111__55_, s_r_111__54_, s_r_111__53_, s_r_111__52_, s_r_111__51_, s_r_111__50_, s_r_111__49_, s_r_111__48_, s_r_111__47_, s_r_111__46_, s_r_111__45_, s_r_111__44_, s_r_111__43_, s_r_111__42_, s_r_111__41_, s_r_111__40_, s_r_111__39_, s_r_111__38_, s_r_111__37_, s_r_111__36_, s_r_111__35_, s_r_111__34_, s_r_111__33_, s_r_111__32_, s_r_111__31_, s_r_111__30_, s_r_111__29_, s_r_111__28_, s_r_111__27_, s_r_111__26_, s_r_111__25_, s_r_111__24_, s_r_111__23_, s_r_111__22_, s_r_111__21_, s_r_111__20_, s_r_111__19_, s_r_111__18_, s_r_111__17_, s_r_111__16_, s_r_111__15_, s_r_111__14_, s_r_111__13_, s_r_111__12_, s_r_111__11_, s_r_111__10_, s_r_111__9_, s_r_111__8_, s_r_111__7_, s_r_111__6_, s_r_111__5_, s_r_111__4_, s_r_111__3_, s_r_111__2_, s_r_111__1_, s_r_111__0_ }),
    .c_o(c_r[111]),
    .prod_accum_o({ prod_accum_111__112_, prod_accum_111__111_, prod_accum_111__110_, prod_accum_111__109_, prod_accum_111__108_, prod_accum_111__107_, prod_accum_111__106_, prod_accum_111__105_, prod_accum_111__104_, prod_accum_111__103_, prod_accum_111__102_, prod_accum_111__101_, prod_accum_111__100_, prod_accum_111__99_, prod_accum_111__98_, prod_accum_111__97_, prod_accum_111__96_, prod_accum_111__95_, prod_accum_111__94_, prod_accum_111__93_, prod_accum_111__92_, prod_accum_111__91_, prod_accum_111__90_, prod_accum_111__89_, prod_accum_111__88_, prod_accum_111__87_, prod_accum_111__86_, prod_accum_111__85_, prod_accum_111__84_, prod_accum_111__83_, prod_accum_111__82_, prod_accum_111__81_, prod_accum_111__80_, prod_accum_111__79_, prod_accum_111__78_, prod_accum_111__77_, prod_accum_111__76_, prod_accum_111__75_, prod_accum_111__74_, prod_accum_111__73_, prod_accum_111__72_, prod_accum_111__71_, prod_accum_111__70_, prod_accum_111__69_, prod_accum_111__68_, prod_accum_111__67_, prod_accum_111__66_, prod_accum_111__65_, prod_accum_111__64_, prod_accum_111__63_, prod_accum_111__62_, prod_accum_111__61_, prod_accum_111__60_, prod_accum_111__59_, prod_accum_111__58_, prod_accum_111__57_, prod_accum_111__56_, prod_accum_111__55_, prod_accum_111__54_, prod_accum_111__53_, prod_accum_111__52_, prod_accum_111__51_, prod_accum_111__50_, prod_accum_111__49_, prod_accum_111__48_, prod_accum_111__47_, prod_accum_111__46_, prod_accum_111__45_, prod_accum_111__44_, prod_accum_111__43_, prod_accum_111__42_, prod_accum_111__41_, prod_accum_111__40_, prod_accum_111__39_, prod_accum_111__38_, prod_accum_111__37_, prod_accum_111__36_, prod_accum_111__35_, prod_accum_111__34_, prod_accum_111__33_, prod_accum_111__32_, prod_accum_111__31_, prod_accum_111__30_, prod_accum_111__29_, prod_accum_111__28_, prod_accum_111__27_, prod_accum_111__26_, prod_accum_111__25_, prod_accum_111__24_, prod_accum_111__23_, prod_accum_111__22_, prod_accum_111__21_, prod_accum_111__20_, prod_accum_111__19_, prod_accum_111__18_, prod_accum_111__17_, prod_accum_111__16_, prod_accum_111__15_, prod_accum_111__14_, prod_accum_111__13_, prod_accum_111__12_, prod_accum_111__11_, prod_accum_111__10_, prod_accum_111__9_, prod_accum_111__8_, prod_accum_111__7_, prod_accum_111__6_, prod_accum_111__5_, prod_accum_111__4_, prod_accum_111__3_, prod_accum_111__2_, prod_accum_111__1_, prod_accum_111__0_ })
  );


  bsg_mul_array_row_128_112_x
  genblk1_112__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[14335:14208]),
    .b_i(b_r[14335:14208]),
    .s_i({ s_r_111__127_, s_r_111__126_, s_r_111__125_, s_r_111__124_, s_r_111__123_, s_r_111__122_, s_r_111__121_, s_r_111__120_, s_r_111__119_, s_r_111__118_, s_r_111__117_, s_r_111__116_, s_r_111__115_, s_r_111__114_, s_r_111__113_, s_r_111__112_, s_r_111__111_, s_r_111__110_, s_r_111__109_, s_r_111__108_, s_r_111__107_, s_r_111__106_, s_r_111__105_, s_r_111__104_, s_r_111__103_, s_r_111__102_, s_r_111__101_, s_r_111__100_, s_r_111__99_, s_r_111__98_, s_r_111__97_, s_r_111__96_, s_r_111__95_, s_r_111__94_, s_r_111__93_, s_r_111__92_, s_r_111__91_, s_r_111__90_, s_r_111__89_, s_r_111__88_, s_r_111__87_, s_r_111__86_, s_r_111__85_, s_r_111__84_, s_r_111__83_, s_r_111__82_, s_r_111__81_, s_r_111__80_, s_r_111__79_, s_r_111__78_, s_r_111__77_, s_r_111__76_, s_r_111__75_, s_r_111__74_, s_r_111__73_, s_r_111__72_, s_r_111__71_, s_r_111__70_, s_r_111__69_, s_r_111__68_, s_r_111__67_, s_r_111__66_, s_r_111__65_, s_r_111__64_, s_r_111__63_, s_r_111__62_, s_r_111__61_, s_r_111__60_, s_r_111__59_, s_r_111__58_, s_r_111__57_, s_r_111__56_, s_r_111__55_, s_r_111__54_, s_r_111__53_, s_r_111__52_, s_r_111__51_, s_r_111__50_, s_r_111__49_, s_r_111__48_, s_r_111__47_, s_r_111__46_, s_r_111__45_, s_r_111__44_, s_r_111__43_, s_r_111__42_, s_r_111__41_, s_r_111__40_, s_r_111__39_, s_r_111__38_, s_r_111__37_, s_r_111__36_, s_r_111__35_, s_r_111__34_, s_r_111__33_, s_r_111__32_, s_r_111__31_, s_r_111__30_, s_r_111__29_, s_r_111__28_, s_r_111__27_, s_r_111__26_, s_r_111__25_, s_r_111__24_, s_r_111__23_, s_r_111__22_, s_r_111__21_, s_r_111__20_, s_r_111__19_, s_r_111__18_, s_r_111__17_, s_r_111__16_, s_r_111__15_, s_r_111__14_, s_r_111__13_, s_r_111__12_, s_r_111__11_, s_r_111__10_, s_r_111__9_, s_r_111__8_, s_r_111__7_, s_r_111__6_, s_r_111__5_, s_r_111__4_, s_r_111__3_, s_r_111__2_, s_r_111__1_, s_r_111__0_ }),
    .c_i(c_r[111]),
    .prod_accum_i({ prod_accum_111__112_, prod_accum_111__111_, prod_accum_111__110_, prod_accum_111__109_, prod_accum_111__108_, prod_accum_111__107_, prod_accum_111__106_, prod_accum_111__105_, prod_accum_111__104_, prod_accum_111__103_, prod_accum_111__102_, prod_accum_111__101_, prod_accum_111__100_, prod_accum_111__99_, prod_accum_111__98_, prod_accum_111__97_, prod_accum_111__96_, prod_accum_111__95_, prod_accum_111__94_, prod_accum_111__93_, prod_accum_111__92_, prod_accum_111__91_, prod_accum_111__90_, prod_accum_111__89_, prod_accum_111__88_, prod_accum_111__87_, prod_accum_111__86_, prod_accum_111__85_, prod_accum_111__84_, prod_accum_111__83_, prod_accum_111__82_, prod_accum_111__81_, prod_accum_111__80_, prod_accum_111__79_, prod_accum_111__78_, prod_accum_111__77_, prod_accum_111__76_, prod_accum_111__75_, prod_accum_111__74_, prod_accum_111__73_, prod_accum_111__72_, prod_accum_111__71_, prod_accum_111__70_, prod_accum_111__69_, prod_accum_111__68_, prod_accum_111__67_, prod_accum_111__66_, prod_accum_111__65_, prod_accum_111__64_, prod_accum_111__63_, prod_accum_111__62_, prod_accum_111__61_, prod_accum_111__60_, prod_accum_111__59_, prod_accum_111__58_, prod_accum_111__57_, prod_accum_111__56_, prod_accum_111__55_, prod_accum_111__54_, prod_accum_111__53_, prod_accum_111__52_, prod_accum_111__51_, prod_accum_111__50_, prod_accum_111__49_, prod_accum_111__48_, prod_accum_111__47_, prod_accum_111__46_, prod_accum_111__45_, prod_accum_111__44_, prod_accum_111__43_, prod_accum_111__42_, prod_accum_111__41_, prod_accum_111__40_, prod_accum_111__39_, prod_accum_111__38_, prod_accum_111__37_, prod_accum_111__36_, prod_accum_111__35_, prod_accum_111__34_, prod_accum_111__33_, prod_accum_111__32_, prod_accum_111__31_, prod_accum_111__30_, prod_accum_111__29_, prod_accum_111__28_, prod_accum_111__27_, prod_accum_111__26_, prod_accum_111__25_, prod_accum_111__24_, prod_accum_111__23_, prod_accum_111__22_, prod_accum_111__21_, prod_accum_111__20_, prod_accum_111__19_, prod_accum_111__18_, prod_accum_111__17_, prod_accum_111__16_, prod_accum_111__15_, prod_accum_111__14_, prod_accum_111__13_, prod_accum_111__12_, prod_accum_111__11_, prod_accum_111__10_, prod_accum_111__9_, prod_accum_111__8_, prod_accum_111__7_, prod_accum_111__6_, prod_accum_111__5_, prod_accum_111__4_, prod_accum_111__3_, prod_accum_111__2_, prod_accum_111__1_, prod_accum_111__0_ }),
    .a_o(a_r[14463:14336]),
    .b_o(b_r[14463:14336]),
    .s_o({ s_r_112__127_, s_r_112__126_, s_r_112__125_, s_r_112__124_, s_r_112__123_, s_r_112__122_, s_r_112__121_, s_r_112__120_, s_r_112__119_, s_r_112__118_, s_r_112__117_, s_r_112__116_, s_r_112__115_, s_r_112__114_, s_r_112__113_, s_r_112__112_, s_r_112__111_, s_r_112__110_, s_r_112__109_, s_r_112__108_, s_r_112__107_, s_r_112__106_, s_r_112__105_, s_r_112__104_, s_r_112__103_, s_r_112__102_, s_r_112__101_, s_r_112__100_, s_r_112__99_, s_r_112__98_, s_r_112__97_, s_r_112__96_, s_r_112__95_, s_r_112__94_, s_r_112__93_, s_r_112__92_, s_r_112__91_, s_r_112__90_, s_r_112__89_, s_r_112__88_, s_r_112__87_, s_r_112__86_, s_r_112__85_, s_r_112__84_, s_r_112__83_, s_r_112__82_, s_r_112__81_, s_r_112__80_, s_r_112__79_, s_r_112__78_, s_r_112__77_, s_r_112__76_, s_r_112__75_, s_r_112__74_, s_r_112__73_, s_r_112__72_, s_r_112__71_, s_r_112__70_, s_r_112__69_, s_r_112__68_, s_r_112__67_, s_r_112__66_, s_r_112__65_, s_r_112__64_, s_r_112__63_, s_r_112__62_, s_r_112__61_, s_r_112__60_, s_r_112__59_, s_r_112__58_, s_r_112__57_, s_r_112__56_, s_r_112__55_, s_r_112__54_, s_r_112__53_, s_r_112__52_, s_r_112__51_, s_r_112__50_, s_r_112__49_, s_r_112__48_, s_r_112__47_, s_r_112__46_, s_r_112__45_, s_r_112__44_, s_r_112__43_, s_r_112__42_, s_r_112__41_, s_r_112__40_, s_r_112__39_, s_r_112__38_, s_r_112__37_, s_r_112__36_, s_r_112__35_, s_r_112__34_, s_r_112__33_, s_r_112__32_, s_r_112__31_, s_r_112__30_, s_r_112__29_, s_r_112__28_, s_r_112__27_, s_r_112__26_, s_r_112__25_, s_r_112__24_, s_r_112__23_, s_r_112__22_, s_r_112__21_, s_r_112__20_, s_r_112__19_, s_r_112__18_, s_r_112__17_, s_r_112__16_, s_r_112__15_, s_r_112__14_, s_r_112__13_, s_r_112__12_, s_r_112__11_, s_r_112__10_, s_r_112__9_, s_r_112__8_, s_r_112__7_, s_r_112__6_, s_r_112__5_, s_r_112__4_, s_r_112__3_, s_r_112__2_, s_r_112__1_, s_r_112__0_ }),
    .c_o(c_r[112]),
    .prod_accum_o({ prod_accum_112__113_, prod_accum_112__112_, prod_accum_112__111_, prod_accum_112__110_, prod_accum_112__109_, prod_accum_112__108_, prod_accum_112__107_, prod_accum_112__106_, prod_accum_112__105_, prod_accum_112__104_, prod_accum_112__103_, prod_accum_112__102_, prod_accum_112__101_, prod_accum_112__100_, prod_accum_112__99_, prod_accum_112__98_, prod_accum_112__97_, prod_accum_112__96_, prod_accum_112__95_, prod_accum_112__94_, prod_accum_112__93_, prod_accum_112__92_, prod_accum_112__91_, prod_accum_112__90_, prod_accum_112__89_, prod_accum_112__88_, prod_accum_112__87_, prod_accum_112__86_, prod_accum_112__85_, prod_accum_112__84_, prod_accum_112__83_, prod_accum_112__82_, prod_accum_112__81_, prod_accum_112__80_, prod_accum_112__79_, prod_accum_112__78_, prod_accum_112__77_, prod_accum_112__76_, prod_accum_112__75_, prod_accum_112__74_, prod_accum_112__73_, prod_accum_112__72_, prod_accum_112__71_, prod_accum_112__70_, prod_accum_112__69_, prod_accum_112__68_, prod_accum_112__67_, prod_accum_112__66_, prod_accum_112__65_, prod_accum_112__64_, prod_accum_112__63_, prod_accum_112__62_, prod_accum_112__61_, prod_accum_112__60_, prod_accum_112__59_, prod_accum_112__58_, prod_accum_112__57_, prod_accum_112__56_, prod_accum_112__55_, prod_accum_112__54_, prod_accum_112__53_, prod_accum_112__52_, prod_accum_112__51_, prod_accum_112__50_, prod_accum_112__49_, prod_accum_112__48_, prod_accum_112__47_, prod_accum_112__46_, prod_accum_112__45_, prod_accum_112__44_, prod_accum_112__43_, prod_accum_112__42_, prod_accum_112__41_, prod_accum_112__40_, prod_accum_112__39_, prod_accum_112__38_, prod_accum_112__37_, prod_accum_112__36_, prod_accum_112__35_, prod_accum_112__34_, prod_accum_112__33_, prod_accum_112__32_, prod_accum_112__31_, prod_accum_112__30_, prod_accum_112__29_, prod_accum_112__28_, prod_accum_112__27_, prod_accum_112__26_, prod_accum_112__25_, prod_accum_112__24_, prod_accum_112__23_, prod_accum_112__22_, prod_accum_112__21_, prod_accum_112__20_, prod_accum_112__19_, prod_accum_112__18_, prod_accum_112__17_, prod_accum_112__16_, prod_accum_112__15_, prod_accum_112__14_, prod_accum_112__13_, prod_accum_112__12_, prod_accum_112__11_, prod_accum_112__10_, prod_accum_112__9_, prod_accum_112__8_, prod_accum_112__7_, prod_accum_112__6_, prod_accum_112__5_, prod_accum_112__4_, prod_accum_112__3_, prod_accum_112__2_, prod_accum_112__1_, prod_accum_112__0_ })
  );


  bsg_mul_array_row_128_113_x
  genblk1_113__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[14463:14336]),
    .b_i(b_r[14463:14336]),
    .s_i({ s_r_112__127_, s_r_112__126_, s_r_112__125_, s_r_112__124_, s_r_112__123_, s_r_112__122_, s_r_112__121_, s_r_112__120_, s_r_112__119_, s_r_112__118_, s_r_112__117_, s_r_112__116_, s_r_112__115_, s_r_112__114_, s_r_112__113_, s_r_112__112_, s_r_112__111_, s_r_112__110_, s_r_112__109_, s_r_112__108_, s_r_112__107_, s_r_112__106_, s_r_112__105_, s_r_112__104_, s_r_112__103_, s_r_112__102_, s_r_112__101_, s_r_112__100_, s_r_112__99_, s_r_112__98_, s_r_112__97_, s_r_112__96_, s_r_112__95_, s_r_112__94_, s_r_112__93_, s_r_112__92_, s_r_112__91_, s_r_112__90_, s_r_112__89_, s_r_112__88_, s_r_112__87_, s_r_112__86_, s_r_112__85_, s_r_112__84_, s_r_112__83_, s_r_112__82_, s_r_112__81_, s_r_112__80_, s_r_112__79_, s_r_112__78_, s_r_112__77_, s_r_112__76_, s_r_112__75_, s_r_112__74_, s_r_112__73_, s_r_112__72_, s_r_112__71_, s_r_112__70_, s_r_112__69_, s_r_112__68_, s_r_112__67_, s_r_112__66_, s_r_112__65_, s_r_112__64_, s_r_112__63_, s_r_112__62_, s_r_112__61_, s_r_112__60_, s_r_112__59_, s_r_112__58_, s_r_112__57_, s_r_112__56_, s_r_112__55_, s_r_112__54_, s_r_112__53_, s_r_112__52_, s_r_112__51_, s_r_112__50_, s_r_112__49_, s_r_112__48_, s_r_112__47_, s_r_112__46_, s_r_112__45_, s_r_112__44_, s_r_112__43_, s_r_112__42_, s_r_112__41_, s_r_112__40_, s_r_112__39_, s_r_112__38_, s_r_112__37_, s_r_112__36_, s_r_112__35_, s_r_112__34_, s_r_112__33_, s_r_112__32_, s_r_112__31_, s_r_112__30_, s_r_112__29_, s_r_112__28_, s_r_112__27_, s_r_112__26_, s_r_112__25_, s_r_112__24_, s_r_112__23_, s_r_112__22_, s_r_112__21_, s_r_112__20_, s_r_112__19_, s_r_112__18_, s_r_112__17_, s_r_112__16_, s_r_112__15_, s_r_112__14_, s_r_112__13_, s_r_112__12_, s_r_112__11_, s_r_112__10_, s_r_112__9_, s_r_112__8_, s_r_112__7_, s_r_112__6_, s_r_112__5_, s_r_112__4_, s_r_112__3_, s_r_112__2_, s_r_112__1_, s_r_112__0_ }),
    .c_i(c_r[112]),
    .prod_accum_i({ prod_accum_112__113_, prod_accum_112__112_, prod_accum_112__111_, prod_accum_112__110_, prod_accum_112__109_, prod_accum_112__108_, prod_accum_112__107_, prod_accum_112__106_, prod_accum_112__105_, prod_accum_112__104_, prod_accum_112__103_, prod_accum_112__102_, prod_accum_112__101_, prod_accum_112__100_, prod_accum_112__99_, prod_accum_112__98_, prod_accum_112__97_, prod_accum_112__96_, prod_accum_112__95_, prod_accum_112__94_, prod_accum_112__93_, prod_accum_112__92_, prod_accum_112__91_, prod_accum_112__90_, prod_accum_112__89_, prod_accum_112__88_, prod_accum_112__87_, prod_accum_112__86_, prod_accum_112__85_, prod_accum_112__84_, prod_accum_112__83_, prod_accum_112__82_, prod_accum_112__81_, prod_accum_112__80_, prod_accum_112__79_, prod_accum_112__78_, prod_accum_112__77_, prod_accum_112__76_, prod_accum_112__75_, prod_accum_112__74_, prod_accum_112__73_, prod_accum_112__72_, prod_accum_112__71_, prod_accum_112__70_, prod_accum_112__69_, prod_accum_112__68_, prod_accum_112__67_, prod_accum_112__66_, prod_accum_112__65_, prod_accum_112__64_, prod_accum_112__63_, prod_accum_112__62_, prod_accum_112__61_, prod_accum_112__60_, prod_accum_112__59_, prod_accum_112__58_, prod_accum_112__57_, prod_accum_112__56_, prod_accum_112__55_, prod_accum_112__54_, prod_accum_112__53_, prod_accum_112__52_, prod_accum_112__51_, prod_accum_112__50_, prod_accum_112__49_, prod_accum_112__48_, prod_accum_112__47_, prod_accum_112__46_, prod_accum_112__45_, prod_accum_112__44_, prod_accum_112__43_, prod_accum_112__42_, prod_accum_112__41_, prod_accum_112__40_, prod_accum_112__39_, prod_accum_112__38_, prod_accum_112__37_, prod_accum_112__36_, prod_accum_112__35_, prod_accum_112__34_, prod_accum_112__33_, prod_accum_112__32_, prod_accum_112__31_, prod_accum_112__30_, prod_accum_112__29_, prod_accum_112__28_, prod_accum_112__27_, prod_accum_112__26_, prod_accum_112__25_, prod_accum_112__24_, prod_accum_112__23_, prod_accum_112__22_, prod_accum_112__21_, prod_accum_112__20_, prod_accum_112__19_, prod_accum_112__18_, prod_accum_112__17_, prod_accum_112__16_, prod_accum_112__15_, prod_accum_112__14_, prod_accum_112__13_, prod_accum_112__12_, prod_accum_112__11_, prod_accum_112__10_, prod_accum_112__9_, prod_accum_112__8_, prod_accum_112__7_, prod_accum_112__6_, prod_accum_112__5_, prod_accum_112__4_, prod_accum_112__3_, prod_accum_112__2_, prod_accum_112__1_, prod_accum_112__0_ }),
    .a_o(a_r[14591:14464]),
    .b_o(b_r[14591:14464]),
    .s_o({ s_r_113__127_, s_r_113__126_, s_r_113__125_, s_r_113__124_, s_r_113__123_, s_r_113__122_, s_r_113__121_, s_r_113__120_, s_r_113__119_, s_r_113__118_, s_r_113__117_, s_r_113__116_, s_r_113__115_, s_r_113__114_, s_r_113__113_, s_r_113__112_, s_r_113__111_, s_r_113__110_, s_r_113__109_, s_r_113__108_, s_r_113__107_, s_r_113__106_, s_r_113__105_, s_r_113__104_, s_r_113__103_, s_r_113__102_, s_r_113__101_, s_r_113__100_, s_r_113__99_, s_r_113__98_, s_r_113__97_, s_r_113__96_, s_r_113__95_, s_r_113__94_, s_r_113__93_, s_r_113__92_, s_r_113__91_, s_r_113__90_, s_r_113__89_, s_r_113__88_, s_r_113__87_, s_r_113__86_, s_r_113__85_, s_r_113__84_, s_r_113__83_, s_r_113__82_, s_r_113__81_, s_r_113__80_, s_r_113__79_, s_r_113__78_, s_r_113__77_, s_r_113__76_, s_r_113__75_, s_r_113__74_, s_r_113__73_, s_r_113__72_, s_r_113__71_, s_r_113__70_, s_r_113__69_, s_r_113__68_, s_r_113__67_, s_r_113__66_, s_r_113__65_, s_r_113__64_, s_r_113__63_, s_r_113__62_, s_r_113__61_, s_r_113__60_, s_r_113__59_, s_r_113__58_, s_r_113__57_, s_r_113__56_, s_r_113__55_, s_r_113__54_, s_r_113__53_, s_r_113__52_, s_r_113__51_, s_r_113__50_, s_r_113__49_, s_r_113__48_, s_r_113__47_, s_r_113__46_, s_r_113__45_, s_r_113__44_, s_r_113__43_, s_r_113__42_, s_r_113__41_, s_r_113__40_, s_r_113__39_, s_r_113__38_, s_r_113__37_, s_r_113__36_, s_r_113__35_, s_r_113__34_, s_r_113__33_, s_r_113__32_, s_r_113__31_, s_r_113__30_, s_r_113__29_, s_r_113__28_, s_r_113__27_, s_r_113__26_, s_r_113__25_, s_r_113__24_, s_r_113__23_, s_r_113__22_, s_r_113__21_, s_r_113__20_, s_r_113__19_, s_r_113__18_, s_r_113__17_, s_r_113__16_, s_r_113__15_, s_r_113__14_, s_r_113__13_, s_r_113__12_, s_r_113__11_, s_r_113__10_, s_r_113__9_, s_r_113__8_, s_r_113__7_, s_r_113__6_, s_r_113__5_, s_r_113__4_, s_r_113__3_, s_r_113__2_, s_r_113__1_, s_r_113__0_ }),
    .c_o(c_r[113]),
    .prod_accum_o({ prod_accum_113__114_, prod_accum_113__113_, prod_accum_113__112_, prod_accum_113__111_, prod_accum_113__110_, prod_accum_113__109_, prod_accum_113__108_, prod_accum_113__107_, prod_accum_113__106_, prod_accum_113__105_, prod_accum_113__104_, prod_accum_113__103_, prod_accum_113__102_, prod_accum_113__101_, prod_accum_113__100_, prod_accum_113__99_, prod_accum_113__98_, prod_accum_113__97_, prod_accum_113__96_, prod_accum_113__95_, prod_accum_113__94_, prod_accum_113__93_, prod_accum_113__92_, prod_accum_113__91_, prod_accum_113__90_, prod_accum_113__89_, prod_accum_113__88_, prod_accum_113__87_, prod_accum_113__86_, prod_accum_113__85_, prod_accum_113__84_, prod_accum_113__83_, prod_accum_113__82_, prod_accum_113__81_, prod_accum_113__80_, prod_accum_113__79_, prod_accum_113__78_, prod_accum_113__77_, prod_accum_113__76_, prod_accum_113__75_, prod_accum_113__74_, prod_accum_113__73_, prod_accum_113__72_, prod_accum_113__71_, prod_accum_113__70_, prod_accum_113__69_, prod_accum_113__68_, prod_accum_113__67_, prod_accum_113__66_, prod_accum_113__65_, prod_accum_113__64_, prod_accum_113__63_, prod_accum_113__62_, prod_accum_113__61_, prod_accum_113__60_, prod_accum_113__59_, prod_accum_113__58_, prod_accum_113__57_, prod_accum_113__56_, prod_accum_113__55_, prod_accum_113__54_, prod_accum_113__53_, prod_accum_113__52_, prod_accum_113__51_, prod_accum_113__50_, prod_accum_113__49_, prod_accum_113__48_, prod_accum_113__47_, prod_accum_113__46_, prod_accum_113__45_, prod_accum_113__44_, prod_accum_113__43_, prod_accum_113__42_, prod_accum_113__41_, prod_accum_113__40_, prod_accum_113__39_, prod_accum_113__38_, prod_accum_113__37_, prod_accum_113__36_, prod_accum_113__35_, prod_accum_113__34_, prod_accum_113__33_, prod_accum_113__32_, prod_accum_113__31_, prod_accum_113__30_, prod_accum_113__29_, prod_accum_113__28_, prod_accum_113__27_, prod_accum_113__26_, prod_accum_113__25_, prod_accum_113__24_, prod_accum_113__23_, prod_accum_113__22_, prod_accum_113__21_, prod_accum_113__20_, prod_accum_113__19_, prod_accum_113__18_, prod_accum_113__17_, prod_accum_113__16_, prod_accum_113__15_, prod_accum_113__14_, prod_accum_113__13_, prod_accum_113__12_, prod_accum_113__11_, prod_accum_113__10_, prod_accum_113__9_, prod_accum_113__8_, prod_accum_113__7_, prod_accum_113__6_, prod_accum_113__5_, prod_accum_113__4_, prod_accum_113__3_, prod_accum_113__2_, prod_accum_113__1_, prod_accum_113__0_ })
  );


  bsg_mul_array_row_128_114_x
  genblk1_114__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[14591:14464]),
    .b_i(b_r[14591:14464]),
    .s_i({ s_r_113__127_, s_r_113__126_, s_r_113__125_, s_r_113__124_, s_r_113__123_, s_r_113__122_, s_r_113__121_, s_r_113__120_, s_r_113__119_, s_r_113__118_, s_r_113__117_, s_r_113__116_, s_r_113__115_, s_r_113__114_, s_r_113__113_, s_r_113__112_, s_r_113__111_, s_r_113__110_, s_r_113__109_, s_r_113__108_, s_r_113__107_, s_r_113__106_, s_r_113__105_, s_r_113__104_, s_r_113__103_, s_r_113__102_, s_r_113__101_, s_r_113__100_, s_r_113__99_, s_r_113__98_, s_r_113__97_, s_r_113__96_, s_r_113__95_, s_r_113__94_, s_r_113__93_, s_r_113__92_, s_r_113__91_, s_r_113__90_, s_r_113__89_, s_r_113__88_, s_r_113__87_, s_r_113__86_, s_r_113__85_, s_r_113__84_, s_r_113__83_, s_r_113__82_, s_r_113__81_, s_r_113__80_, s_r_113__79_, s_r_113__78_, s_r_113__77_, s_r_113__76_, s_r_113__75_, s_r_113__74_, s_r_113__73_, s_r_113__72_, s_r_113__71_, s_r_113__70_, s_r_113__69_, s_r_113__68_, s_r_113__67_, s_r_113__66_, s_r_113__65_, s_r_113__64_, s_r_113__63_, s_r_113__62_, s_r_113__61_, s_r_113__60_, s_r_113__59_, s_r_113__58_, s_r_113__57_, s_r_113__56_, s_r_113__55_, s_r_113__54_, s_r_113__53_, s_r_113__52_, s_r_113__51_, s_r_113__50_, s_r_113__49_, s_r_113__48_, s_r_113__47_, s_r_113__46_, s_r_113__45_, s_r_113__44_, s_r_113__43_, s_r_113__42_, s_r_113__41_, s_r_113__40_, s_r_113__39_, s_r_113__38_, s_r_113__37_, s_r_113__36_, s_r_113__35_, s_r_113__34_, s_r_113__33_, s_r_113__32_, s_r_113__31_, s_r_113__30_, s_r_113__29_, s_r_113__28_, s_r_113__27_, s_r_113__26_, s_r_113__25_, s_r_113__24_, s_r_113__23_, s_r_113__22_, s_r_113__21_, s_r_113__20_, s_r_113__19_, s_r_113__18_, s_r_113__17_, s_r_113__16_, s_r_113__15_, s_r_113__14_, s_r_113__13_, s_r_113__12_, s_r_113__11_, s_r_113__10_, s_r_113__9_, s_r_113__8_, s_r_113__7_, s_r_113__6_, s_r_113__5_, s_r_113__4_, s_r_113__3_, s_r_113__2_, s_r_113__1_, s_r_113__0_ }),
    .c_i(c_r[113]),
    .prod_accum_i({ prod_accum_113__114_, prod_accum_113__113_, prod_accum_113__112_, prod_accum_113__111_, prod_accum_113__110_, prod_accum_113__109_, prod_accum_113__108_, prod_accum_113__107_, prod_accum_113__106_, prod_accum_113__105_, prod_accum_113__104_, prod_accum_113__103_, prod_accum_113__102_, prod_accum_113__101_, prod_accum_113__100_, prod_accum_113__99_, prod_accum_113__98_, prod_accum_113__97_, prod_accum_113__96_, prod_accum_113__95_, prod_accum_113__94_, prod_accum_113__93_, prod_accum_113__92_, prod_accum_113__91_, prod_accum_113__90_, prod_accum_113__89_, prod_accum_113__88_, prod_accum_113__87_, prod_accum_113__86_, prod_accum_113__85_, prod_accum_113__84_, prod_accum_113__83_, prod_accum_113__82_, prod_accum_113__81_, prod_accum_113__80_, prod_accum_113__79_, prod_accum_113__78_, prod_accum_113__77_, prod_accum_113__76_, prod_accum_113__75_, prod_accum_113__74_, prod_accum_113__73_, prod_accum_113__72_, prod_accum_113__71_, prod_accum_113__70_, prod_accum_113__69_, prod_accum_113__68_, prod_accum_113__67_, prod_accum_113__66_, prod_accum_113__65_, prod_accum_113__64_, prod_accum_113__63_, prod_accum_113__62_, prod_accum_113__61_, prod_accum_113__60_, prod_accum_113__59_, prod_accum_113__58_, prod_accum_113__57_, prod_accum_113__56_, prod_accum_113__55_, prod_accum_113__54_, prod_accum_113__53_, prod_accum_113__52_, prod_accum_113__51_, prod_accum_113__50_, prod_accum_113__49_, prod_accum_113__48_, prod_accum_113__47_, prod_accum_113__46_, prod_accum_113__45_, prod_accum_113__44_, prod_accum_113__43_, prod_accum_113__42_, prod_accum_113__41_, prod_accum_113__40_, prod_accum_113__39_, prod_accum_113__38_, prod_accum_113__37_, prod_accum_113__36_, prod_accum_113__35_, prod_accum_113__34_, prod_accum_113__33_, prod_accum_113__32_, prod_accum_113__31_, prod_accum_113__30_, prod_accum_113__29_, prod_accum_113__28_, prod_accum_113__27_, prod_accum_113__26_, prod_accum_113__25_, prod_accum_113__24_, prod_accum_113__23_, prod_accum_113__22_, prod_accum_113__21_, prod_accum_113__20_, prod_accum_113__19_, prod_accum_113__18_, prod_accum_113__17_, prod_accum_113__16_, prod_accum_113__15_, prod_accum_113__14_, prod_accum_113__13_, prod_accum_113__12_, prod_accum_113__11_, prod_accum_113__10_, prod_accum_113__9_, prod_accum_113__8_, prod_accum_113__7_, prod_accum_113__6_, prod_accum_113__5_, prod_accum_113__4_, prod_accum_113__3_, prod_accum_113__2_, prod_accum_113__1_, prod_accum_113__0_ }),
    .a_o(a_r[14719:14592]),
    .b_o(b_r[14719:14592]),
    .s_o({ s_r_114__127_, s_r_114__126_, s_r_114__125_, s_r_114__124_, s_r_114__123_, s_r_114__122_, s_r_114__121_, s_r_114__120_, s_r_114__119_, s_r_114__118_, s_r_114__117_, s_r_114__116_, s_r_114__115_, s_r_114__114_, s_r_114__113_, s_r_114__112_, s_r_114__111_, s_r_114__110_, s_r_114__109_, s_r_114__108_, s_r_114__107_, s_r_114__106_, s_r_114__105_, s_r_114__104_, s_r_114__103_, s_r_114__102_, s_r_114__101_, s_r_114__100_, s_r_114__99_, s_r_114__98_, s_r_114__97_, s_r_114__96_, s_r_114__95_, s_r_114__94_, s_r_114__93_, s_r_114__92_, s_r_114__91_, s_r_114__90_, s_r_114__89_, s_r_114__88_, s_r_114__87_, s_r_114__86_, s_r_114__85_, s_r_114__84_, s_r_114__83_, s_r_114__82_, s_r_114__81_, s_r_114__80_, s_r_114__79_, s_r_114__78_, s_r_114__77_, s_r_114__76_, s_r_114__75_, s_r_114__74_, s_r_114__73_, s_r_114__72_, s_r_114__71_, s_r_114__70_, s_r_114__69_, s_r_114__68_, s_r_114__67_, s_r_114__66_, s_r_114__65_, s_r_114__64_, s_r_114__63_, s_r_114__62_, s_r_114__61_, s_r_114__60_, s_r_114__59_, s_r_114__58_, s_r_114__57_, s_r_114__56_, s_r_114__55_, s_r_114__54_, s_r_114__53_, s_r_114__52_, s_r_114__51_, s_r_114__50_, s_r_114__49_, s_r_114__48_, s_r_114__47_, s_r_114__46_, s_r_114__45_, s_r_114__44_, s_r_114__43_, s_r_114__42_, s_r_114__41_, s_r_114__40_, s_r_114__39_, s_r_114__38_, s_r_114__37_, s_r_114__36_, s_r_114__35_, s_r_114__34_, s_r_114__33_, s_r_114__32_, s_r_114__31_, s_r_114__30_, s_r_114__29_, s_r_114__28_, s_r_114__27_, s_r_114__26_, s_r_114__25_, s_r_114__24_, s_r_114__23_, s_r_114__22_, s_r_114__21_, s_r_114__20_, s_r_114__19_, s_r_114__18_, s_r_114__17_, s_r_114__16_, s_r_114__15_, s_r_114__14_, s_r_114__13_, s_r_114__12_, s_r_114__11_, s_r_114__10_, s_r_114__9_, s_r_114__8_, s_r_114__7_, s_r_114__6_, s_r_114__5_, s_r_114__4_, s_r_114__3_, s_r_114__2_, s_r_114__1_, s_r_114__0_ }),
    .c_o(c_r[114]),
    .prod_accum_o({ prod_accum_114__115_, prod_accum_114__114_, prod_accum_114__113_, prod_accum_114__112_, prod_accum_114__111_, prod_accum_114__110_, prod_accum_114__109_, prod_accum_114__108_, prod_accum_114__107_, prod_accum_114__106_, prod_accum_114__105_, prod_accum_114__104_, prod_accum_114__103_, prod_accum_114__102_, prod_accum_114__101_, prod_accum_114__100_, prod_accum_114__99_, prod_accum_114__98_, prod_accum_114__97_, prod_accum_114__96_, prod_accum_114__95_, prod_accum_114__94_, prod_accum_114__93_, prod_accum_114__92_, prod_accum_114__91_, prod_accum_114__90_, prod_accum_114__89_, prod_accum_114__88_, prod_accum_114__87_, prod_accum_114__86_, prod_accum_114__85_, prod_accum_114__84_, prod_accum_114__83_, prod_accum_114__82_, prod_accum_114__81_, prod_accum_114__80_, prod_accum_114__79_, prod_accum_114__78_, prod_accum_114__77_, prod_accum_114__76_, prod_accum_114__75_, prod_accum_114__74_, prod_accum_114__73_, prod_accum_114__72_, prod_accum_114__71_, prod_accum_114__70_, prod_accum_114__69_, prod_accum_114__68_, prod_accum_114__67_, prod_accum_114__66_, prod_accum_114__65_, prod_accum_114__64_, prod_accum_114__63_, prod_accum_114__62_, prod_accum_114__61_, prod_accum_114__60_, prod_accum_114__59_, prod_accum_114__58_, prod_accum_114__57_, prod_accum_114__56_, prod_accum_114__55_, prod_accum_114__54_, prod_accum_114__53_, prod_accum_114__52_, prod_accum_114__51_, prod_accum_114__50_, prod_accum_114__49_, prod_accum_114__48_, prod_accum_114__47_, prod_accum_114__46_, prod_accum_114__45_, prod_accum_114__44_, prod_accum_114__43_, prod_accum_114__42_, prod_accum_114__41_, prod_accum_114__40_, prod_accum_114__39_, prod_accum_114__38_, prod_accum_114__37_, prod_accum_114__36_, prod_accum_114__35_, prod_accum_114__34_, prod_accum_114__33_, prod_accum_114__32_, prod_accum_114__31_, prod_accum_114__30_, prod_accum_114__29_, prod_accum_114__28_, prod_accum_114__27_, prod_accum_114__26_, prod_accum_114__25_, prod_accum_114__24_, prod_accum_114__23_, prod_accum_114__22_, prod_accum_114__21_, prod_accum_114__20_, prod_accum_114__19_, prod_accum_114__18_, prod_accum_114__17_, prod_accum_114__16_, prod_accum_114__15_, prod_accum_114__14_, prod_accum_114__13_, prod_accum_114__12_, prod_accum_114__11_, prod_accum_114__10_, prod_accum_114__9_, prod_accum_114__8_, prod_accum_114__7_, prod_accum_114__6_, prod_accum_114__5_, prod_accum_114__4_, prod_accum_114__3_, prod_accum_114__2_, prod_accum_114__1_, prod_accum_114__0_ })
  );


  bsg_mul_array_row_128_115_x
  genblk1_115__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[14719:14592]),
    .b_i(b_r[14719:14592]),
    .s_i({ s_r_114__127_, s_r_114__126_, s_r_114__125_, s_r_114__124_, s_r_114__123_, s_r_114__122_, s_r_114__121_, s_r_114__120_, s_r_114__119_, s_r_114__118_, s_r_114__117_, s_r_114__116_, s_r_114__115_, s_r_114__114_, s_r_114__113_, s_r_114__112_, s_r_114__111_, s_r_114__110_, s_r_114__109_, s_r_114__108_, s_r_114__107_, s_r_114__106_, s_r_114__105_, s_r_114__104_, s_r_114__103_, s_r_114__102_, s_r_114__101_, s_r_114__100_, s_r_114__99_, s_r_114__98_, s_r_114__97_, s_r_114__96_, s_r_114__95_, s_r_114__94_, s_r_114__93_, s_r_114__92_, s_r_114__91_, s_r_114__90_, s_r_114__89_, s_r_114__88_, s_r_114__87_, s_r_114__86_, s_r_114__85_, s_r_114__84_, s_r_114__83_, s_r_114__82_, s_r_114__81_, s_r_114__80_, s_r_114__79_, s_r_114__78_, s_r_114__77_, s_r_114__76_, s_r_114__75_, s_r_114__74_, s_r_114__73_, s_r_114__72_, s_r_114__71_, s_r_114__70_, s_r_114__69_, s_r_114__68_, s_r_114__67_, s_r_114__66_, s_r_114__65_, s_r_114__64_, s_r_114__63_, s_r_114__62_, s_r_114__61_, s_r_114__60_, s_r_114__59_, s_r_114__58_, s_r_114__57_, s_r_114__56_, s_r_114__55_, s_r_114__54_, s_r_114__53_, s_r_114__52_, s_r_114__51_, s_r_114__50_, s_r_114__49_, s_r_114__48_, s_r_114__47_, s_r_114__46_, s_r_114__45_, s_r_114__44_, s_r_114__43_, s_r_114__42_, s_r_114__41_, s_r_114__40_, s_r_114__39_, s_r_114__38_, s_r_114__37_, s_r_114__36_, s_r_114__35_, s_r_114__34_, s_r_114__33_, s_r_114__32_, s_r_114__31_, s_r_114__30_, s_r_114__29_, s_r_114__28_, s_r_114__27_, s_r_114__26_, s_r_114__25_, s_r_114__24_, s_r_114__23_, s_r_114__22_, s_r_114__21_, s_r_114__20_, s_r_114__19_, s_r_114__18_, s_r_114__17_, s_r_114__16_, s_r_114__15_, s_r_114__14_, s_r_114__13_, s_r_114__12_, s_r_114__11_, s_r_114__10_, s_r_114__9_, s_r_114__8_, s_r_114__7_, s_r_114__6_, s_r_114__5_, s_r_114__4_, s_r_114__3_, s_r_114__2_, s_r_114__1_, s_r_114__0_ }),
    .c_i(c_r[114]),
    .prod_accum_i({ prod_accum_114__115_, prod_accum_114__114_, prod_accum_114__113_, prod_accum_114__112_, prod_accum_114__111_, prod_accum_114__110_, prod_accum_114__109_, prod_accum_114__108_, prod_accum_114__107_, prod_accum_114__106_, prod_accum_114__105_, prod_accum_114__104_, prod_accum_114__103_, prod_accum_114__102_, prod_accum_114__101_, prod_accum_114__100_, prod_accum_114__99_, prod_accum_114__98_, prod_accum_114__97_, prod_accum_114__96_, prod_accum_114__95_, prod_accum_114__94_, prod_accum_114__93_, prod_accum_114__92_, prod_accum_114__91_, prod_accum_114__90_, prod_accum_114__89_, prod_accum_114__88_, prod_accum_114__87_, prod_accum_114__86_, prod_accum_114__85_, prod_accum_114__84_, prod_accum_114__83_, prod_accum_114__82_, prod_accum_114__81_, prod_accum_114__80_, prod_accum_114__79_, prod_accum_114__78_, prod_accum_114__77_, prod_accum_114__76_, prod_accum_114__75_, prod_accum_114__74_, prod_accum_114__73_, prod_accum_114__72_, prod_accum_114__71_, prod_accum_114__70_, prod_accum_114__69_, prod_accum_114__68_, prod_accum_114__67_, prod_accum_114__66_, prod_accum_114__65_, prod_accum_114__64_, prod_accum_114__63_, prod_accum_114__62_, prod_accum_114__61_, prod_accum_114__60_, prod_accum_114__59_, prod_accum_114__58_, prod_accum_114__57_, prod_accum_114__56_, prod_accum_114__55_, prod_accum_114__54_, prod_accum_114__53_, prod_accum_114__52_, prod_accum_114__51_, prod_accum_114__50_, prod_accum_114__49_, prod_accum_114__48_, prod_accum_114__47_, prod_accum_114__46_, prod_accum_114__45_, prod_accum_114__44_, prod_accum_114__43_, prod_accum_114__42_, prod_accum_114__41_, prod_accum_114__40_, prod_accum_114__39_, prod_accum_114__38_, prod_accum_114__37_, prod_accum_114__36_, prod_accum_114__35_, prod_accum_114__34_, prod_accum_114__33_, prod_accum_114__32_, prod_accum_114__31_, prod_accum_114__30_, prod_accum_114__29_, prod_accum_114__28_, prod_accum_114__27_, prod_accum_114__26_, prod_accum_114__25_, prod_accum_114__24_, prod_accum_114__23_, prod_accum_114__22_, prod_accum_114__21_, prod_accum_114__20_, prod_accum_114__19_, prod_accum_114__18_, prod_accum_114__17_, prod_accum_114__16_, prod_accum_114__15_, prod_accum_114__14_, prod_accum_114__13_, prod_accum_114__12_, prod_accum_114__11_, prod_accum_114__10_, prod_accum_114__9_, prod_accum_114__8_, prod_accum_114__7_, prod_accum_114__6_, prod_accum_114__5_, prod_accum_114__4_, prod_accum_114__3_, prod_accum_114__2_, prod_accum_114__1_, prod_accum_114__0_ }),
    .a_o(a_r[14847:14720]),
    .b_o(b_r[14847:14720]),
    .s_o({ s_r_115__127_, s_r_115__126_, s_r_115__125_, s_r_115__124_, s_r_115__123_, s_r_115__122_, s_r_115__121_, s_r_115__120_, s_r_115__119_, s_r_115__118_, s_r_115__117_, s_r_115__116_, s_r_115__115_, s_r_115__114_, s_r_115__113_, s_r_115__112_, s_r_115__111_, s_r_115__110_, s_r_115__109_, s_r_115__108_, s_r_115__107_, s_r_115__106_, s_r_115__105_, s_r_115__104_, s_r_115__103_, s_r_115__102_, s_r_115__101_, s_r_115__100_, s_r_115__99_, s_r_115__98_, s_r_115__97_, s_r_115__96_, s_r_115__95_, s_r_115__94_, s_r_115__93_, s_r_115__92_, s_r_115__91_, s_r_115__90_, s_r_115__89_, s_r_115__88_, s_r_115__87_, s_r_115__86_, s_r_115__85_, s_r_115__84_, s_r_115__83_, s_r_115__82_, s_r_115__81_, s_r_115__80_, s_r_115__79_, s_r_115__78_, s_r_115__77_, s_r_115__76_, s_r_115__75_, s_r_115__74_, s_r_115__73_, s_r_115__72_, s_r_115__71_, s_r_115__70_, s_r_115__69_, s_r_115__68_, s_r_115__67_, s_r_115__66_, s_r_115__65_, s_r_115__64_, s_r_115__63_, s_r_115__62_, s_r_115__61_, s_r_115__60_, s_r_115__59_, s_r_115__58_, s_r_115__57_, s_r_115__56_, s_r_115__55_, s_r_115__54_, s_r_115__53_, s_r_115__52_, s_r_115__51_, s_r_115__50_, s_r_115__49_, s_r_115__48_, s_r_115__47_, s_r_115__46_, s_r_115__45_, s_r_115__44_, s_r_115__43_, s_r_115__42_, s_r_115__41_, s_r_115__40_, s_r_115__39_, s_r_115__38_, s_r_115__37_, s_r_115__36_, s_r_115__35_, s_r_115__34_, s_r_115__33_, s_r_115__32_, s_r_115__31_, s_r_115__30_, s_r_115__29_, s_r_115__28_, s_r_115__27_, s_r_115__26_, s_r_115__25_, s_r_115__24_, s_r_115__23_, s_r_115__22_, s_r_115__21_, s_r_115__20_, s_r_115__19_, s_r_115__18_, s_r_115__17_, s_r_115__16_, s_r_115__15_, s_r_115__14_, s_r_115__13_, s_r_115__12_, s_r_115__11_, s_r_115__10_, s_r_115__9_, s_r_115__8_, s_r_115__7_, s_r_115__6_, s_r_115__5_, s_r_115__4_, s_r_115__3_, s_r_115__2_, s_r_115__1_, s_r_115__0_ }),
    .c_o(c_r[115]),
    .prod_accum_o({ prod_accum_115__116_, prod_accum_115__115_, prod_accum_115__114_, prod_accum_115__113_, prod_accum_115__112_, prod_accum_115__111_, prod_accum_115__110_, prod_accum_115__109_, prod_accum_115__108_, prod_accum_115__107_, prod_accum_115__106_, prod_accum_115__105_, prod_accum_115__104_, prod_accum_115__103_, prod_accum_115__102_, prod_accum_115__101_, prod_accum_115__100_, prod_accum_115__99_, prod_accum_115__98_, prod_accum_115__97_, prod_accum_115__96_, prod_accum_115__95_, prod_accum_115__94_, prod_accum_115__93_, prod_accum_115__92_, prod_accum_115__91_, prod_accum_115__90_, prod_accum_115__89_, prod_accum_115__88_, prod_accum_115__87_, prod_accum_115__86_, prod_accum_115__85_, prod_accum_115__84_, prod_accum_115__83_, prod_accum_115__82_, prod_accum_115__81_, prod_accum_115__80_, prod_accum_115__79_, prod_accum_115__78_, prod_accum_115__77_, prod_accum_115__76_, prod_accum_115__75_, prod_accum_115__74_, prod_accum_115__73_, prod_accum_115__72_, prod_accum_115__71_, prod_accum_115__70_, prod_accum_115__69_, prod_accum_115__68_, prod_accum_115__67_, prod_accum_115__66_, prod_accum_115__65_, prod_accum_115__64_, prod_accum_115__63_, prod_accum_115__62_, prod_accum_115__61_, prod_accum_115__60_, prod_accum_115__59_, prod_accum_115__58_, prod_accum_115__57_, prod_accum_115__56_, prod_accum_115__55_, prod_accum_115__54_, prod_accum_115__53_, prod_accum_115__52_, prod_accum_115__51_, prod_accum_115__50_, prod_accum_115__49_, prod_accum_115__48_, prod_accum_115__47_, prod_accum_115__46_, prod_accum_115__45_, prod_accum_115__44_, prod_accum_115__43_, prod_accum_115__42_, prod_accum_115__41_, prod_accum_115__40_, prod_accum_115__39_, prod_accum_115__38_, prod_accum_115__37_, prod_accum_115__36_, prod_accum_115__35_, prod_accum_115__34_, prod_accum_115__33_, prod_accum_115__32_, prod_accum_115__31_, prod_accum_115__30_, prod_accum_115__29_, prod_accum_115__28_, prod_accum_115__27_, prod_accum_115__26_, prod_accum_115__25_, prod_accum_115__24_, prod_accum_115__23_, prod_accum_115__22_, prod_accum_115__21_, prod_accum_115__20_, prod_accum_115__19_, prod_accum_115__18_, prod_accum_115__17_, prod_accum_115__16_, prod_accum_115__15_, prod_accum_115__14_, prod_accum_115__13_, prod_accum_115__12_, prod_accum_115__11_, prod_accum_115__10_, prod_accum_115__9_, prod_accum_115__8_, prod_accum_115__7_, prod_accum_115__6_, prod_accum_115__5_, prod_accum_115__4_, prod_accum_115__3_, prod_accum_115__2_, prod_accum_115__1_, prod_accum_115__0_ })
  );


  bsg_mul_array_row_128_116_x
  genblk1_116__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[14847:14720]),
    .b_i(b_r[14847:14720]),
    .s_i({ s_r_115__127_, s_r_115__126_, s_r_115__125_, s_r_115__124_, s_r_115__123_, s_r_115__122_, s_r_115__121_, s_r_115__120_, s_r_115__119_, s_r_115__118_, s_r_115__117_, s_r_115__116_, s_r_115__115_, s_r_115__114_, s_r_115__113_, s_r_115__112_, s_r_115__111_, s_r_115__110_, s_r_115__109_, s_r_115__108_, s_r_115__107_, s_r_115__106_, s_r_115__105_, s_r_115__104_, s_r_115__103_, s_r_115__102_, s_r_115__101_, s_r_115__100_, s_r_115__99_, s_r_115__98_, s_r_115__97_, s_r_115__96_, s_r_115__95_, s_r_115__94_, s_r_115__93_, s_r_115__92_, s_r_115__91_, s_r_115__90_, s_r_115__89_, s_r_115__88_, s_r_115__87_, s_r_115__86_, s_r_115__85_, s_r_115__84_, s_r_115__83_, s_r_115__82_, s_r_115__81_, s_r_115__80_, s_r_115__79_, s_r_115__78_, s_r_115__77_, s_r_115__76_, s_r_115__75_, s_r_115__74_, s_r_115__73_, s_r_115__72_, s_r_115__71_, s_r_115__70_, s_r_115__69_, s_r_115__68_, s_r_115__67_, s_r_115__66_, s_r_115__65_, s_r_115__64_, s_r_115__63_, s_r_115__62_, s_r_115__61_, s_r_115__60_, s_r_115__59_, s_r_115__58_, s_r_115__57_, s_r_115__56_, s_r_115__55_, s_r_115__54_, s_r_115__53_, s_r_115__52_, s_r_115__51_, s_r_115__50_, s_r_115__49_, s_r_115__48_, s_r_115__47_, s_r_115__46_, s_r_115__45_, s_r_115__44_, s_r_115__43_, s_r_115__42_, s_r_115__41_, s_r_115__40_, s_r_115__39_, s_r_115__38_, s_r_115__37_, s_r_115__36_, s_r_115__35_, s_r_115__34_, s_r_115__33_, s_r_115__32_, s_r_115__31_, s_r_115__30_, s_r_115__29_, s_r_115__28_, s_r_115__27_, s_r_115__26_, s_r_115__25_, s_r_115__24_, s_r_115__23_, s_r_115__22_, s_r_115__21_, s_r_115__20_, s_r_115__19_, s_r_115__18_, s_r_115__17_, s_r_115__16_, s_r_115__15_, s_r_115__14_, s_r_115__13_, s_r_115__12_, s_r_115__11_, s_r_115__10_, s_r_115__9_, s_r_115__8_, s_r_115__7_, s_r_115__6_, s_r_115__5_, s_r_115__4_, s_r_115__3_, s_r_115__2_, s_r_115__1_, s_r_115__0_ }),
    .c_i(c_r[115]),
    .prod_accum_i({ prod_accum_115__116_, prod_accum_115__115_, prod_accum_115__114_, prod_accum_115__113_, prod_accum_115__112_, prod_accum_115__111_, prod_accum_115__110_, prod_accum_115__109_, prod_accum_115__108_, prod_accum_115__107_, prod_accum_115__106_, prod_accum_115__105_, prod_accum_115__104_, prod_accum_115__103_, prod_accum_115__102_, prod_accum_115__101_, prod_accum_115__100_, prod_accum_115__99_, prod_accum_115__98_, prod_accum_115__97_, prod_accum_115__96_, prod_accum_115__95_, prod_accum_115__94_, prod_accum_115__93_, prod_accum_115__92_, prod_accum_115__91_, prod_accum_115__90_, prod_accum_115__89_, prod_accum_115__88_, prod_accum_115__87_, prod_accum_115__86_, prod_accum_115__85_, prod_accum_115__84_, prod_accum_115__83_, prod_accum_115__82_, prod_accum_115__81_, prod_accum_115__80_, prod_accum_115__79_, prod_accum_115__78_, prod_accum_115__77_, prod_accum_115__76_, prod_accum_115__75_, prod_accum_115__74_, prod_accum_115__73_, prod_accum_115__72_, prod_accum_115__71_, prod_accum_115__70_, prod_accum_115__69_, prod_accum_115__68_, prod_accum_115__67_, prod_accum_115__66_, prod_accum_115__65_, prod_accum_115__64_, prod_accum_115__63_, prod_accum_115__62_, prod_accum_115__61_, prod_accum_115__60_, prod_accum_115__59_, prod_accum_115__58_, prod_accum_115__57_, prod_accum_115__56_, prod_accum_115__55_, prod_accum_115__54_, prod_accum_115__53_, prod_accum_115__52_, prod_accum_115__51_, prod_accum_115__50_, prod_accum_115__49_, prod_accum_115__48_, prod_accum_115__47_, prod_accum_115__46_, prod_accum_115__45_, prod_accum_115__44_, prod_accum_115__43_, prod_accum_115__42_, prod_accum_115__41_, prod_accum_115__40_, prod_accum_115__39_, prod_accum_115__38_, prod_accum_115__37_, prod_accum_115__36_, prod_accum_115__35_, prod_accum_115__34_, prod_accum_115__33_, prod_accum_115__32_, prod_accum_115__31_, prod_accum_115__30_, prod_accum_115__29_, prod_accum_115__28_, prod_accum_115__27_, prod_accum_115__26_, prod_accum_115__25_, prod_accum_115__24_, prod_accum_115__23_, prod_accum_115__22_, prod_accum_115__21_, prod_accum_115__20_, prod_accum_115__19_, prod_accum_115__18_, prod_accum_115__17_, prod_accum_115__16_, prod_accum_115__15_, prod_accum_115__14_, prod_accum_115__13_, prod_accum_115__12_, prod_accum_115__11_, prod_accum_115__10_, prod_accum_115__9_, prod_accum_115__8_, prod_accum_115__7_, prod_accum_115__6_, prod_accum_115__5_, prod_accum_115__4_, prod_accum_115__3_, prod_accum_115__2_, prod_accum_115__1_, prod_accum_115__0_ }),
    .a_o(a_r[14975:14848]),
    .b_o(b_r[14975:14848]),
    .s_o({ s_r_116__127_, s_r_116__126_, s_r_116__125_, s_r_116__124_, s_r_116__123_, s_r_116__122_, s_r_116__121_, s_r_116__120_, s_r_116__119_, s_r_116__118_, s_r_116__117_, s_r_116__116_, s_r_116__115_, s_r_116__114_, s_r_116__113_, s_r_116__112_, s_r_116__111_, s_r_116__110_, s_r_116__109_, s_r_116__108_, s_r_116__107_, s_r_116__106_, s_r_116__105_, s_r_116__104_, s_r_116__103_, s_r_116__102_, s_r_116__101_, s_r_116__100_, s_r_116__99_, s_r_116__98_, s_r_116__97_, s_r_116__96_, s_r_116__95_, s_r_116__94_, s_r_116__93_, s_r_116__92_, s_r_116__91_, s_r_116__90_, s_r_116__89_, s_r_116__88_, s_r_116__87_, s_r_116__86_, s_r_116__85_, s_r_116__84_, s_r_116__83_, s_r_116__82_, s_r_116__81_, s_r_116__80_, s_r_116__79_, s_r_116__78_, s_r_116__77_, s_r_116__76_, s_r_116__75_, s_r_116__74_, s_r_116__73_, s_r_116__72_, s_r_116__71_, s_r_116__70_, s_r_116__69_, s_r_116__68_, s_r_116__67_, s_r_116__66_, s_r_116__65_, s_r_116__64_, s_r_116__63_, s_r_116__62_, s_r_116__61_, s_r_116__60_, s_r_116__59_, s_r_116__58_, s_r_116__57_, s_r_116__56_, s_r_116__55_, s_r_116__54_, s_r_116__53_, s_r_116__52_, s_r_116__51_, s_r_116__50_, s_r_116__49_, s_r_116__48_, s_r_116__47_, s_r_116__46_, s_r_116__45_, s_r_116__44_, s_r_116__43_, s_r_116__42_, s_r_116__41_, s_r_116__40_, s_r_116__39_, s_r_116__38_, s_r_116__37_, s_r_116__36_, s_r_116__35_, s_r_116__34_, s_r_116__33_, s_r_116__32_, s_r_116__31_, s_r_116__30_, s_r_116__29_, s_r_116__28_, s_r_116__27_, s_r_116__26_, s_r_116__25_, s_r_116__24_, s_r_116__23_, s_r_116__22_, s_r_116__21_, s_r_116__20_, s_r_116__19_, s_r_116__18_, s_r_116__17_, s_r_116__16_, s_r_116__15_, s_r_116__14_, s_r_116__13_, s_r_116__12_, s_r_116__11_, s_r_116__10_, s_r_116__9_, s_r_116__8_, s_r_116__7_, s_r_116__6_, s_r_116__5_, s_r_116__4_, s_r_116__3_, s_r_116__2_, s_r_116__1_, s_r_116__0_ }),
    .c_o(c_r[116]),
    .prod_accum_o({ prod_accum_116__117_, prod_accum_116__116_, prod_accum_116__115_, prod_accum_116__114_, prod_accum_116__113_, prod_accum_116__112_, prod_accum_116__111_, prod_accum_116__110_, prod_accum_116__109_, prod_accum_116__108_, prod_accum_116__107_, prod_accum_116__106_, prod_accum_116__105_, prod_accum_116__104_, prod_accum_116__103_, prod_accum_116__102_, prod_accum_116__101_, prod_accum_116__100_, prod_accum_116__99_, prod_accum_116__98_, prod_accum_116__97_, prod_accum_116__96_, prod_accum_116__95_, prod_accum_116__94_, prod_accum_116__93_, prod_accum_116__92_, prod_accum_116__91_, prod_accum_116__90_, prod_accum_116__89_, prod_accum_116__88_, prod_accum_116__87_, prod_accum_116__86_, prod_accum_116__85_, prod_accum_116__84_, prod_accum_116__83_, prod_accum_116__82_, prod_accum_116__81_, prod_accum_116__80_, prod_accum_116__79_, prod_accum_116__78_, prod_accum_116__77_, prod_accum_116__76_, prod_accum_116__75_, prod_accum_116__74_, prod_accum_116__73_, prod_accum_116__72_, prod_accum_116__71_, prod_accum_116__70_, prod_accum_116__69_, prod_accum_116__68_, prod_accum_116__67_, prod_accum_116__66_, prod_accum_116__65_, prod_accum_116__64_, prod_accum_116__63_, prod_accum_116__62_, prod_accum_116__61_, prod_accum_116__60_, prod_accum_116__59_, prod_accum_116__58_, prod_accum_116__57_, prod_accum_116__56_, prod_accum_116__55_, prod_accum_116__54_, prod_accum_116__53_, prod_accum_116__52_, prod_accum_116__51_, prod_accum_116__50_, prod_accum_116__49_, prod_accum_116__48_, prod_accum_116__47_, prod_accum_116__46_, prod_accum_116__45_, prod_accum_116__44_, prod_accum_116__43_, prod_accum_116__42_, prod_accum_116__41_, prod_accum_116__40_, prod_accum_116__39_, prod_accum_116__38_, prod_accum_116__37_, prod_accum_116__36_, prod_accum_116__35_, prod_accum_116__34_, prod_accum_116__33_, prod_accum_116__32_, prod_accum_116__31_, prod_accum_116__30_, prod_accum_116__29_, prod_accum_116__28_, prod_accum_116__27_, prod_accum_116__26_, prod_accum_116__25_, prod_accum_116__24_, prod_accum_116__23_, prod_accum_116__22_, prod_accum_116__21_, prod_accum_116__20_, prod_accum_116__19_, prod_accum_116__18_, prod_accum_116__17_, prod_accum_116__16_, prod_accum_116__15_, prod_accum_116__14_, prod_accum_116__13_, prod_accum_116__12_, prod_accum_116__11_, prod_accum_116__10_, prod_accum_116__9_, prod_accum_116__8_, prod_accum_116__7_, prod_accum_116__6_, prod_accum_116__5_, prod_accum_116__4_, prod_accum_116__3_, prod_accum_116__2_, prod_accum_116__1_, prod_accum_116__0_ })
  );


  bsg_mul_array_row_128_117_x
  genblk1_117__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[14975:14848]),
    .b_i(b_r[14975:14848]),
    .s_i({ s_r_116__127_, s_r_116__126_, s_r_116__125_, s_r_116__124_, s_r_116__123_, s_r_116__122_, s_r_116__121_, s_r_116__120_, s_r_116__119_, s_r_116__118_, s_r_116__117_, s_r_116__116_, s_r_116__115_, s_r_116__114_, s_r_116__113_, s_r_116__112_, s_r_116__111_, s_r_116__110_, s_r_116__109_, s_r_116__108_, s_r_116__107_, s_r_116__106_, s_r_116__105_, s_r_116__104_, s_r_116__103_, s_r_116__102_, s_r_116__101_, s_r_116__100_, s_r_116__99_, s_r_116__98_, s_r_116__97_, s_r_116__96_, s_r_116__95_, s_r_116__94_, s_r_116__93_, s_r_116__92_, s_r_116__91_, s_r_116__90_, s_r_116__89_, s_r_116__88_, s_r_116__87_, s_r_116__86_, s_r_116__85_, s_r_116__84_, s_r_116__83_, s_r_116__82_, s_r_116__81_, s_r_116__80_, s_r_116__79_, s_r_116__78_, s_r_116__77_, s_r_116__76_, s_r_116__75_, s_r_116__74_, s_r_116__73_, s_r_116__72_, s_r_116__71_, s_r_116__70_, s_r_116__69_, s_r_116__68_, s_r_116__67_, s_r_116__66_, s_r_116__65_, s_r_116__64_, s_r_116__63_, s_r_116__62_, s_r_116__61_, s_r_116__60_, s_r_116__59_, s_r_116__58_, s_r_116__57_, s_r_116__56_, s_r_116__55_, s_r_116__54_, s_r_116__53_, s_r_116__52_, s_r_116__51_, s_r_116__50_, s_r_116__49_, s_r_116__48_, s_r_116__47_, s_r_116__46_, s_r_116__45_, s_r_116__44_, s_r_116__43_, s_r_116__42_, s_r_116__41_, s_r_116__40_, s_r_116__39_, s_r_116__38_, s_r_116__37_, s_r_116__36_, s_r_116__35_, s_r_116__34_, s_r_116__33_, s_r_116__32_, s_r_116__31_, s_r_116__30_, s_r_116__29_, s_r_116__28_, s_r_116__27_, s_r_116__26_, s_r_116__25_, s_r_116__24_, s_r_116__23_, s_r_116__22_, s_r_116__21_, s_r_116__20_, s_r_116__19_, s_r_116__18_, s_r_116__17_, s_r_116__16_, s_r_116__15_, s_r_116__14_, s_r_116__13_, s_r_116__12_, s_r_116__11_, s_r_116__10_, s_r_116__9_, s_r_116__8_, s_r_116__7_, s_r_116__6_, s_r_116__5_, s_r_116__4_, s_r_116__3_, s_r_116__2_, s_r_116__1_, s_r_116__0_ }),
    .c_i(c_r[116]),
    .prod_accum_i({ prod_accum_116__117_, prod_accum_116__116_, prod_accum_116__115_, prod_accum_116__114_, prod_accum_116__113_, prod_accum_116__112_, prod_accum_116__111_, prod_accum_116__110_, prod_accum_116__109_, prod_accum_116__108_, prod_accum_116__107_, prod_accum_116__106_, prod_accum_116__105_, prod_accum_116__104_, prod_accum_116__103_, prod_accum_116__102_, prod_accum_116__101_, prod_accum_116__100_, prod_accum_116__99_, prod_accum_116__98_, prod_accum_116__97_, prod_accum_116__96_, prod_accum_116__95_, prod_accum_116__94_, prod_accum_116__93_, prod_accum_116__92_, prod_accum_116__91_, prod_accum_116__90_, prod_accum_116__89_, prod_accum_116__88_, prod_accum_116__87_, prod_accum_116__86_, prod_accum_116__85_, prod_accum_116__84_, prod_accum_116__83_, prod_accum_116__82_, prod_accum_116__81_, prod_accum_116__80_, prod_accum_116__79_, prod_accum_116__78_, prod_accum_116__77_, prod_accum_116__76_, prod_accum_116__75_, prod_accum_116__74_, prod_accum_116__73_, prod_accum_116__72_, prod_accum_116__71_, prod_accum_116__70_, prod_accum_116__69_, prod_accum_116__68_, prod_accum_116__67_, prod_accum_116__66_, prod_accum_116__65_, prod_accum_116__64_, prod_accum_116__63_, prod_accum_116__62_, prod_accum_116__61_, prod_accum_116__60_, prod_accum_116__59_, prod_accum_116__58_, prod_accum_116__57_, prod_accum_116__56_, prod_accum_116__55_, prod_accum_116__54_, prod_accum_116__53_, prod_accum_116__52_, prod_accum_116__51_, prod_accum_116__50_, prod_accum_116__49_, prod_accum_116__48_, prod_accum_116__47_, prod_accum_116__46_, prod_accum_116__45_, prod_accum_116__44_, prod_accum_116__43_, prod_accum_116__42_, prod_accum_116__41_, prod_accum_116__40_, prod_accum_116__39_, prod_accum_116__38_, prod_accum_116__37_, prod_accum_116__36_, prod_accum_116__35_, prod_accum_116__34_, prod_accum_116__33_, prod_accum_116__32_, prod_accum_116__31_, prod_accum_116__30_, prod_accum_116__29_, prod_accum_116__28_, prod_accum_116__27_, prod_accum_116__26_, prod_accum_116__25_, prod_accum_116__24_, prod_accum_116__23_, prod_accum_116__22_, prod_accum_116__21_, prod_accum_116__20_, prod_accum_116__19_, prod_accum_116__18_, prod_accum_116__17_, prod_accum_116__16_, prod_accum_116__15_, prod_accum_116__14_, prod_accum_116__13_, prod_accum_116__12_, prod_accum_116__11_, prod_accum_116__10_, prod_accum_116__9_, prod_accum_116__8_, prod_accum_116__7_, prod_accum_116__6_, prod_accum_116__5_, prod_accum_116__4_, prod_accum_116__3_, prod_accum_116__2_, prod_accum_116__1_, prod_accum_116__0_ }),
    .a_o(a_r[15103:14976]),
    .b_o(b_r[15103:14976]),
    .s_o({ s_r_117__127_, s_r_117__126_, s_r_117__125_, s_r_117__124_, s_r_117__123_, s_r_117__122_, s_r_117__121_, s_r_117__120_, s_r_117__119_, s_r_117__118_, s_r_117__117_, s_r_117__116_, s_r_117__115_, s_r_117__114_, s_r_117__113_, s_r_117__112_, s_r_117__111_, s_r_117__110_, s_r_117__109_, s_r_117__108_, s_r_117__107_, s_r_117__106_, s_r_117__105_, s_r_117__104_, s_r_117__103_, s_r_117__102_, s_r_117__101_, s_r_117__100_, s_r_117__99_, s_r_117__98_, s_r_117__97_, s_r_117__96_, s_r_117__95_, s_r_117__94_, s_r_117__93_, s_r_117__92_, s_r_117__91_, s_r_117__90_, s_r_117__89_, s_r_117__88_, s_r_117__87_, s_r_117__86_, s_r_117__85_, s_r_117__84_, s_r_117__83_, s_r_117__82_, s_r_117__81_, s_r_117__80_, s_r_117__79_, s_r_117__78_, s_r_117__77_, s_r_117__76_, s_r_117__75_, s_r_117__74_, s_r_117__73_, s_r_117__72_, s_r_117__71_, s_r_117__70_, s_r_117__69_, s_r_117__68_, s_r_117__67_, s_r_117__66_, s_r_117__65_, s_r_117__64_, s_r_117__63_, s_r_117__62_, s_r_117__61_, s_r_117__60_, s_r_117__59_, s_r_117__58_, s_r_117__57_, s_r_117__56_, s_r_117__55_, s_r_117__54_, s_r_117__53_, s_r_117__52_, s_r_117__51_, s_r_117__50_, s_r_117__49_, s_r_117__48_, s_r_117__47_, s_r_117__46_, s_r_117__45_, s_r_117__44_, s_r_117__43_, s_r_117__42_, s_r_117__41_, s_r_117__40_, s_r_117__39_, s_r_117__38_, s_r_117__37_, s_r_117__36_, s_r_117__35_, s_r_117__34_, s_r_117__33_, s_r_117__32_, s_r_117__31_, s_r_117__30_, s_r_117__29_, s_r_117__28_, s_r_117__27_, s_r_117__26_, s_r_117__25_, s_r_117__24_, s_r_117__23_, s_r_117__22_, s_r_117__21_, s_r_117__20_, s_r_117__19_, s_r_117__18_, s_r_117__17_, s_r_117__16_, s_r_117__15_, s_r_117__14_, s_r_117__13_, s_r_117__12_, s_r_117__11_, s_r_117__10_, s_r_117__9_, s_r_117__8_, s_r_117__7_, s_r_117__6_, s_r_117__5_, s_r_117__4_, s_r_117__3_, s_r_117__2_, s_r_117__1_, s_r_117__0_ }),
    .c_o(c_r[117]),
    .prod_accum_o({ prod_accum_117__118_, prod_accum_117__117_, prod_accum_117__116_, prod_accum_117__115_, prod_accum_117__114_, prod_accum_117__113_, prod_accum_117__112_, prod_accum_117__111_, prod_accum_117__110_, prod_accum_117__109_, prod_accum_117__108_, prod_accum_117__107_, prod_accum_117__106_, prod_accum_117__105_, prod_accum_117__104_, prod_accum_117__103_, prod_accum_117__102_, prod_accum_117__101_, prod_accum_117__100_, prod_accum_117__99_, prod_accum_117__98_, prod_accum_117__97_, prod_accum_117__96_, prod_accum_117__95_, prod_accum_117__94_, prod_accum_117__93_, prod_accum_117__92_, prod_accum_117__91_, prod_accum_117__90_, prod_accum_117__89_, prod_accum_117__88_, prod_accum_117__87_, prod_accum_117__86_, prod_accum_117__85_, prod_accum_117__84_, prod_accum_117__83_, prod_accum_117__82_, prod_accum_117__81_, prod_accum_117__80_, prod_accum_117__79_, prod_accum_117__78_, prod_accum_117__77_, prod_accum_117__76_, prod_accum_117__75_, prod_accum_117__74_, prod_accum_117__73_, prod_accum_117__72_, prod_accum_117__71_, prod_accum_117__70_, prod_accum_117__69_, prod_accum_117__68_, prod_accum_117__67_, prod_accum_117__66_, prod_accum_117__65_, prod_accum_117__64_, prod_accum_117__63_, prod_accum_117__62_, prod_accum_117__61_, prod_accum_117__60_, prod_accum_117__59_, prod_accum_117__58_, prod_accum_117__57_, prod_accum_117__56_, prod_accum_117__55_, prod_accum_117__54_, prod_accum_117__53_, prod_accum_117__52_, prod_accum_117__51_, prod_accum_117__50_, prod_accum_117__49_, prod_accum_117__48_, prod_accum_117__47_, prod_accum_117__46_, prod_accum_117__45_, prod_accum_117__44_, prod_accum_117__43_, prod_accum_117__42_, prod_accum_117__41_, prod_accum_117__40_, prod_accum_117__39_, prod_accum_117__38_, prod_accum_117__37_, prod_accum_117__36_, prod_accum_117__35_, prod_accum_117__34_, prod_accum_117__33_, prod_accum_117__32_, prod_accum_117__31_, prod_accum_117__30_, prod_accum_117__29_, prod_accum_117__28_, prod_accum_117__27_, prod_accum_117__26_, prod_accum_117__25_, prod_accum_117__24_, prod_accum_117__23_, prod_accum_117__22_, prod_accum_117__21_, prod_accum_117__20_, prod_accum_117__19_, prod_accum_117__18_, prod_accum_117__17_, prod_accum_117__16_, prod_accum_117__15_, prod_accum_117__14_, prod_accum_117__13_, prod_accum_117__12_, prod_accum_117__11_, prod_accum_117__10_, prod_accum_117__9_, prod_accum_117__8_, prod_accum_117__7_, prod_accum_117__6_, prod_accum_117__5_, prod_accum_117__4_, prod_accum_117__3_, prod_accum_117__2_, prod_accum_117__1_, prod_accum_117__0_ })
  );


  bsg_mul_array_row_128_118_x
  genblk1_118__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[15103:14976]),
    .b_i(b_r[15103:14976]),
    .s_i({ s_r_117__127_, s_r_117__126_, s_r_117__125_, s_r_117__124_, s_r_117__123_, s_r_117__122_, s_r_117__121_, s_r_117__120_, s_r_117__119_, s_r_117__118_, s_r_117__117_, s_r_117__116_, s_r_117__115_, s_r_117__114_, s_r_117__113_, s_r_117__112_, s_r_117__111_, s_r_117__110_, s_r_117__109_, s_r_117__108_, s_r_117__107_, s_r_117__106_, s_r_117__105_, s_r_117__104_, s_r_117__103_, s_r_117__102_, s_r_117__101_, s_r_117__100_, s_r_117__99_, s_r_117__98_, s_r_117__97_, s_r_117__96_, s_r_117__95_, s_r_117__94_, s_r_117__93_, s_r_117__92_, s_r_117__91_, s_r_117__90_, s_r_117__89_, s_r_117__88_, s_r_117__87_, s_r_117__86_, s_r_117__85_, s_r_117__84_, s_r_117__83_, s_r_117__82_, s_r_117__81_, s_r_117__80_, s_r_117__79_, s_r_117__78_, s_r_117__77_, s_r_117__76_, s_r_117__75_, s_r_117__74_, s_r_117__73_, s_r_117__72_, s_r_117__71_, s_r_117__70_, s_r_117__69_, s_r_117__68_, s_r_117__67_, s_r_117__66_, s_r_117__65_, s_r_117__64_, s_r_117__63_, s_r_117__62_, s_r_117__61_, s_r_117__60_, s_r_117__59_, s_r_117__58_, s_r_117__57_, s_r_117__56_, s_r_117__55_, s_r_117__54_, s_r_117__53_, s_r_117__52_, s_r_117__51_, s_r_117__50_, s_r_117__49_, s_r_117__48_, s_r_117__47_, s_r_117__46_, s_r_117__45_, s_r_117__44_, s_r_117__43_, s_r_117__42_, s_r_117__41_, s_r_117__40_, s_r_117__39_, s_r_117__38_, s_r_117__37_, s_r_117__36_, s_r_117__35_, s_r_117__34_, s_r_117__33_, s_r_117__32_, s_r_117__31_, s_r_117__30_, s_r_117__29_, s_r_117__28_, s_r_117__27_, s_r_117__26_, s_r_117__25_, s_r_117__24_, s_r_117__23_, s_r_117__22_, s_r_117__21_, s_r_117__20_, s_r_117__19_, s_r_117__18_, s_r_117__17_, s_r_117__16_, s_r_117__15_, s_r_117__14_, s_r_117__13_, s_r_117__12_, s_r_117__11_, s_r_117__10_, s_r_117__9_, s_r_117__8_, s_r_117__7_, s_r_117__6_, s_r_117__5_, s_r_117__4_, s_r_117__3_, s_r_117__2_, s_r_117__1_, s_r_117__0_ }),
    .c_i(c_r[117]),
    .prod_accum_i({ prod_accum_117__118_, prod_accum_117__117_, prod_accum_117__116_, prod_accum_117__115_, prod_accum_117__114_, prod_accum_117__113_, prod_accum_117__112_, prod_accum_117__111_, prod_accum_117__110_, prod_accum_117__109_, prod_accum_117__108_, prod_accum_117__107_, prod_accum_117__106_, prod_accum_117__105_, prod_accum_117__104_, prod_accum_117__103_, prod_accum_117__102_, prod_accum_117__101_, prod_accum_117__100_, prod_accum_117__99_, prod_accum_117__98_, prod_accum_117__97_, prod_accum_117__96_, prod_accum_117__95_, prod_accum_117__94_, prod_accum_117__93_, prod_accum_117__92_, prod_accum_117__91_, prod_accum_117__90_, prod_accum_117__89_, prod_accum_117__88_, prod_accum_117__87_, prod_accum_117__86_, prod_accum_117__85_, prod_accum_117__84_, prod_accum_117__83_, prod_accum_117__82_, prod_accum_117__81_, prod_accum_117__80_, prod_accum_117__79_, prod_accum_117__78_, prod_accum_117__77_, prod_accum_117__76_, prod_accum_117__75_, prod_accum_117__74_, prod_accum_117__73_, prod_accum_117__72_, prod_accum_117__71_, prod_accum_117__70_, prod_accum_117__69_, prod_accum_117__68_, prod_accum_117__67_, prod_accum_117__66_, prod_accum_117__65_, prod_accum_117__64_, prod_accum_117__63_, prod_accum_117__62_, prod_accum_117__61_, prod_accum_117__60_, prod_accum_117__59_, prod_accum_117__58_, prod_accum_117__57_, prod_accum_117__56_, prod_accum_117__55_, prod_accum_117__54_, prod_accum_117__53_, prod_accum_117__52_, prod_accum_117__51_, prod_accum_117__50_, prod_accum_117__49_, prod_accum_117__48_, prod_accum_117__47_, prod_accum_117__46_, prod_accum_117__45_, prod_accum_117__44_, prod_accum_117__43_, prod_accum_117__42_, prod_accum_117__41_, prod_accum_117__40_, prod_accum_117__39_, prod_accum_117__38_, prod_accum_117__37_, prod_accum_117__36_, prod_accum_117__35_, prod_accum_117__34_, prod_accum_117__33_, prod_accum_117__32_, prod_accum_117__31_, prod_accum_117__30_, prod_accum_117__29_, prod_accum_117__28_, prod_accum_117__27_, prod_accum_117__26_, prod_accum_117__25_, prod_accum_117__24_, prod_accum_117__23_, prod_accum_117__22_, prod_accum_117__21_, prod_accum_117__20_, prod_accum_117__19_, prod_accum_117__18_, prod_accum_117__17_, prod_accum_117__16_, prod_accum_117__15_, prod_accum_117__14_, prod_accum_117__13_, prod_accum_117__12_, prod_accum_117__11_, prod_accum_117__10_, prod_accum_117__9_, prod_accum_117__8_, prod_accum_117__7_, prod_accum_117__6_, prod_accum_117__5_, prod_accum_117__4_, prod_accum_117__3_, prod_accum_117__2_, prod_accum_117__1_, prod_accum_117__0_ }),
    .a_o(a_r[15231:15104]),
    .b_o(b_r[15231:15104]),
    .s_o({ s_r_118__127_, s_r_118__126_, s_r_118__125_, s_r_118__124_, s_r_118__123_, s_r_118__122_, s_r_118__121_, s_r_118__120_, s_r_118__119_, s_r_118__118_, s_r_118__117_, s_r_118__116_, s_r_118__115_, s_r_118__114_, s_r_118__113_, s_r_118__112_, s_r_118__111_, s_r_118__110_, s_r_118__109_, s_r_118__108_, s_r_118__107_, s_r_118__106_, s_r_118__105_, s_r_118__104_, s_r_118__103_, s_r_118__102_, s_r_118__101_, s_r_118__100_, s_r_118__99_, s_r_118__98_, s_r_118__97_, s_r_118__96_, s_r_118__95_, s_r_118__94_, s_r_118__93_, s_r_118__92_, s_r_118__91_, s_r_118__90_, s_r_118__89_, s_r_118__88_, s_r_118__87_, s_r_118__86_, s_r_118__85_, s_r_118__84_, s_r_118__83_, s_r_118__82_, s_r_118__81_, s_r_118__80_, s_r_118__79_, s_r_118__78_, s_r_118__77_, s_r_118__76_, s_r_118__75_, s_r_118__74_, s_r_118__73_, s_r_118__72_, s_r_118__71_, s_r_118__70_, s_r_118__69_, s_r_118__68_, s_r_118__67_, s_r_118__66_, s_r_118__65_, s_r_118__64_, s_r_118__63_, s_r_118__62_, s_r_118__61_, s_r_118__60_, s_r_118__59_, s_r_118__58_, s_r_118__57_, s_r_118__56_, s_r_118__55_, s_r_118__54_, s_r_118__53_, s_r_118__52_, s_r_118__51_, s_r_118__50_, s_r_118__49_, s_r_118__48_, s_r_118__47_, s_r_118__46_, s_r_118__45_, s_r_118__44_, s_r_118__43_, s_r_118__42_, s_r_118__41_, s_r_118__40_, s_r_118__39_, s_r_118__38_, s_r_118__37_, s_r_118__36_, s_r_118__35_, s_r_118__34_, s_r_118__33_, s_r_118__32_, s_r_118__31_, s_r_118__30_, s_r_118__29_, s_r_118__28_, s_r_118__27_, s_r_118__26_, s_r_118__25_, s_r_118__24_, s_r_118__23_, s_r_118__22_, s_r_118__21_, s_r_118__20_, s_r_118__19_, s_r_118__18_, s_r_118__17_, s_r_118__16_, s_r_118__15_, s_r_118__14_, s_r_118__13_, s_r_118__12_, s_r_118__11_, s_r_118__10_, s_r_118__9_, s_r_118__8_, s_r_118__7_, s_r_118__6_, s_r_118__5_, s_r_118__4_, s_r_118__3_, s_r_118__2_, s_r_118__1_, s_r_118__0_ }),
    .c_o(c_r[118]),
    .prod_accum_o({ prod_accum_118__119_, prod_accum_118__118_, prod_accum_118__117_, prod_accum_118__116_, prod_accum_118__115_, prod_accum_118__114_, prod_accum_118__113_, prod_accum_118__112_, prod_accum_118__111_, prod_accum_118__110_, prod_accum_118__109_, prod_accum_118__108_, prod_accum_118__107_, prod_accum_118__106_, prod_accum_118__105_, prod_accum_118__104_, prod_accum_118__103_, prod_accum_118__102_, prod_accum_118__101_, prod_accum_118__100_, prod_accum_118__99_, prod_accum_118__98_, prod_accum_118__97_, prod_accum_118__96_, prod_accum_118__95_, prod_accum_118__94_, prod_accum_118__93_, prod_accum_118__92_, prod_accum_118__91_, prod_accum_118__90_, prod_accum_118__89_, prod_accum_118__88_, prod_accum_118__87_, prod_accum_118__86_, prod_accum_118__85_, prod_accum_118__84_, prod_accum_118__83_, prod_accum_118__82_, prod_accum_118__81_, prod_accum_118__80_, prod_accum_118__79_, prod_accum_118__78_, prod_accum_118__77_, prod_accum_118__76_, prod_accum_118__75_, prod_accum_118__74_, prod_accum_118__73_, prod_accum_118__72_, prod_accum_118__71_, prod_accum_118__70_, prod_accum_118__69_, prod_accum_118__68_, prod_accum_118__67_, prod_accum_118__66_, prod_accum_118__65_, prod_accum_118__64_, prod_accum_118__63_, prod_accum_118__62_, prod_accum_118__61_, prod_accum_118__60_, prod_accum_118__59_, prod_accum_118__58_, prod_accum_118__57_, prod_accum_118__56_, prod_accum_118__55_, prod_accum_118__54_, prod_accum_118__53_, prod_accum_118__52_, prod_accum_118__51_, prod_accum_118__50_, prod_accum_118__49_, prod_accum_118__48_, prod_accum_118__47_, prod_accum_118__46_, prod_accum_118__45_, prod_accum_118__44_, prod_accum_118__43_, prod_accum_118__42_, prod_accum_118__41_, prod_accum_118__40_, prod_accum_118__39_, prod_accum_118__38_, prod_accum_118__37_, prod_accum_118__36_, prod_accum_118__35_, prod_accum_118__34_, prod_accum_118__33_, prod_accum_118__32_, prod_accum_118__31_, prod_accum_118__30_, prod_accum_118__29_, prod_accum_118__28_, prod_accum_118__27_, prod_accum_118__26_, prod_accum_118__25_, prod_accum_118__24_, prod_accum_118__23_, prod_accum_118__22_, prod_accum_118__21_, prod_accum_118__20_, prod_accum_118__19_, prod_accum_118__18_, prod_accum_118__17_, prod_accum_118__16_, prod_accum_118__15_, prod_accum_118__14_, prod_accum_118__13_, prod_accum_118__12_, prod_accum_118__11_, prod_accum_118__10_, prod_accum_118__9_, prod_accum_118__8_, prod_accum_118__7_, prod_accum_118__6_, prod_accum_118__5_, prod_accum_118__4_, prod_accum_118__3_, prod_accum_118__2_, prod_accum_118__1_, prod_accum_118__0_ })
  );


  bsg_mul_array_row_128_119_x
  genblk1_119__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[15231:15104]),
    .b_i(b_r[15231:15104]),
    .s_i({ s_r_118__127_, s_r_118__126_, s_r_118__125_, s_r_118__124_, s_r_118__123_, s_r_118__122_, s_r_118__121_, s_r_118__120_, s_r_118__119_, s_r_118__118_, s_r_118__117_, s_r_118__116_, s_r_118__115_, s_r_118__114_, s_r_118__113_, s_r_118__112_, s_r_118__111_, s_r_118__110_, s_r_118__109_, s_r_118__108_, s_r_118__107_, s_r_118__106_, s_r_118__105_, s_r_118__104_, s_r_118__103_, s_r_118__102_, s_r_118__101_, s_r_118__100_, s_r_118__99_, s_r_118__98_, s_r_118__97_, s_r_118__96_, s_r_118__95_, s_r_118__94_, s_r_118__93_, s_r_118__92_, s_r_118__91_, s_r_118__90_, s_r_118__89_, s_r_118__88_, s_r_118__87_, s_r_118__86_, s_r_118__85_, s_r_118__84_, s_r_118__83_, s_r_118__82_, s_r_118__81_, s_r_118__80_, s_r_118__79_, s_r_118__78_, s_r_118__77_, s_r_118__76_, s_r_118__75_, s_r_118__74_, s_r_118__73_, s_r_118__72_, s_r_118__71_, s_r_118__70_, s_r_118__69_, s_r_118__68_, s_r_118__67_, s_r_118__66_, s_r_118__65_, s_r_118__64_, s_r_118__63_, s_r_118__62_, s_r_118__61_, s_r_118__60_, s_r_118__59_, s_r_118__58_, s_r_118__57_, s_r_118__56_, s_r_118__55_, s_r_118__54_, s_r_118__53_, s_r_118__52_, s_r_118__51_, s_r_118__50_, s_r_118__49_, s_r_118__48_, s_r_118__47_, s_r_118__46_, s_r_118__45_, s_r_118__44_, s_r_118__43_, s_r_118__42_, s_r_118__41_, s_r_118__40_, s_r_118__39_, s_r_118__38_, s_r_118__37_, s_r_118__36_, s_r_118__35_, s_r_118__34_, s_r_118__33_, s_r_118__32_, s_r_118__31_, s_r_118__30_, s_r_118__29_, s_r_118__28_, s_r_118__27_, s_r_118__26_, s_r_118__25_, s_r_118__24_, s_r_118__23_, s_r_118__22_, s_r_118__21_, s_r_118__20_, s_r_118__19_, s_r_118__18_, s_r_118__17_, s_r_118__16_, s_r_118__15_, s_r_118__14_, s_r_118__13_, s_r_118__12_, s_r_118__11_, s_r_118__10_, s_r_118__9_, s_r_118__8_, s_r_118__7_, s_r_118__6_, s_r_118__5_, s_r_118__4_, s_r_118__3_, s_r_118__2_, s_r_118__1_, s_r_118__0_ }),
    .c_i(c_r[118]),
    .prod_accum_i({ prod_accum_118__119_, prod_accum_118__118_, prod_accum_118__117_, prod_accum_118__116_, prod_accum_118__115_, prod_accum_118__114_, prod_accum_118__113_, prod_accum_118__112_, prod_accum_118__111_, prod_accum_118__110_, prod_accum_118__109_, prod_accum_118__108_, prod_accum_118__107_, prod_accum_118__106_, prod_accum_118__105_, prod_accum_118__104_, prod_accum_118__103_, prod_accum_118__102_, prod_accum_118__101_, prod_accum_118__100_, prod_accum_118__99_, prod_accum_118__98_, prod_accum_118__97_, prod_accum_118__96_, prod_accum_118__95_, prod_accum_118__94_, prod_accum_118__93_, prod_accum_118__92_, prod_accum_118__91_, prod_accum_118__90_, prod_accum_118__89_, prod_accum_118__88_, prod_accum_118__87_, prod_accum_118__86_, prod_accum_118__85_, prod_accum_118__84_, prod_accum_118__83_, prod_accum_118__82_, prod_accum_118__81_, prod_accum_118__80_, prod_accum_118__79_, prod_accum_118__78_, prod_accum_118__77_, prod_accum_118__76_, prod_accum_118__75_, prod_accum_118__74_, prod_accum_118__73_, prod_accum_118__72_, prod_accum_118__71_, prod_accum_118__70_, prod_accum_118__69_, prod_accum_118__68_, prod_accum_118__67_, prod_accum_118__66_, prod_accum_118__65_, prod_accum_118__64_, prod_accum_118__63_, prod_accum_118__62_, prod_accum_118__61_, prod_accum_118__60_, prod_accum_118__59_, prod_accum_118__58_, prod_accum_118__57_, prod_accum_118__56_, prod_accum_118__55_, prod_accum_118__54_, prod_accum_118__53_, prod_accum_118__52_, prod_accum_118__51_, prod_accum_118__50_, prod_accum_118__49_, prod_accum_118__48_, prod_accum_118__47_, prod_accum_118__46_, prod_accum_118__45_, prod_accum_118__44_, prod_accum_118__43_, prod_accum_118__42_, prod_accum_118__41_, prod_accum_118__40_, prod_accum_118__39_, prod_accum_118__38_, prod_accum_118__37_, prod_accum_118__36_, prod_accum_118__35_, prod_accum_118__34_, prod_accum_118__33_, prod_accum_118__32_, prod_accum_118__31_, prod_accum_118__30_, prod_accum_118__29_, prod_accum_118__28_, prod_accum_118__27_, prod_accum_118__26_, prod_accum_118__25_, prod_accum_118__24_, prod_accum_118__23_, prod_accum_118__22_, prod_accum_118__21_, prod_accum_118__20_, prod_accum_118__19_, prod_accum_118__18_, prod_accum_118__17_, prod_accum_118__16_, prod_accum_118__15_, prod_accum_118__14_, prod_accum_118__13_, prod_accum_118__12_, prod_accum_118__11_, prod_accum_118__10_, prod_accum_118__9_, prod_accum_118__8_, prod_accum_118__7_, prod_accum_118__6_, prod_accum_118__5_, prod_accum_118__4_, prod_accum_118__3_, prod_accum_118__2_, prod_accum_118__1_, prod_accum_118__0_ }),
    .a_o(a_r[15359:15232]),
    .b_o(b_r[15359:15232]),
    .s_o({ s_r_119__127_, s_r_119__126_, s_r_119__125_, s_r_119__124_, s_r_119__123_, s_r_119__122_, s_r_119__121_, s_r_119__120_, s_r_119__119_, s_r_119__118_, s_r_119__117_, s_r_119__116_, s_r_119__115_, s_r_119__114_, s_r_119__113_, s_r_119__112_, s_r_119__111_, s_r_119__110_, s_r_119__109_, s_r_119__108_, s_r_119__107_, s_r_119__106_, s_r_119__105_, s_r_119__104_, s_r_119__103_, s_r_119__102_, s_r_119__101_, s_r_119__100_, s_r_119__99_, s_r_119__98_, s_r_119__97_, s_r_119__96_, s_r_119__95_, s_r_119__94_, s_r_119__93_, s_r_119__92_, s_r_119__91_, s_r_119__90_, s_r_119__89_, s_r_119__88_, s_r_119__87_, s_r_119__86_, s_r_119__85_, s_r_119__84_, s_r_119__83_, s_r_119__82_, s_r_119__81_, s_r_119__80_, s_r_119__79_, s_r_119__78_, s_r_119__77_, s_r_119__76_, s_r_119__75_, s_r_119__74_, s_r_119__73_, s_r_119__72_, s_r_119__71_, s_r_119__70_, s_r_119__69_, s_r_119__68_, s_r_119__67_, s_r_119__66_, s_r_119__65_, s_r_119__64_, s_r_119__63_, s_r_119__62_, s_r_119__61_, s_r_119__60_, s_r_119__59_, s_r_119__58_, s_r_119__57_, s_r_119__56_, s_r_119__55_, s_r_119__54_, s_r_119__53_, s_r_119__52_, s_r_119__51_, s_r_119__50_, s_r_119__49_, s_r_119__48_, s_r_119__47_, s_r_119__46_, s_r_119__45_, s_r_119__44_, s_r_119__43_, s_r_119__42_, s_r_119__41_, s_r_119__40_, s_r_119__39_, s_r_119__38_, s_r_119__37_, s_r_119__36_, s_r_119__35_, s_r_119__34_, s_r_119__33_, s_r_119__32_, s_r_119__31_, s_r_119__30_, s_r_119__29_, s_r_119__28_, s_r_119__27_, s_r_119__26_, s_r_119__25_, s_r_119__24_, s_r_119__23_, s_r_119__22_, s_r_119__21_, s_r_119__20_, s_r_119__19_, s_r_119__18_, s_r_119__17_, s_r_119__16_, s_r_119__15_, s_r_119__14_, s_r_119__13_, s_r_119__12_, s_r_119__11_, s_r_119__10_, s_r_119__9_, s_r_119__8_, s_r_119__7_, s_r_119__6_, s_r_119__5_, s_r_119__4_, s_r_119__3_, s_r_119__2_, s_r_119__1_, s_r_119__0_ }),
    .c_o(c_r[119]),
    .prod_accum_o({ prod_accum_119__120_, prod_accum_119__119_, prod_accum_119__118_, prod_accum_119__117_, prod_accum_119__116_, prod_accum_119__115_, prod_accum_119__114_, prod_accum_119__113_, prod_accum_119__112_, prod_accum_119__111_, prod_accum_119__110_, prod_accum_119__109_, prod_accum_119__108_, prod_accum_119__107_, prod_accum_119__106_, prod_accum_119__105_, prod_accum_119__104_, prod_accum_119__103_, prod_accum_119__102_, prod_accum_119__101_, prod_accum_119__100_, prod_accum_119__99_, prod_accum_119__98_, prod_accum_119__97_, prod_accum_119__96_, prod_accum_119__95_, prod_accum_119__94_, prod_accum_119__93_, prod_accum_119__92_, prod_accum_119__91_, prod_accum_119__90_, prod_accum_119__89_, prod_accum_119__88_, prod_accum_119__87_, prod_accum_119__86_, prod_accum_119__85_, prod_accum_119__84_, prod_accum_119__83_, prod_accum_119__82_, prod_accum_119__81_, prod_accum_119__80_, prod_accum_119__79_, prod_accum_119__78_, prod_accum_119__77_, prod_accum_119__76_, prod_accum_119__75_, prod_accum_119__74_, prod_accum_119__73_, prod_accum_119__72_, prod_accum_119__71_, prod_accum_119__70_, prod_accum_119__69_, prod_accum_119__68_, prod_accum_119__67_, prod_accum_119__66_, prod_accum_119__65_, prod_accum_119__64_, prod_accum_119__63_, prod_accum_119__62_, prod_accum_119__61_, prod_accum_119__60_, prod_accum_119__59_, prod_accum_119__58_, prod_accum_119__57_, prod_accum_119__56_, prod_accum_119__55_, prod_accum_119__54_, prod_accum_119__53_, prod_accum_119__52_, prod_accum_119__51_, prod_accum_119__50_, prod_accum_119__49_, prod_accum_119__48_, prod_accum_119__47_, prod_accum_119__46_, prod_accum_119__45_, prod_accum_119__44_, prod_accum_119__43_, prod_accum_119__42_, prod_accum_119__41_, prod_accum_119__40_, prod_accum_119__39_, prod_accum_119__38_, prod_accum_119__37_, prod_accum_119__36_, prod_accum_119__35_, prod_accum_119__34_, prod_accum_119__33_, prod_accum_119__32_, prod_accum_119__31_, prod_accum_119__30_, prod_accum_119__29_, prod_accum_119__28_, prod_accum_119__27_, prod_accum_119__26_, prod_accum_119__25_, prod_accum_119__24_, prod_accum_119__23_, prod_accum_119__22_, prod_accum_119__21_, prod_accum_119__20_, prod_accum_119__19_, prod_accum_119__18_, prod_accum_119__17_, prod_accum_119__16_, prod_accum_119__15_, prod_accum_119__14_, prod_accum_119__13_, prod_accum_119__12_, prod_accum_119__11_, prod_accum_119__10_, prod_accum_119__9_, prod_accum_119__8_, prod_accum_119__7_, prod_accum_119__6_, prod_accum_119__5_, prod_accum_119__4_, prod_accum_119__3_, prod_accum_119__2_, prod_accum_119__1_, prod_accum_119__0_ })
  );


  bsg_mul_array_row_128_120_x
  genblk1_120__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[15359:15232]),
    .b_i(b_r[15359:15232]),
    .s_i({ s_r_119__127_, s_r_119__126_, s_r_119__125_, s_r_119__124_, s_r_119__123_, s_r_119__122_, s_r_119__121_, s_r_119__120_, s_r_119__119_, s_r_119__118_, s_r_119__117_, s_r_119__116_, s_r_119__115_, s_r_119__114_, s_r_119__113_, s_r_119__112_, s_r_119__111_, s_r_119__110_, s_r_119__109_, s_r_119__108_, s_r_119__107_, s_r_119__106_, s_r_119__105_, s_r_119__104_, s_r_119__103_, s_r_119__102_, s_r_119__101_, s_r_119__100_, s_r_119__99_, s_r_119__98_, s_r_119__97_, s_r_119__96_, s_r_119__95_, s_r_119__94_, s_r_119__93_, s_r_119__92_, s_r_119__91_, s_r_119__90_, s_r_119__89_, s_r_119__88_, s_r_119__87_, s_r_119__86_, s_r_119__85_, s_r_119__84_, s_r_119__83_, s_r_119__82_, s_r_119__81_, s_r_119__80_, s_r_119__79_, s_r_119__78_, s_r_119__77_, s_r_119__76_, s_r_119__75_, s_r_119__74_, s_r_119__73_, s_r_119__72_, s_r_119__71_, s_r_119__70_, s_r_119__69_, s_r_119__68_, s_r_119__67_, s_r_119__66_, s_r_119__65_, s_r_119__64_, s_r_119__63_, s_r_119__62_, s_r_119__61_, s_r_119__60_, s_r_119__59_, s_r_119__58_, s_r_119__57_, s_r_119__56_, s_r_119__55_, s_r_119__54_, s_r_119__53_, s_r_119__52_, s_r_119__51_, s_r_119__50_, s_r_119__49_, s_r_119__48_, s_r_119__47_, s_r_119__46_, s_r_119__45_, s_r_119__44_, s_r_119__43_, s_r_119__42_, s_r_119__41_, s_r_119__40_, s_r_119__39_, s_r_119__38_, s_r_119__37_, s_r_119__36_, s_r_119__35_, s_r_119__34_, s_r_119__33_, s_r_119__32_, s_r_119__31_, s_r_119__30_, s_r_119__29_, s_r_119__28_, s_r_119__27_, s_r_119__26_, s_r_119__25_, s_r_119__24_, s_r_119__23_, s_r_119__22_, s_r_119__21_, s_r_119__20_, s_r_119__19_, s_r_119__18_, s_r_119__17_, s_r_119__16_, s_r_119__15_, s_r_119__14_, s_r_119__13_, s_r_119__12_, s_r_119__11_, s_r_119__10_, s_r_119__9_, s_r_119__8_, s_r_119__7_, s_r_119__6_, s_r_119__5_, s_r_119__4_, s_r_119__3_, s_r_119__2_, s_r_119__1_, s_r_119__0_ }),
    .c_i(c_r[119]),
    .prod_accum_i({ prod_accum_119__120_, prod_accum_119__119_, prod_accum_119__118_, prod_accum_119__117_, prod_accum_119__116_, prod_accum_119__115_, prod_accum_119__114_, prod_accum_119__113_, prod_accum_119__112_, prod_accum_119__111_, prod_accum_119__110_, prod_accum_119__109_, prod_accum_119__108_, prod_accum_119__107_, prod_accum_119__106_, prod_accum_119__105_, prod_accum_119__104_, prod_accum_119__103_, prod_accum_119__102_, prod_accum_119__101_, prod_accum_119__100_, prod_accum_119__99_, prod_accum_119__98_, prod_accum_119__97_, prod_accum_119__96_, prod_accum_119__95_, prod_accum_119__94_, prod_accum_119__93_, prod_accum_119__92_, prod_accum_119__91_, prod_accum_119__90_, prod_accum_119__89_, prod_accum_119__88_, prod_accum_119__87_, prod_accum_119__86_, prod_accum_119__85_, prod_accum_119__84_, prod_accum_119__83_, prod_accum_119__82_, prod_accum_119__81_, prod_accum_119__80_, prod_accum_119__79_, prod_accum_119__78_, prod_accum_119__77_, prod_accum_119__76_, prod_accum_119__75_, prod_accum_119__74_, prod_accum_119__73_, prod_accum_119__72_, prod_accum_119__71_, prod_accum_119__70_, prod_accum_119__69_, prod_accum_119__68_, prod_accum_119__67_, prod_accum_119__66_, prod_accum_119__65_, prod_accum_119__64_, prod_accum_119__63_, prod_accum_119__62_, prod_accum_119__61_, prod_accum_119__60_, prod_accum_119__59_, prod_accum_119__58_, prod_accum_119__57_, prod_accum_119__56_, prod_accum_119__55_, prod_accum_119__54_, prod_accum_119__53_, prod_accum_119__52_, prod_accum_119__51_, prod_accum_119__50_, prod_accum_119__49_, prod_accum_119__48_, prod_accum_119__47_, prod_accum_119__46_, prod_accum_119__45_, prod_accum_119__44_, prod_accum_119__43_, prod_accum_119__42_, prod_accum_119__41_, prod_accum_119__40_, prod_accum_119__39_, prod_accum_119__38_, prod_accum_119__37_, prod_accum_119__36_, prod_accum_119__35_, prod_accum_119__34_, prod_accum_119__33_, prod_accum_119__32_, prod_accum_119__31_, prod_accum_119__30_, prod_accum_119__29_, prod_accum_119__28_, prod_accum_119__27_, prod_accum_119__26_, prod_accum_119__25_, prod_accum_119__24_, prod_accum_119__23_, prod_accum_119__22_, prod_accum_119__21_, prod_accum_119__20_, prod_accum_119__19_, prod_accum_119__18_, prod_accum_119__17_, prod_accum_119__16_, prod_accum_119__15_, prod_accum_119__14_, prod_accum_119__13_, prod_accum_119__12_, prod_accum_119__11_, prod_accum_119__10_, prod_accum_119__9_, prod_accum_119__8_, prod_accum_119__7_, prod_accum_119__6_, prod_accum_119__5_, prod_accum_119__4_, prod_accum_119__3_, prod_accum_119__2_, prod_accum_119__1_, prod_accum_119__0_ }),
    .a_o(a_r[15487:15360]),
    .b_o(b_r[15487:15360]),
    .s_o({ s_r_120__127_, s_r_120__126_, s_r_120__125_, s_r_120__124_, s_r_120__123_, s_r_120__122_, s_r_120__121_, s_r_120__120_, s_r_120__119_, s_r_120__118_, s_r_120__117_, s_r_120__116_, s_r_120__115_, s_r_120__114_, s_r_120__113_, s_r_120__112_, s_r_120__111_, s_r_120__110_, s_r_120__109_, s_r_120__108_, s_r_120__107_, s_r_120__106_, s_r_120__105_, s_r_120__104_, s_r_120__103_, s_r_120__102_, s_r_120__101_, s_r_120__100_, s_r_120__99_, s_r_120__98_, s_r_120__97_, s_r_120__96_, s_r_120__95_, s_r_120__94_, s_r_120__93_, s_r_120__92_, s_r_120__91_, s_r_120__90_, s_r_120__89_, s_r_120__88_, s_r_120__87_, s_r_120__86_, s_r_120__85_, s_r_120__84_, s_r_120__83_, s_r_120__82_, s_r_120__81_, s_r_120__80_, s_r_120__79_, s_r_120__78_, s_r_120__77_, s_r_120__76_, s_r_120__75_, s_r_120__74_, s_r_120__73_, s_r_120__72_, s_r_120__71_, s_r_120__70_, s_r_120__69_, s_r_120__68_, s_r_120__67_, s_r_120__66_, s_r_120__65_, s_r_120__64_, s_r_120__63_, s_r_120__62_, s_r_120__61_, s_r_120__60_, s_r_120__59_, s_r_120__58_, s_r_120__57_, s_r_120__56_, s_r_120__55_, s_r_120__54_, s_r_120__53_, s_r_120__52_, s_r_120__51_, s_r_120__50_, s_r_120__49_, s_r_120__48_, s_r_120__47_, s_r_120__46_, s_r_120__45_, s_r_120__44_, s_r_120__43_, s_r_120__42_, s_r_120__41_, s_r_120__40_, s_r_120__39_, s_r_120__38_, s_r_120__37_, s_r_120__36_, s_r_120__35_, s_r_120__34_, s_r_120__33_, s_r_120__32_, s_r_120__31_, s_r_120__30_, s_r_120__29_, s_r_120__28_, s_r_120__27_, s_r_120__26_, s_r_120__25_, s_r_120__24_, s_r_120__23_, s_r_120__22_, s_r_120__21_, s_r_120__20_, s_r_120__19_, s_r_120__18_, s_r_120__17_, s_r_120__16_, s_r_120__15_, s_r_120__14_, s_r_120__13_, s_r_120__12_, s_r_120__11_, s_r_120__10_, s_r_120__9_, s_r_120__8_, s_r_120__7_, s_r_120__6_, s_r_120__5_, s_r_120__4_, s_r_120__3_, s_r_120__2_, s_r_120__1_, s_r_120__0_ }),
    .c_o(c_r[120]),
    .prod_accum_o({ prod_accum_120__121_, prod_accum_120__120_, prod_accum_120__119_, prod_accum_120__118_, prod_accum_120__117_, prod_accum_120__116_, prod_accum_120__115_, prod_accum_120__114_, prod_accum_120__113_, prod_accum_120__112_, prod_accum_120__111_, prod_accum_120__110_, prod_accum_120__109_, prod_accum_120__108_, prod_accum_120__107_, prod_accum_120__106_, prod_accum_120__105_, prod_accum_120__104_, prod_accum_120__103_, prod_accum_120__102_, prod_accum_120__101_, prod_accum_120__100_, prod_accum_120__99_, prod_accum_120__98_, prod_accum_120__97_, prod_accum_120__96_, prod_accum_120__95_, prod_accum_120__94_, prod_accum_120__93_, prod_accum_120__92_, prod_accum_120__91_, prod_accum_120__90_, prod_accum_120__89_, prod_accum_120__88_, prod_accum_120__87_, prod_accum_120__86_, prod_accum_120__85_, prod_accum_120__84_, prod_accum_120__83_, prod_accum_120__82_, prod_accum_120__81_, prod_accum_120__80_, prod_accum_120__79_, prod_accum_120__78_, prod_accum_120__77_, prod_accum_120__76_, prod_accum_120__75_, prod_accum_120__74_, prod_accum_120__73_, prod_accum_120__72_, prod_accum_120__71_, prod_accum_120__70_, prod_accum_120__69_, prod_accum_120__68_, prod_accum_120__67_, prod_accum_120__66_, prod_accum_120__65_, prod_accum_120__64_, prod_accum_120__63_, prod_accum_120__62_, prod_accum_120__61_, prod_accum_120__60_, prod_accum_120__59_, prod_accum_120__58_, prod_accum_120__57_, prod_accum_120__56_, prod_accum_120__55_, prod_accum_120__54_, prod_accum_120__53_, prod_accum_120__52_, prod_accum_120__51_, prod_accum_120__50_, prod_accum_120__49_, prod_accum_120__48_, prod_accum_120__47_, prod_accum_120__46_, prod_accum_120__45_, prod_accum_120__44_, prod_accum_120__43_, prod_accum_120__42_, prod_accum_120__41_, prod_accum_120__40_, prod_accum_120__39_, prod_accum_120__38_, prod_accum_120__37_, prod_accum_120__36_, prod_accum_120__35_, prod_accum_120__34_, prod_accum_120__33_, prod_accum_120__32_, prod_accum_120__31_, prod_accum_120__30_, prod_accum_120__29_, prod_accum_120__28_, prod_accum_120__27_, prod_accum_120__26_, prod_accum_120__25_, prod_accum_120__24_, prod_accum_120__23_, prod_accum_120__22_, prod_accum_120__21_, prod_accum_120__20_, prod_accum_120__19_, prod_accum_120__18_, prod_accum_120__17_, prod_accum_120__16_, prod_accum_120__15_, prod_accum_120__14_, prod_accum_120__13_, prod_accum_120__12_, prod_accum_120__11_, prod_accum_120__10_, prod_accum_120__9_, prod_accum_120__8_, prod_accum_120__7_, prod_accum_120__6_, prod_accum_120__5_, prod_accum_120__4_, prod_accum_120__3_, prod_accum_120__2_, prod_accum_120__1_, prod_accum_120__0_ })
  );


  bsg_mul_array_row_128_121_x
  genblk1_121__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[15487:15360]),
    .b_i(b_r[15487:15360]),
    .s_i({ s_r_120__127_, s_r_120__126_, s_r_120__125_, s_r_120__124_, s_r_120__123_, s_r_120__122_, s_r_120__121_, s_r_120__120_, s_r_120__119_, s_r_120__118_, s_r_120__117_, s_r_120__116_, s_r_120__115_, s_r_120__114_, s_r_120__113_, s_r_120__112_, s_r_120__111_, s_r_120__110_, s_r_120__109_, s_r_120__108_, s_r_120__107_, s_r_120__106_, s_r_120__105_, s_r_120__104_, s_r_120__103_, s_r_120__102_, s_r_120__101_, s_r_120__100_, s_r_120__99_, s_r_120__98_, s_r_120__97_, s_r_120__96_, s_r_120__95_, s_r_120__94_, s_r_120__93_, s_r_120__92_, s_r_120__91_, s_r_120__90_, s_r_120__89_, s_r_120__88_, s_r_120__87_, s_r_120__86_, s_r_120__85_, s_r_120__84_, s_r_120__83_, s_r_120__82_, s_r_120__81_, s_r_120__80_, s_r_120__79_, s_r_120__78_, s_r_120__77_, s_r_120__76_, s_r_120__75_, s_r_120__74_, s_r_120__73_, s_r_120__72_, s_r_120__71_, s_r_120__70_, s_r_120__69_, s_r_120__68_, s_r_120__67_, s_r_120__66_, s_r_120__65_, s_r_120__64_, s_r_120__63_, s_r_120__62_, s_r_120__61_, s_r_120__60_, s_r_120__59_, s_r_120__58_, s_r_120__57_, s_r_120__56_, s_r_120__55_, s_r_120__54_, s_r_120__53_, s_r_120__52_, s_r_120__51_, s_r_120__50_, s_r_120__49_, s_r_120__48_, s_r_120__47_, s_r_120__46_, s_r_120__45_, s_r_120__44_, s_r_120__43_, s_r_120__42_, s_r_120__41_, s_r_120__40_, s_r_120__39_, s_r_120__38_, s_r_120__37_, s_r_120__36_, s_r_120__35_, s_r_120__34_, s_r_120__33_, s_r_120__32_, s_r_120__31_, s_r_120__30_, s_r_120__29_, s_r_120__28_, s_r_120__27_, s_r_120__26_, s_r_120__25_, s_r_120__24_, s_r_120__23_, s_r_120__22_, s_r_120__21_, s_r_120__20_, s_r_120__19_, s_r_120__18_, s_r_120__17_, s_r_120__16_, s_r_120__15_, s_r_120__14_, s_r_120__13_, s_r_120__12_, s_r_120__11_, s_r_120__10_, s_r_120__9_, s_r_120__8_, s_r_120__7_, s_r_120__6_, s_r_120__5_, s_r_120__4_, s_r_120__3_, s_r_120__2_, s_r_120__1_, s_r_120__0_ }),
    .c_i(c_r[120]),
    .prod_accum_i({ prod_accum_120__121_, prod_accum_120__120_, prod_accum_120__119_, prod_accum_120__118_, prod_accum_120__117_, prod_accum_120__116_, prod_accum_120__115_, prod_accum_120__114_, prod_accum_120__113_, prod_accum_120__112_, prod_accum_120__111_, prod_accum_120__110_, prod_accum_120__109_, prod_accum_120__108_, prod_accum_120__107_, prod_accum_120__106_, prod_accum_120__105_, prod_accum_120__104_, prod_accum_120__103_, prod_accum_120__102_, prod_accum_120__101_, prod_accum_120__100_, prod_accum_120__99_, prod_accum_120__98_, prod_accum_120__97_, prod_accum_120__96_, prod_accum_120__95_, prod_accum_120__94_, prod_accum_120__93_, prod_accum_120__92_, prod_accum_120__91_, prod_accum_120__90_, prod_accum_120__89_, prod_accum_120__88_, prod_accum_120__87_, prod_accum_120__86_, prod_accum_120__85_, prod_accum_120__84_, prod_accum_120__83_, prod_accum_120__82_, prod_accum_120__81_, prod_accum_120__80_, prod_accum_120__79_, prod_accum_120__78_, prod_accum_120__77_, prod_accum_120__76_, prod_accum_120__75_, prod_accum_120__74_, prod_accum_120__73_, prod_accum_120__72_, prod_accum_120__71_, prod_accum_120__70_, prod_accum_120__69_, prod_accum_120__68_, prod_accum_120__67_, prod_accum_120__66_, prod_accum_120__65_, prod_accum_120__64_, prod_accum_120__63_, prod_accum_120__62_, prod_accum_120__61_, prod_accum_120__60_, prod_accum_120__59_, prod_accum_120__58_, prod_accum_120__57_, prod_accum_120__56_, prod_accum_120__55_, prod_accum_120__54_, prod_accum_120__53_, prod_accum_120__52_, prod_accum_120__51_, prod_accum_120__50_, prod_accum_120__49_, prod_accum_120__48_, prod_accum_120__47_, prod_accum_120__46_, prod_accum_120__45_, prod_accum_120__44_, prod_accum_120__43_, prod_accum_120__42_, prod_accum_120__41_, prod_accum_120__40_, prod_accum_120__39_, prod_accum_120__38_, prod_accum_120__37_, prod_accum_120__36_, prod_accum_120__35_, prod_accum_120__34_, prod_accum_120__33_, prod_accum_120__32_, prod_accum_120__31_, prod_accum_120__30_, prod_accum_120__29_, prod_accum_120__28_, prod_accum_120__27_, prod_accum_120__26_, prod_accum_120__25_, prod_accum_120__24_, prod_accum_120__23_, prod_accum_120__22_, prod_accum_120__21_, prod_accum_120__20_, prod_accum_120__19_, prod_accum_120__18_, prod_accum_120__17_, prod_accum_120__16_, prod_accum_120__15_, prod_accum_120__14_, prod_accum_120__13_, prod_accum_120__12_, prod_accum_120__11_, prod_accum_120__10_, prod_accum_120__9_, prod_accum_120__8_, prod_accum_120__7_, prod_accum_120__6_, prod_accum_120__5_, prod_accum_120__4_, prod_accum_120__3_, prod_accum_120__2_, prod_accum_120__1_, prod_accum_120__0_ }),
    .a_o(a_r[15615:15488]),
    .b_o(b_r[15615:15488]),
    .s_o({ s_r_121__127_, s_r_121__126_, s_r_121__125_, s_r_121__124_, s_r_121__123_, s_r_121__122_, s_r_121__121_, s_r_121__120_, s_r_121__119_, s_r_121__118_, s_r_121__117_, s_r_121__116_, s_r_121__115_, s_r_121__114_, s_r_121__113_, s_r_121__112_, s_r_121__111_, s_r_121__110_, s_r_121__109_, s_r_121__108_, s_r_121__107_, s_r_121__106_, s_r_121__105_, s_r_121__104_, s_r_121__103_, s_r_121__102_, s_r_121__101_, s_r_121__100_, s_r_121__99_, s_r_121__98_, s_r_121__97_, s_r_121__96_, s_r_121__95_, s_r_121__94_, s_r_121__93_, s_r_121__92_, s_r_121__91_, s_r_121__90_, s_r_121__89_, s_r_121__88_, s_r_121__87_, s_r_121__86_, s_r_121__85_, s_r_121__84_, s_r_121__83_, s_r_121__82_, s_r_121__81_, s_r_121__80_, s_r_121__79_, s_r_121__78_, s_r_121__77_, s_r_121__76_, s_r_121__75_, s_r_121__74_, s_r_121__73_, s_r_121__72_, s_r_121__71_, s_r_121__70_, s_r_121__69_, s_r_121__68_, s_r_121__67_, s_r_121__66_, s_r_121__65_, s_r_121__64_, s_r_121__63_, s_r_121__62_, s_r_121__61_, s_r_121__60_, s_r_121__59_, s_r_121__58_, s_r_121__57_, s_r_121__56_, s_r_121__55_, s_r_121__54_, s_r_121__53_, s_r_121__52_, s_r_121__51_, s_r_121__50_, s_r_121__49_, s_r_121__48_, s_r_121__47_, s_r_121__46_, s_r_121__45_, s_r_121__44_, s_r_121__43_, s_r_121__42_, s_r_121__41_, s_r_121__40_, s_r_121__39_, s_r_121__38_, s_r_121__37_, s_r_121__36_, s_r_121__35_, s_r_121__34_, s_r_121__33_, s_r_121__32_, s_r_121__31_, s_r_121__30_, s_r_121__29_, s_r_121__28_, s_r_121__27_, s_r_121__26_, s_r_121__25_, s_r_121__24_, s_r_121__23_, s_r_121__22_, s_r_121__21_, s_r_121__20_, s_r_121__19_, s_r_121__18_, s_r_121__17_, s_r_121__16_, s_r_121__15_, s_r_121__14_, s_r_121__13_, s_r_121__12_, s_r_121__11_, s_r_121__10_, s_r_121__9_, s_r_121__8_, s_r_121__7_, s_r_121__6_, s_r_121__5_, s_r_121__4_, s_r_121__3_, s_r_121__2_, s_r_121__1_, s_r_121__0_ }),
    .c_o(c_r[121]),
    .prod_accum_o({ prod_accum_121__122_, prod_accum_121__121_, prod_accum_121__120_, prod_accum_121__119_, prod_accum_121__118_, prod_accum_121__117_, prod_accum_121__116_, prod_accum_121__115_, prod_accum_121__114_, prod_accum_121__113_, prod_accum_121__112_, prod_accum_121__111_, prod_accum_121__110_, prod_accum_121__109_, prod_accum_121__108_, prod_accum_121__107_, prod_accum_121__106_, prod_accum_121__105_, prod_accum_121__104_, prod_accum_121__103_, prod_accum_121__102_, prod_accum_121__101_, prod_accum_121__100_, prod_accum_121__99_, prod_accum_121__98_, prod_accum_121__97_, prod_accum_121__96_, prod_accum_121__95_, prod_accum_121__94_, prod_accum_121__93_, prod_accum_121__92_, prod_accum_121__91_, prod_accum_121__90_, prod_accum_121__89_, prod_accum_121__88_, prod_accum_121__87_, prod_accum_121__86_, prod_accum_121__85_, prod_accum_121__84_, prod_accum_121__83_, prod_accum_121__82_, prod_accum_121__81_, prod_accum_121__80_, prod_accum_121__79_, prod_accum_121__78_, prod_accum_121__77_, prod_accum_121__76_, prod_accum_121__75_, prod_accum_121__74_, prod_accum_121__73_, prod_accum_121__72_, prod_accum_121__71_, prod_accum_121__70_, prod_accum_121__69_, prod_accum_121__68_, prod_accum_121__67_, prod_accum_121__66_, prod_accum_121__65_, prod_accum_121__64_, prod_accum_121__63_, prod_accum_121__62_, prod_accum_121__61_, prod_accum_121__60_, prod_accum_121__59_, prod_accum_121__58_, prod_accum_121__57_, prod_accum_121__56_, prod_accum_121__55_, prod_accum_121__54_, prod_accum_121__53_, prod_accum_121__52_, prod_accum_121__51_, prod_accum_121__50_, prod_accum_121__49_, prod_accum_121__48_, prod_accum_121__47_, prod_accum_121__46_, prod_accum_121__45_, prod_accum_121__44_, prod_accum_121__43_, prod_accum_121__42_, prod_accum_121__41_, prod_accum_121__40_, prod_accum_121__39_, prod_accum_121__38_, prod_accum_121__37_, prod_accum_121__36_, prod_accum_121__35_, prod_accum_121__34_, prod_accum_121__33_, prod_accum_121__32_, prod_accum_121__31_, prod_accum_121__30_, prod_accum_121__29_, prod_accum_121__28_, prod_accum_121__27_, prod_accum_121__26_, prod_accum_121__25_, prod_accum_121__24_, prod_accum_121__23_, prod_accum_121__22_, prod_accum_121__21_, prod_accum_121__20_, prod_accum_121__19_, prod_accum_121__18_, prod_accum_121__17_, prod_accum_121__16_, prod_accum_121__15_, prod_accum_121__14_, prod_accum_121__13_, prod_accum_121__12_, prod_accum_121__11_, prod_accum_121__10_, prod_accum_121__9_, prod_accum_121__8_, prod_accum_121__7_, prod_accum_121__6_, prod_accum_121__5_, prod_accum_121__4_, prod_accum_121__3_, prod_accum_121__2_, prod_accum_121__1_, prod_accum_121__0_ })
  );


  bsg_mul_array_row_128_122_x
  genblk1_122__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[15615:15488]),
    .b_i(b_r[15615:15488]),
    .s_i({ s_r_121__127_, s_r_121__126_, s_r_121__125_, s_r_121__124_, s_r_121__123_, s_r_121__122_, s_r_121__121_, s_r_121__120_, s_r_121__119_, s_r_121__118_, s_r_121__117_, s_r_121__116_, s_r_121__115_, s_r_121__114_, s_r_121__113_, s_r_121__112_, s_r_121__111_, s_r_121__110_, s_r_121__109_, s_r_121__108_, s_r_121__107_, s_r_121__106_, s_r_121__105_, s_r_121__104_, s_r_121__103_, s_r_121__102_, s_r_121__101_, s_r_121__100_, s_r_121__99_, s_r_121__98_, s_r_121__97_, s_r_121__96_, s_r_121__95_, s_r_121__94_, s_r_121__93_, s_r_121__92_, s_r_121__91_, s_r_121__90_, s_r_121__89_, s_r_121__88_, s_r_121__87_, s_r_121__86_, s_r_121__85_, s_r_121__84_, s_r_121__83_, s_r_121__82_, s_r_121__81_, s_r_121__80_, s_r_121__79_, s_r_121__78_, s_r_121__77_, s_r_121__76_, s_r_121__75_, s_r_121__74_, s_r_121__73_, s_r_121__72_, s_r_121__71_, s_r_121__70_, s_r_121__69_, s_r_121__68_, s_r_121__67_, s_r_121__66_, s_r_121__65_, s_r_121__64_, s_r_121__63_, s_r_121__62_, s_r_121__61_, s_r_121__60_, s_r_121__59_, s_r_121__58_, s_r_121__57_, s_r_121__56_, s_r_121__55_, s_r_121__54_, s_r_121__53_, s_r_121__52_, s_r_121__51_, s_r_121__50_, s_r_121__49_, s_r_121__48_, s_r_121__47_, s_r_121__46_, s_r_121__45_, s_r_121__44_, s_r_121__43_, s_r_121__42_, s_r_121__41_, s_r_121__40_, s_r_121__39_, s_r_121__38_, s_r_121__37_, s_r_121__36_, s_r_121__35_, s_r_121__34_, s_r_121__33_, s_r_121__32_, s_r_121__31_, s_r_121__30_, s_r_121__29_, s_r_121__28_, s_r_121__27_, s_r_121__26_, s_r_121__25_, s_r_121__24_, s_r_121__23_, s_r_121__22_, s_r_121__21_, s_r_121__20_, s_r_121__19_, s_r_121__18_, s_r_121__17_, s_r_121__16_, s_r_121__15_, s_r_121__14_, s_r_121__13_, s_r_121__12_, s_r_121__11_, s_r_121__10_, s_r_121__9_, s_r_121__8_, s_r_121__7_, s_r_121__6_, s_r_121__5_, s_r_121__4_, s_r_121__3_, s_r_121__2_, s_r_121__1_, s_r_121__0_ }),
    .c_i(c_r[121]),
    .prod_accum_i({ prod_accum_121__122_, prod_accum_121__121_, prod_accum_121__120_, prod_accum_121__119_, prod_accum_121__118_, prod_accum_121__117_, prod_accum_121__116_, prod_accum_121__115_, prod_accum_121__114_, prod_accum_121__113_, prod_accum_121__112_, prod_accum_121__111_, prod_accum_121__110_, prod_accum_121__109_, prod_accum_121__108_, prod_accum_121__107_, prod_accum_121__106_, prod_accum_121__105_, prod_accum_121__104_, prod_accum_121__103_, prod_accum_121__102_, prod_accum_121__101_, prod_accum_121__100_, prod_accum_121__99_, prod_accum_121__98_, prod_accum_121__97_, prod_accum_121__96_, prod_accum_121__95_, prod_accum_121__94_, prod_accum_121__93_, prod_accum_121__92_, prod_accum_121__91_, prod_accum_121__90_, prod_accum_121__89_, prod_accum_121__88_, prod_accum_121__87_, prod_accum_121__86_, prod_accum_121__85_, prod_accum_121__84_, prod_accum_121__83_, prod_accum_121__82_, prod_accum_121__81_, prod_accum_121__80_, prod_accum_121__79_, prod_accum_121__78_, prod_accum_121__77_, prod_accum_121__76_, prod_accum_121__75_, prod_accum_121__74_, prod_accum_121__73_, prod_accum_121__72_, prod_accum_121__71_, prod_accum_121__70_, prod_accum_121__69_, prod_accum_121__68_, prod_accum_121__67_, prod_accum_121__66_, prod_accum_121__65_, prod_accum_121__64_, prod_accum_121__63_, prod_accum_121__62_, prod_accum_121__61_, prod_accum_121__60_, prod_accum_121__59_, prod_accum_121__58_, prod_accum_121__57_, prod_accum_121__56_, prod_accum_121__55_, prod_accum_121__54_, prod_accum_121__53_, prod_accum_121__52_, prod_accum_121__51_, prod_accum_121__50_, prod_accum_121__49_, prod_accum_121__48_, prod_accum_121__47_, prod_accum_121__46_, prod_accum_121__45_, prod_accum_121__44_, prod_accum_121__43_, prod_accum_121__42_, prod_accum_121__41_, prod_accum_121__40_, prod_accum_121__39_, prod_accum_121__38_, prod_accum_121__37_, prod_accum_121__36_, prod_accum_121__35_, prod_accum_121__34_, prod_accum_121__33_, prod_accum_121__32_, prod_accum_121__31_, prod_accum_121__30_, prod_accum_121__29_, prod_accum_121__28_, prod_accum_121__27_, prod_accum_121__26_, prod_accum_121__25_, prod_accum_121__24_, prod_accum_121__23_, prod_accum_121__22_, prod_accum_121__21_, prod_accum_121__20_, prod_accum_121__19_, prod_accum_121__18_, prod_accum_121__17_, prod_accum_121__16_, prod_accum_121__15_, prod_accum_121__14_, prod_accum_121__13_, prod_accum_121__12_, prod_accum_121__11_, prod_accum_121__10_, prod_accum_121__9_, prod_accum_121__8_, prod_accum_121__7_, prod_accum_121__6_, prod_accum_121__5_, prod_accum_121__4_, prod_accum_121__3_, prod_accum_121__2_, prod_accum_121__1_, prod_accum_121__0_ }),
    .a_o(a_r[15743:15616]),
    .b_o(b_r[15743:15616]),
    .s_o({ s_r_122__127_, s_r_122__126_, s_r_122__125_, s_r_122__124_, s_r_122__123_, s_r_122__122_, s_r_122__121_, s_r_122__120_, s_r_122__119_, s_r_122__118_, s_r_122__117_, s_r_122__116_, s_r_122__115_, s_r_122__114_, s_r_122__113_, s_r_122__112_, s_r_122__111_, s_r_122__110_, s_r_122__109_, s_r_122__108_, s_r_122__107_, s_r_122__106_, s_r_122__105_, s_r_122__104_, s_r_122__103_, s_r_122__102_, s_r_122__101_, s_r_122__100_, s_r_122__99_, s_r_122__98_, s_r_122__97_, s_r_122__96_, s_r_122__95_, s_r_122__94_, s_r_122__93_, s_r_122__92_, s_r_122__91_, s_r_122__90_, s_r_122__89_, s_r_122__88_, s_r_122__87_, s_r_122__86_, s_r_122__85_, s_r_122__84_, s_r_122__83_, s_r_122__82_, s_r_122__81_, s_r_122__80_, s_r_122__79_, s_r_122__78_, s_r_122__77_, s_r_122__76_, s_r_122__75_, s_r_122__74_, s_r_122__73_, s_r_122__72_, s_r_122__71_, s_r_122__70_, s_r_122__69_, s_r_122__68_, s_r_122__67_, s_r_122__66_, s_r_122__65_, s_r_122__64_, s_r_122__63_, s_r_122__62_, s_r_122__61_, s_r_122__60_, s_r_122__59_, s_r_122__58_, s_r_122__57_, s_r_122__56_, s_r_122__55_, s_r_122__54_, s_r_122__53_, s_r_122__52_, s_r_122__51_, s_r_122__50_, s_r_122__49_, s_r_122__48_, s_r_122__47_, s_r_122__46_, s_r_122__45_, s_r_122__44_, s_r_122__43_, s_r_122__42_, s_r_122__41_, s_r_122__40_, s_r_122__39_, s_r_122__38_, s_r_122__37_, s_r_122__36_, s_r_122__35_, s_r_122__34_, s_r_122__33_, s_r_122__32_, s_r_122__31_, s_r_122__30_, s_r_122__29_, s_r_122__28_, s_r_122__27_, s_r_122__26_, s_r_122__25_, s_r_122__24_, s_r_122__23_, s_r_122__22_, s_r_122__21_, s_r_122__20_, s_r_122__19_, s_r_122__18_, s_r_122__17_, s_r_122__16_, s_r_122__15_, s_r_122__14_, s_r_122__13_, s_r_122__12_, s_r_122__11_, s_r_122__10_, s_r_122__9_, s_r_122__8_, s_r_122__7_, s_r_122__6_, s_r_122__5_, s_r_122__4_, s_r_122__3_, s_r_122__2_, s_r_122__1_, s_r_122__0_ }),
    .c_o(c_r[122]),
    .prod_accum_o({ prod_accum_122__123_, prod_accum_122__122_, prod_accum_122__121_, prod_accum_122__120_, prod_accum_122__119_, prod_accum_122__118_, prod_accum_122__117_, prod_accum_122__116_, prod_accum_122__115_, prod_accum_122__114_, prod_accum_122__113_, prod_accum_122__112_, prod_accum_122__111_, prod_accum_122__110_, prod_accum_122__109_, prod_accum_122__108_, prod_accum_122__107_, prod_accum_122__106_, prod_accum_122__105_, prod_accum_122__104_, prod_accum_122__103_, prod_accum_122__102_, prod_accum_122__101_, prod_accum_122__100_, prod_accum_122__99_, prod_accum_122__98_, prod_accum_122__97_, prod_accum_122__96_, prod_accum_122__95_, prod_accum_122__94_, prod_accum_122__93_, prod_accum_122__92_, prod_accum_122__91_, prod_accum_122__90_, prod_accum_122__89_, prod_accum_122__88_, prod_accum_122__87_, prod_accum_122__86_, prod_accum_122__85_, prod_accum_122__84_, prod_accum_122__83_, prod_accum_122__82_, prod_accum_122__81_, prod_accum_122__80_, prod_accum_122__79_, prod_accum_122__78_, prod_accum_122__77_, prod_accum_122__76_, prod_accum_122__75_, prod_accum_122__74_, prod_accum_122__73_, prod_accum_122__72_, prod_accum_122__71_, prod_accum_122__70_, prod_accum_122__69_, prod_accum_122__68_, prod_accum_122__67_, prod_accum_122__66_, prod_accum_122__65_, prod_accum_122__64_, prod_accum_122__63_, prod_accum_122__62_, prod_accum_122__61_, prod_accum_122__60_, prod_accum_122__59_, prod_accum_122__58_, prod_accum_122__57_, prod_accum_122__56_, prod_accum_122__55_, prod_accum_122__54_, prod_accum_122__53_, prod_accum_122__52_, prod_accum_122__51_, prod_accum_122__50_, prod_accum_122__49_, prod_accum_122__48_, prod_accum_122__47_, prod_accum_122__46_, prod_accum_122__45_, prod_accum_122__44_, prod_accum_122__43_, prod_accum_122__42_, prod_accum_122__41_, prod_accum_122__40_, prod_accum_122__39_, prod_accum_122__38_, prod_accum_122__37_, prod_accum_122__36_, prod_accum_122__35_, prod_accum_122__34_, prod_accum_122__33_, prod_accum_122__32_, prod_accum_122__31_, prod_accum_122__30_, prod_accum_122__29_, prod_accum_122__28_, prod_accum_122__27_, prod_accum_122__26_, prod_accum_122__25_, prod_accum_122__24_, prod_accum_122__23_, prod_accum_122__22_, prod_accum_122__21_, prod_accum_122__20_, prod_accum_122__19_, prod_accum_122__18_, prod_accum_122__17_, prod_accum_122__16_, prod_accum_122__15_, prod_accum_122__14_, prod_accum_122__13_, prod_accum_122__12_, prod_accum_122__11_, prod_accum_122__10_, prod_accum_122__9_, prod_accum_122__8_, prod_accum_122__7_, prod_accum_122__6_, prod_accum_122__5_, prod_accum_122__4_, prod_accum_122__3_, prod_accum_122__2_, prod_accum_122__1_, prod_accum_122__0_ })
  );


  bsg_mul_array_row_128_123_x
  genblk1_123__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[15743:15616]),
    .b_i(b_r[15743:15616]),
    .s_i({ s_r_122__127_, s_r_122__126_, s_r_122__125_, s_r_122__124_, s_r_122__123_, s_r_122__122_, s_r_122__121_, s_r_122__120_, s_r_122__119_, s_r_122__118_, s_r_122__117_, s_r_122__116_, s_r_122__115_, s_r_122__114_, s_r_122__113_, s_r_122__112_, s_r_122__111_, s_r_122__110_, s_r_122__109_, s_r_122__108_, s_r_122__107_, s_r_122__106_, s_r_122__105_, s_r_122__104_, s_r_122__103_, s_r_122__102_, s_r_122__101_, s_r_122__100_, s_r_122__99_, s_r_122__98_, s_r_122__97_, s_r_122__96_, s_r_122__95_, s_r_122__94_, s_r_122__93_, s_r_122__92_, s_r_122__91_, s_r_122__90_, s_r_122__89_, s_r_122__88_, s_r_122__87_, s_r_122__86_, s_r_122__85_, s_r_122__84_, s_r_122__83_, s_r_122__82_, s_r_122__81_, s_r_122__80_, s_r_122__79_, s_r_122__78_, s_r_122__77_, s_r_122__76_, s_r_122__75_, s_r_122__74_, s_r_122__73_, s_r_122__72_, s_r_122__71_, s_r_122__70_, s_r_122__69_, s_r_122__68_, s_r_122__67_, s_r_122__66_, s_r_122__65_, s_r_122__64_, s_r_122__63_, s_r_122__62_, s_r_122__61_, s_r_122__60_, s_r_122__59_, s_r_122__58_, s_r_122__57_, s_r_122__56_, s_r_122__55_, s_r_122__54_, s_r_122__53_, s_r_122__52_, s_r_122__51_, s_r_122__50_, s_r_122__49_, s_r_122__48_, s_r_122__47_, s_r_122__46_, s_r_122__45_, s_r_122__44_, s_r_122__43_, s_r_122__42_, s_r_122__41_, s_r_122__40_, s_r_122__39_, s_r_122__38_, s_r_122__37_, s_r_122__36_, s_r_122__35_, s_r_122__34_, s_r_122__33_, s_r_122__32_, s_r_122__31_, s_r_122__30_, s_r_122__29_, s_r_122__28_, s_r_122__27_, s_r_122__26_, s_r_122__25_, s_r_122__24_, s_r_122__23_, s_r_122__22_, s_r_122__21_, s_r_122__20_, s_r_122__19_, s_r_122__18_, s_r_122__17_, s_r_122__16_, s_r_122__15_, s_r_122__14_, s_r_122__13_, s_r_122__12_, s_r_122__11_, s_r_122__10_, s_r_122__9_, s_r_122__8_, s_r_122__7_, s_r_122__6_, s_r_122__5_, s_r_122__4_, s_r_122__3_, s_r_122__2_, s_r_122__1_, s_r_122__0_ }),
    .c_i(c_r[122]),
    .prod_accum_i({ prod_accum_122__123_, prod_accum_122__122_, prod_accum_122__121_, prod_accum_122__120_, prod_accum_122__119_, prod_accum_122__118_, prod_accum_122__117_, prod_accum_122__116_, prod_accum_122__115_, prod_accum_122__114_, prod_accum_122__113_, prod_accum_122__112_, prod_accum_122__111_, prod_accum_122__110_, prod_accum_122__109_, prod_accum_122__108_, prod_accum_122__107_, prod_accum_122__106_, prod_accum_122__105_, prod_accum_122__104_, prod_accum_122__103_, prod_accum_122__102_, prod_accum_122__101_, prod_accum_122__100_, prod_accum_122__99_, prod_accum_122__98_, prod_accum_122__97_, prod_accum_122__96_, prod_accum_122__95_, prod_accum_122__94_, prod_accum_122__93_, prod_accum_122__92_, prod_accum_122__91_, prod_accum_122__90_, prod_accum_122__89_, prod_accum_122__88_, prod_accum_122__87_, prod_accum_122__86_, prod_accum_122__85_, prod_accum_122__84_, prod_accum_122__83_, prod_accum_122__82_, prod_accum_122__81_, prod_accum_122__80_, prod_accum_122__79_, prod_accum_122__78_, prod_accum_122__77_, prod_accum_122__76_, prod_accum_122__75_, prod_accum_122__74_, prod_accum_122__73_, prod_accum_122__72_, prod_accum_122__71_, prod_accum_122__70_, prod_accum_122__69_, prod_accum_122__68_, prod_accum_122__67_, prod_accum_122__66_, prod_accum_122__65_, prod_accum_122__64_, prod_accum_122__63_, prod_accum_122__62_, prod_accum_122__61_, prod_accum_122__60_, prod_accum_122__59_, prod_accum_122__58_, prod_accum_122__57_, prod_accum_122__56_, prod_accum_122__55_, prod_accum_122__54_, prod_accum_122__53_, prod_accum_122__52_, prod_accum_122__51_, prod_accum_122__50_, prod_accum_122__49_, prod_accum_122__48_, prod_accum_122__47_, prod_accum_122__46_, prod_accum_122__45_, prod_accum_122__44_, prod_accum_122__43_, prod_accum_122__42_, prod_accum_122__41_, prod_accum_122__40_, prod_accum_122__39_, prod_accum_122__38_, prod_accum_122__37_, prod_accum_122__36_, prod_accum_122__35_, prod_accum_122__34_, prod_accum_122__33_, prod_accum_122__32_, prod_accum_122__31_, prod_accum_122__30_, prod_accum_122__29_, prod_accum_122__28_, prod_accum_122__27_, prod_accum_122__26_, prod_accum_122__25_, prod_accum_122__24_, prod_accum_122__23_, prod_accum_122__22_, prod_accum_122__21_, prod_accum_122__20_, prod_accum_122__19_, prod_accum_122__18_, prod_accum_122__17_, prod_accum_122__16_, prod_accum_122__15_, prod_accum_122__14_, prod_accum_122__13_, prod_accum_122__12_, prod_accum_122__11_, prod_accum_122__10_, prod_accum_122__9_, prod_accum_122__8_, prod_accum_122__7_, prod_accum_122__6_, prod_accum_122__5_, prod_accum_122__4_, prod_accum_122__3_, prod_accum_122__2_, prod_accum_122__1_, prod_accum_122__0_ }),
    .a_o(a_r[15871:15744]),
    .b_o(b_r[15871:15744]),
    .s_o({ s_r_123__127_, s_r_123__126_, s_r_123__125_, s_r_123__124_, s_r_123__123_, s_r_123__122_, s_r_123__121_, s_r_123__120_, s_r_123__119_, s_r_123__118_, s_r_123__117_, s_r_123__116_, s_r_123__115_, s_r_123__114_, s_r_123__113_, s_r_123__112_, s_r_123__111_, s_r_123__110_, s_r_123__109_, s_r_123__108_, s_r_123__107_, s_r_123__106_, s_r_123__105_, s_r_123__104_, s_r_123__103_, s_r_123__102_, s_r_123__101_, s_r_123__100_, s_r_123__99_, s_r_123__98_, s_r_123__97_, s_r_123__96_, s_r_123__95_, s_r_123__94_, s_r_123__93_, s_r_123__92_, s_r_123__91_, s_r_123__90_, s_r_123__89_, s_r_123__88_, s_r_123__87_, s_r_123__86_, s_r_123__85_, s_r_123__84_, s_r_123__83_, s_r_123__82_, s_r_123__81_, s_r_123__80_, s_r_123__79_, s_r_123__78_, s_r_123__77_, s_r_123__76_, s_r_123__75_, s_r_123__74_, s_r_123__73_, s_r_123__72_, s_r_123__71_, s_r_123__70_, s_r_123__69_, s_r_123__68_, s_r_123__67_, s_r_123__66_, s_r_123__65_, s_r_123__64_, s_r_123__63_, s_r_123__62_, s_r_123__61_, s_r_123__60_, s_r_123__59_, s_r_123__58_, s_r_123__57_, s_r_123__56_, s_r_123__55_, s_r_123__54_, s_r_123__53_, s_r_123__52_, s_r_123__51_, s_r_123__50_, s_r_123__49_, s_r_123__48_, s_r_123__47_, s_r_123__46_, s_r_123__45_, s_r_123__44_, s_r_123__43_, s_r_123__42_, s_r_123__41_, s_r_123__40_, s_r_123__39_, s_r_123__38_, s_r_123__37_, s_r_123__36_, s_r_123__35_, s_r_123__34_, s_r_123__33_, s_r_123__32_, s_r_123__31_, s_r_123__30_, s_r_123__29_, s_r_123__28_, s_r_123__27_, s_r_123__26_, s_r_123__25_, s_r_123__24_, s_r_123__23_, s_r_123__22_, s_r_123__21_, s_r_123__20_, s_r_123__19_, s_r_123__18_, s_r_123__17_, s_r_123__16_, s_r_123__15_, s_r_123__14_, s_r_123__13_, s_r_123__12_, s_r_123__11_, s_r_123__10_, s_r_123__9_, s_r_123__8_, s_r_123__7_, s_r_123__6_, s_r_123__5_, s_r_123__4_, s_r_123__3_, s_r_123__2_, s_r_123__1_, s_r_123__0_ }),
    .c_o(c_r[123]),
    .prod_accum_o({ prod_accum_123__124_, prod_accum_123__123_, prod_accum_123__122_, prod_accum_123__121_, prod_accum_123__120_, prod_accum_123__119_, prod_accum_123__118_, prod_accum_123__117_, prod_accum_123__116_, prod_accum_123__115_, prod_accum_123__114_, prod_accum_123__113_, prod_accum_123__112_, prod_accum_123__111_, prod_accum_123__110_, prod_accum_123__109_, prod_accum_123__108_, prod_accum_123__107_, prod_accum_123__106_, prod_accum_123__105_, prod_accum_123__104_, prod_accum_123__103_, prod_accum_123__102_, prod_accum_123__101_, prod_accum_123__100_, prod_accum_123__99_, prod_accum_123__98_, prod_accum_123__97_, prod_accum_123__96_, prod_accum_123__95_, prod_accum_123__94_, prod_accum_123__93_, prod_accum_123__92_, prod_accum_123__91_, prod_accum_123__90_, prod_accum_123__89_, prod_accum_123__88_, prod_accum_123__87_, prod_accum_123__86_, prod_accum_123__85_, prod_accum_123__84_, prod_accum_123__83_, prod_accum_123__82_, prod_accum_123__81_, prod_accum_123__80_, prod_accum_123__79_, prod_accum_123__78_, prod_accum_123__77_, prod_accum_123__76_, prod_accum_123__75_, prod_accum_123__74_, prod_accum_123__73_, prod_accum_123__72_, prod_accum_123__71_, prod_accum_123__70_, prod_accum_123__69_, prod_accum_123__68_, prod_accum_123__67_, prod_accum_123__66_, prod_accum_123__65_, prod_accum_123__64_, prod_accum_123__63_, prod_accum_123__62_, prod_accum_123__61_, prod_accum_123__60_, prod_accum_123__59_, prod_accum_123__58_, prod_accum_123__57_, prod_accum_123__56_, prod_accum_123__55_, prod_accum_123__54_, prod_accum_123__53_, prod_accum_123__52_, prod_accum_123__51_, prod_accum_123__50_, prod_accum_123__49_, prod_accum_123__48_, prod_accum_123__47_, prod_accum_123__46_, prod_accum_123__45_, prod_accum_123__44_, prod_accum_123__43_, prod_accum_123__42_, prod_accum_123__41_, prod_accum_123__40_, prod_accum_123__39_, prod_accum_123__38_, prod_accum_123__37_, prod_accum_123__36_, prod_accum_123__35_, prod_accum_123__34_, prod_accum_123__33_, prod_accum_123__32_, prod_accum_123__31_, prod_accum_123__30_, prod_accum_123__29_, prod_accum_123__28_, prod_accum_123__27_, prod_accum_123__26_, prod_accum_123__25_, prod_accum_123__24_, prod_accum_123__23_, prod_accum_123__22_, prod_accum_123__21_, prod_accum_123__20_, prod_accum_123__19_, prod_accum_123__18_, prod_accum_123__17_, prod_accum_123__16_, prod_accum_123__15_, prod_accum_123__14_, prod_accum_123__13_, prod_accum_123__12_, prod_accum_123__11_, prod_accum_123__10_, prod_accum_123__9_, prod_accum_123__8_, prod_accum_123__7_, prod_accum_123__6_, prod_accum_123__5_, prod_accum_123__4_, prod_accum_123__3_, prod_accum_123__2_, prod_accum_123__1_, prod_accum_123__0_ })
  );


  bsg_mul_array_row_128_124_x
  genblk1_124__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[15871:15744]),
    .b_i(b_r[15871:15744]),
    .s_i({ s_r_123__127_, s_r_123__126_, s_r_123__125_, s_r_123__124_, s_r_123__123_, s_r_123__122_, s_r_123__121_, s_r_123__120_, s_r_123__119_, s_r_123__118_, s_r_123__117_, s_r_123__116_, s_r_123__115_, s_r_123__114_, s_r_123__113_, s_r_123__112_, s_r_123__111_, s_r_123__110_, s_r_123__109_, s_r_123__108_, s_r_123__107_, s_r_123__106_, s_r_123__105_, s_r_123__104_, s_r_123__103_, s_r_123__102_, s_r_123__101_, s_r_123__100_, s_r_123__99_, s_r_123__98_, s_r_123__97_, s_r_123__96_, s_r_123__95_, s_r_123__94_, s_r_123__93_, s_r_123__92_, s_r_123__91_, s_r_123__90_, s_r_123__89_, s_r_123__88_, s_r_123__87_, s_r_123__86_, s_r_123__85_, s_r_123__84_, s_r_123__83_, s_r_123__82_, s_r_123__81_, s_r_123__80_, s_r_123__79_, s_r_123__78_, s_r_123__77_, s_r_123__76_, s_r_123__75_, s_r_123__74_, s_r_123__73_, s_r_123__72_, s_r_123__71_, s_r_123__70_, s_r_123__69_, s_r_123__68_, s_r_123__67_, s_r_123__66_, s_r_123__65_, s_r_123__64_, s_r_123__63_, s_r_123__62_, s_r_123__61_, s_r_123__60_, s_r_123__59_, s_r_123__58_, s_r_123__57_, s_r_123__56_, s_r_123__55_, s_r_123__54_, s_r_123__53_, s_r_123__52_, s_r_123__51_, s_r_123__50_, s_r_123__49_, s_r_123__48_, s_r_123__47_, s_r_123__46_, s_r_123__45_, s_r_123__44_, s_r_123__43_, s_r_123__42_, s_r_123__41_, s_r_123__40_, s_r_123__39_, s_r_123__38_, s_r_123__37_, s_r_123__36_, s_r_123__35_, s_r_123__34_, s_r_123__33_, s_r_123__32_, s_r_123__31_, s_r_123__30_, s_r_123__29_, s_r_123__28_, s_r_123__27_, s_r_123__26_, s_r_123__25_, s_r_123__24_, s_r_123__23_, s_r_123__22_, s_r_123__21_, s_r_123__20_, s_r_123__19_, s_r_123__18_, s_r_123__17_, s_r_123__16_, s_r_123__15_, s_r_123__14_, s_r_123__13_, s_r_123__12_, s_r_123__11_, s_r_123__10_, s_r_123__9_, s_r_123__8_, s_r_123__7_, s_r_123__6_, s_r_123__5_, s_r_123__4_, s_r_123__3_, s_r_123__2_, s_r_123__1_, s_r_123__0_ }),
    .c_i(c_r[123]),
    .prod_accum_i({ prod_accum_123__124_, prod_accum_123__123_, prod_accum_123__122_, prod_accum_123__121_, prod_accum_123__120_, prod_accum_123__119_, prod_accum_123__118_, prod_accum_123__117_, prod_accum_123__116_, prod_accum_123__115_, prod_accum_123__114_, prod_accum_123__113_, prod_accum_123__112_, prod_accum_123__111_, prod_accum_123__110_, prod_accum_123__109_, prod_accum_123__108_, prod_accum_123__107_, prod_accum_123__106_, prod_accum_123__105_, prod_accum_123__104_, prod_accum_123__103_, prod_accum_123__102_, prod_accum_123__101_, prod_accum_123__100_, prod_accum_123__99_, prod_accum_123__98_, prod_accum_123__97_, prod_accum_123__96_, prod_accum_123__95_, prod_accum_123__94_, prod_accum_123__93_, prod_accum_123__92_, prod_accum_123__91_, prod_accum_123__90_, prod_accum_123__89_, prod_accum_123__88_, prod_accum_123__87_, prod_accum_123__86_, prod_accum_123__85_, prod_accum_123__84_, prod_accum_123__83_, prod_accum_123__82_, prod_accum_123__81_, prod_accum_123__80_, prod_accum_123__79_, prod_accum_123__78_, prod_accum_123__77_, prod_accum_123__76_, prod_accum_123__75_, prod_accum_123__74_, prod_accum_123__73_, prod_accum_123__72_, prod_accum_123__71_, prod_accum_123__70_, prod_accum_123__69_, prod_accum_123__68_, prod_accum_123__67_, prod_accum_123__66_, prod_accum_123__65_, prod_accum_123__64_, prod_accum_123__63_, prod_accum_123__62_, prod_accum_123__61_, prod_accum_123__60_, prod_accum_123__59_, prod_accum_123__58_, prod_accum_123__57_, prod_accum_123__56_, prod_accum_123__55_, prod_accum_123__54_, prod_accum_123__53_, prod_accum_123__52_, prod_accum_123__51_, prod_accum_123__50_, prod_accum_123__49_, prod_accum_123__48_, prod_accum_123__47_, prod_accum_123__46_, prod_accum_123__45_, prod_accum_123__44_, prod_accum_123__43_, prod_accum_123__42_, prod_accum_123__41_, prod_accum_123__40_, prod_accum_123__39_, prod_accum_123__38_, prod_accum_123__37_, prod_accum_123__36_, prod_accum_123__35_, prod_accum_123__34_, prod_accum_123__33_, prod_accum_123__32_, prod_accum_123__31_, prod_accum_123__30_, prod_accum_123__29_, prod_accum_123__28_, prod_accum_123__27_, prod_accum_123__26_, prod_accum_123__25_, prod_accum_123__24_, prod_accum_123__23_, prod_accum_123__22_, prod_accum_123__21_, prod_accum_123__20_, prod_accum_123__19_, prod_accum_123__18_, prod_accum_123__17_, prod_accum_123__16_, prod_accum_123__15_, prod_accum_123__14_, prod_accum_123__13_, prod_accum_123__12_, prod_accum_123__11_, prod_accum_123__10_, prod_accum_123__9_, prod_accum_123__8_, prod_accum_123__7_, prod_accum_123__6_, prod_accum_123__5_, prod_accum_123__4_, prod_accum_123__3_, prod_accum_123__2_, prod_accum_123__1_, prod_accum_123__0_ }),
    .a_o(a_r[15999:15872]),
    .b_o(b_r[15999:15872]),
    .s_o({ s_r_124__127_, s_r_124__126_, s_r_124__125_, s_r_124__124_, s_r_124__123_, s_r_124__122_, s_r_124__121_, s_r_124__120_, s_r_124__119_, s_r_124__118_, s_r_124__117_, s_r_124__116_, s_r_124__115_, s_r_124__114_, s_r_124__113_, s_r_124__112_, s_r_124__111_, s_r_124__110_, s_r_124__109_, s_r_124__108_, s_r_124__107_, s_r_124__106_, s_r_124__105_, s_r_124__104_, s_r_124__103_, s_r_124__102_, s_r_124__101_, s_r_124__100_, s_r_124__99_, s_r_124__98_, s_r_124__97_, s_r_124__96_, s_r_124__95_, s_r_124__94_, s_r_124__93_, s_r_124__92_, s_r_124__91_, s_r_124__90_, s_r_124__89_, s_r_124__88_, s_r_124__87_, s_r_124__86_, s_r_124__85_, s_r_124__84_, s_r_124__83_, s_r_124__82_, s_r_124__81_, s_r_124__80_, s_r_124__79_, s_r_124__78_, s_r_124__77_, s_r_124__76_, s_r_124__75_, s_r_124__74_, s_r_124__73_, s_r_124__72_, s_r_124__71_, s_r_124__70_, s_r_124__69_, s_r_124__68_, s_r_124__67_, s_r_124__66_, s_r_124__65_, s_r_124__64_, s_r_124__63_, s_r_124__62_, s_r_124__61_, s_r_124__60_, s_r_124__59_, s_r_124__58_, s_r_124__57_, s_r_124__56_, s_r_124__55_, s_r_124__54_, s_r_124__53_, s_r_124__52_, s_r_124__51_, s_r_124__50_, s_r_124__49_, s_r_124__48_, s_r_124__47_, s_r_124__46_, s_r_124__45_, s_r_124__44_, s_r_124__43_, s_r_124__42_, s_r_124__41_, s_r_124__40_, s_r_124__39_, s_r_124__38_, s_r_124__37_, s_r_124__36_, s_r_124__35_, s_r_124__34_, s_r_124__33_, s_r_124__32_, s_r_124__31_, s_r_124__30_, s_r_124__29_, s_r_124__28_, s_r_124__27_, s_r_124__26_, s_r_124__25_, s_r_124__24_, s_r_124__23_, s_r_124__22_, s_r_124__21_, s_r_124__20_, s_r_124__19_, s_r_124__18_, s_r_124__17_, s_r_124__16_, s_r_124__15_, s_r_124__14_, s_r_124__13_, s_r_124__12_, s_r_124__11_, s_r_124__10_, s_r_124__9_, s_r_124__8_, s_r_124__7_, s_r_124__6_, s_r_124__5_, s_r_124__4_, s_r_124__3_, s_r_124__2_, s_r_124__1_, s_r_124__0_ }),
    .c_o(c_r[124]),
    .prod_accum_o({ prod_accum_124__125_, prod_accum_124__124_, prod_accum_124__123_, prod_accum_124__122_, prod_accum_124__121_, prod_accum_124__120_, prod_accum_124__119_, prod_accum_124__118_, prod_accum_124__117_, prod_accum_124__116_, prod_accum_124__115_, prod_accum_124__114_, prod_accum_124__113_, prod_accum_124__112_, prod_accum_124__111_, prod_accum_124__110_, prod_accum_124__109_, prod_accum_124__108_, prod_accum_124__107_, prod_accum_124__106_, prod_accum_124__105_, prod_accum_124__104_, prod_accum_124__103_, prod_accum_124__102_, prod_accum_124__101_, prod_accum_124__100_, prod_accum_124__99_, prod_accum_124__98_, prod_accum_124__97_, prod_accum_124__96_, prod_accum_124__95_, prod_accum_124__94_, prod_accum_124__93_, prod_accum_124__92_, prod_accum_124__91_, prod_accum_124__90_, prod_accum_124__89_, prod_accum_124__88_, prod_accum_124__87_, prod_accum_124__86_, prod_accum_124__85_, prod_accum_124__84_, prod_accum_124__83_, prod_accum_124__82_, prod_accum_124__81_, prod_accum_124__80_, prod_accum_124__79_, prod_accum_124__78_, prod_accum_124__77_, prod_accum_124__76_, prod_accum_124__75_, prod_accum_124__74_, prod_accum_124__73_, prod_accum_124__72_, prod_accum_124__71_, prod_accum_124__70_, prod_accum_124__69_, prod_accum_124__68_, prod_accum_124__67_, prod_accum_124__66_, prod_accum_124__65_, prod_accum_124__64_, prod_accum_124__63_, prod_accum_124__62_, prod_accum_124__61_, prod_accum_124__60_, prod_accum_124__59_, prod_accum_124__58_, prod_accum_124__57_, prod_accum_124__56_, prod_accum_124__55_, prod_accum_124__54_, prod_accum_124__53_, prod_accum_124__52_, prod_accum_124__51_, prod_accum_124__50_, prod_accum_124__49_, prod_accum_124__48_, prod_accum_124__47_, prod_accum_124__46_, prod_accum_124__45_, prod_accum_124__44_, prod_accum_124__43_, prod_accum_124__42_, prod_accum_124__41_, prod_accum_124__40_, prod_accum_124__39_, prod_accum_124__38_, prod_accum_124__37_, prod_accum_124__36_, prod_accum_124__35_, prod_accum_124__34_, prod_accum_124__33_, prod_accum_124__32_, prod_accum_124__31_, prod_accum_124__30_, prod_accum_124__29_, prod_accum_124__28_, prod_accum_124__27_, prod_accum_124__26_, prod_accum_124__25_, prod_accum_124__24_, prod_accum_124__23_, prod_accum_124__22_, prod_accum_124__21_, prod_accum_124__20_, prod_accum_124__19_, prod_accum_124__18_, prod_accum_124__17_, prod_accum_124__16_, prod_accum_124__15_, prod_accum_124__14_, prod_accum_124__13_, prod_accum_124__12_, prod_accum_124__11_, prod_accum_124__10_, prod_accum_124__9_, prod_accum_124__8_, prod_accum_124__7_, prod_accum_124__6_, prod_accum_124__5_, prod_accum_124__4_, prod_accum_124__3_, prod_accum_124__2_, prod_accum_124__1_, prod_accum_124__0_ })
  );


  bsg_mul_array_row_128_125_x
  genblk1_125__genblk1_mid_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[15999:15872]),
    .b_i(b_r[15999:15872]),
    .s_i({ s_r_124__127_, s_r_124__126_, s_r_124__125_, s_r_124__124_, s_r_124__123_, s_r_124__122_, s_r_124__121_, s_r_124__120_, s_r_124__119_, s_r_124__118_, s_r_124__117_, s_r_124__116_, s_r_124__115_, s_r_124__114_, s_r_124__113_, s_r_124__112_, s_r_124__111_, s_r_124__110_, s_r_124__109_, s_r_124__108_, s_r_124__107_, s_r_124__106_, s_r_124__105_, s_r_124__104_, s_r_124__103_, s_r_124__102_, s_r_124__101_, s_r_124__100_, s_r_124__99_, s_r_124__98_, s_r_124__97_, s_r_124__96_, s_r_124__95_, s_r_124__94_, s_r_124__93_, s_r_124__92_, s_r_124__91_, s_r_124__90_, s_r_124__89_, s_r_124__88_, s_r_124__87_, s_r_124__86_, s_r_124__85_, s_r_124__84_, s_r_124__83_, s_r_124__82_, s_r_124__81_, s_r_124__80_, s_r_124__79_, s_r_124__78_, s_r_124__77_, s_r_124__76_, s_r_124__75_, s_r_124__74_, s_r_124__73_, s_r_124__72_, s_r_124__71_, s_r_124__70_, s_r_124__69_, s_r_124__68_, s_r_124__67_, s_r_124__66_, s_r_124__65_, s_r_124__64_, s_r_124__63_, s_r_124__62_, s_r_124__61_, s_r_124__60_, s_r_124__59_, s_r_124__58_, s_r_124__57_, s_r_124__56_, s_r_124__55_, s_r_124__54_, s_r_124__53_, s_r_124__52_, s_r_124__51_, s_r_124__50_, s_r_124__49_, s_r_124__48_, s_r_124__47_, s_r_124__46_, s_r_124__45_, s_r_124__44_, s_r_124__43_, s_r_124__42_, s_r_124__41_, s_r_124__40_, s_r_124__39_, s_r_124__38_, s_r_124__37_, s_r_124__36_, s_r_124__35_, s_r_124__34_, s_r_124__33_, s_r_124__32_, s_r_124__31_, s_r_124__30_, s_r_124__29_, s_r_124__28_, s_r_124__27_, s_r_124__26_, s_r_124__25_, s_r_124__24_, s_r_124__23_, s_r_124__22_, s_r_124__21_, s_r_124__20_, s_r_124__19_, s_r_124__18_, s_r_124__17_, s_r_124__16_, s_r_124__15_, s_r_124__14_, s_r_124__13_, s_r_124__12_, s_r_124__11_, s_r_124__10_, s_r_124__9_, s_r_124__8_, s_r_124__7_, s_r_124__6_, s_r_124__5_, s_r_124__4_, s_r_124__3_, s_r_124__2_, s_r_124__1_, s_r_124__0_ }),
    .c_i(c_r[124]),
    .prod_accum_i({ prod_accum_124__125_, prod_accum_124__124_, prod_accum_124__123_, prod_accum_124__122_, prod_accum_124__121_, prod_accum_124__120_, prod_accum_124__119_, prod_accum_124__118_, prod_accum_124__117_, prod_accum_124__116_, prod_accum_124__115_, prod_accum_124__114_, prod_accum_124__113_, prod_accum_124__112_, prod_accum_124__111_, prod_accum_124__110_, prod_accum_124__109_, prod_accum_124__108_, prod_accum_124__107_, prod_accum_124__106_, prod_accum_124__105_, prod_accum_124__104_, prod_accum_124__103_, prod_accum_124__102_, prod_accum_124__101_, prod_accum_124__100_, prod_accum_124__99_, prod_accum_124__98_, prod_accum_124__97_, prod_accum_124__96_, prod_accum_124__95_, prod_accum_124__94_, prod_accum_124__93_, prod_accum_124__92_, prod_accum_124__91_, prod_accum_124__90_, prod_accum_124__89_, prod_accum_124__88_, prod_accum_124__87_, prod_accum_124__86_, prod_accum_124__85_, prod_accum_124__84_, prod_accum_124__83_, prod_accum_124__82_, prod_accum_124__81_, prod_accum_124__80_, prod_accum_124__79_, prod_accum_124__78_, prod_accum_124__77_, prod_accum_124__76_, prod_accum_124__75_, prod_accum_124__74_, prod_accum_124__73_, prod_accum_124__72_, prod_accum_124__71_, prod_accum_124__70_, prod_accum_124__69_, prod_accum_124__68_, prod_accum_124__67_, prod_accum_124__66_, prod_accum_124__65_, prod_accum_124__64_, prod_accum_124__63_, prod_accum_124__62_, prod_accum_124__61_, prod_accum_124__60_, prod_accum_124__59_, prod_accum_124__58_, prod_accum_124__57_, prod_accum_124__56_, prod_accum_124__55_, prod_accum_124__54_, prod_accum_124__53_, prod_accum_124__52_, prod_accum_124__51_, prod_accum_124__50_, prod_accum_124__49_, prod_accum_124__48_, prod_accum_124__47_, prod_accum_124__46_, prod_accum_124__45_, prod_accum_124__44_, prod_accum_124__43_, prod_accum_124__42_, prod_accum_124__41_, prod_accum_124__40_, prod_accum_124__39_, prod_accum_124__38_, prod_accum_124__37_, prod_accum_124__36_, prod_accum_124__35_, prod_accum_124__34_, prod_accum_124__33_, prod_accum_124__32_, prod_accum_124__31_, prod_accum_124__30_, prod_accum_124__29_, prod_accum_124__28_, prod_accum_124__27_, prod_accum_124__26_, prod_accum_124__25_, prod_accum_124__24_, prod_accum_124__23_, prod_accum_124__22_, prod_accum_124__21_, prod_accum_124__20_, prod_accum_124__19_, prod_accum_124__18_, prod_accum_124__17_, prod_accum_124__16_, prod_accum_124__15_, prod_accum_124__14_, prod_accum_124__13_, prod_accum_124__12_, prod_accum_124__11_, prod_accum_124__10_, prod_accum_124__9_, prod_accum_124__8_, prod_accum_124__7_, prod_accum_124__6_, prod_accum_124__5_, prod_accum_124__4_, prod_accum_124__3_, prod_accum_124__2_, prod_accum_124__1_, prod_accum_124__0_ }),
    .a_o(a_r[16127:16000]),
    .b_o(b_r[16127:16000]),
    .s_o({ s_r_125__127_, s_r_125__126_, s_r_125__125_, s_r_125__124_, s_r_125__123_, s_r_125__122_, s_r_125__121_, s_r_125__120_, s_r_125__119_, s_r_125__118_, s_r_125__117_, s_r_125__116_, s_r_125__115_, s_r_125__114_, s_r_125__113_, s_r_125__112_, s_r_125__111_, s_r_125__110_, s_r_125__109_, s_r_125__108_, s_r_125__107_, s_r_125__106_, s_r_125__105_, s_r_125__104_, s_r_125__103_, s_r_125__102_, s_r_125__101_, s_r_125__100_, s_r_125__99_, s_r_125__98_, s_r_125__97_, s_r_125__96_, s_r_125__95_, s_r_125__94_, s_r_125__93_, s_r_125__92_, s_r_125__91_, s_r_125__90_, s_r_125__89_, s_r_125__88_, s_r_125__87_, s_r_125__86_, s_r_125__85_, s_r_125__84_, s_r_125__83_, s_r_125__82_, s_r_125__81_, s_r_125__80_, s_r_125__79_, s_r_125__78_, s_r_125__77_, s_r_125__76_, s_r_125__75_, s_r_125__74_, s_r_125__73_, s_r_125__72_, s_r_125__71_, s_r_125__70_, s_r_125__69_, s_r_125__68_, s_r_125__67_, s_r_125__66_, s_r_125__65_, s_r_125__64_, s_r_125__63_, s_r_125__62_, s_r_125__61_, s_r_125__60_, s_r_125__59_, s_r_125__58_, s_r_125__57_, s_r_125__56_, s_r_125__55_, s_r_125__54_, s_r_125__53_, s_r_125__52_, s_r_125__51_, s_r_125__50_, s_r_125__49_, s_r_125__48_, s_r_125__47_, s_r_125__46_, s_r_125__45_, s_r_125__44_, s_r_125__43_, s_r_125__42_, s_r_125__41_, s_r_125__40_, s_r_125__39_, s_r_125__38_, s_r_125__37_, s_r_125__36_, s_r_125__35_, s_r_125__34_, s_r_125__33_, s_r_125__32_, s_r_125__31_, s_r_125__30_, s_r_125__29_, s_r_125__28_, s_r_125__27_, s_r_125__26_, s_r_125__25_, s_r_125__24_, s_r_125__23_, s_r_125__22_, s_r_125__21_, s_r_125__20_, s_r_125__19_, s_r_125__18_, s_r_125__17_, s_r_125__16_, s_r_125__15_, s_r_125__14_, s_r_125__13_, s_r_125__12_, s_r_125__11_, s_r_125__10_, s_r_125__9_, s_r_125__8_, s_r_125__7_, s_r_125__6_, s_r_125__5_, s_r_125__4_, s_r_125__3_, s_r_125__2_, s_r_125__1_, s_r_125__0_ }),
    .c_o(c_r[125]),
    .prod_accum_o({ prod_accum_125__126_, prod_accum_125__125_, prod_accum_125__124_, prod_accum_125__123_, prod_accum_125__122_, prod_accum_125__121_, prod_accum_125__120_, prod_accum_125__119_, prod_accum_125__118_, prod_accum_125__117_, prod_accum_125__116_, prod_accum_125__115_, prod_accum_125__114_, prod_accum_125__113_, prod_accum_125__112_, prod_accum_125__111_, prod_accum_125__110_, prod_accum_125__109_, prod_accum_125__108_, prod_accum_125__107_, prod_accum_125__106_, prod_accum_125__105_, prod_accum_125__104_, prod_accum_125__103_, prod_accum_125__102_, prod_accum_125__101_, prod_accum_125__100_, prod_accum_125__99_, prod_accum_125__98_, prod_accum_125__97_, prod_accum_125__96_, prod_accum_125__95_, prod_accum_125__94_, prod_accum_125__93_, prod_accum_125__92_, prod_accum_125__91_, prod_accum_125__90_, prod_accum_125__89_, prod_accum_125__88_, prod_accum_125__87_, prod_accum_125__86_, prod_accum_125__85_, prod_accum_125__84_, prod_accum_125__83_, prod_accum_125__82_, prod_accum_125__81_, prod_accum_125__80_, prod_accum_125__79_, prod_accum_125__78_, prod_accum_125__77_, prod_accum_125__76_, prod_accum_125__75_, prod_accum_125__74_, prod_accum_125__73_, prod_accum_125__72_, prod_accum_125__71_, prod_accum_125__70_, prod_accum_125__69_, prod_accum_125__68_, prod_accum_125__67_, prod_accum_125__66_, prod_accum_125__65_, prod_accum_125__64_, prod_accum_125__63_, prod_accum_125__62_, prod_accum_125__61_, prod_accum_125__60_, prod_accum_125__59_, prod_accum_125__58_, prod_accum_125__57_, prod_accum_125__56_, prod_accum_125__55_, prod_accum_125__54_, prod_accum_125__53_, prod_accum_125__52_, prod_accum_125__51_, prod_accum_125__50_, prod_accum_125__49_, prod_accum_125__48_, prod_accum_125__47_, prod_accum_125__46_, prod_accum_125__45_, prod_accum_125__44_, prod_accum_125__43_, prod_accum_125__42_, prod_accum_125__41_, prod_accum_125__40_, prod_accum_125__39_, prod_accum_125__38_, prod_accum_125__37_, prod_accum_125__36_, prod_accum_125__35_, prod_accum_125__34_, prod_accum_125__33_, prod_accum_125__32_, prod_accum_125__31_, prod_accum_125__30_, prod_accum_125__29_, prod_accum_125__28_, prod_accum_125__27_, prod_accum_125__26_, prod_accum_125__25_, prod_accum_125__24_, prod_accum_125__23_, prod_accum_125__22_, prod_accum_125__21_, prod_accum_125__20_, prod_accum_125__19_, prod_accum_125__18_, prod_accum_125__17_, prod_accum_125__16_, prod_accum_125__15_, prod_accum_125__14_, prod_accum_125__13_, prod_accum_125__12_, prod_accum_125__11_, prod_accum_125__10_, prod_accum_125__9_, prod_accum_125__8_, prod_accum_125__7_, prod_accum_125__6_, prod_accum_125__5_, prod_accum_125__4_, prod_accum_125__3_, prod_accum_125__2_, prod_accum_125__1_, prod_accum_125__0_ })
  );


  bsg_mul_array_row_128_126_x
  genblk1_126__genblk1_last_row
  (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .v_i(v_i),
    .a_i(a_r[16127:16000]),
    .b_i(b_r[16127:16000]),
    .s_i({ s_r_125__127_, s_r_125__126_, s_r_125__125_, s_r_125__124_, s_r_125__123_, s_r_125__122_, s_r_125__121_, s_r_125__120_, s_r_125__119_, s_r_125__118_, s_r_125__117_, s_r_125__116_, s_r_125__115_, s_r_125__114_, s_r_125__113_, s_r_125__112_, s_r_125__111_, s_r_125__110_, s_r_125__109_, s_r_125__108_, s_r_125__107_, s_r_125__106_, s_r_125__105_, s_r_125__104_, s_r_125__103_, s_r_125__102_, s_r_125__101_, s_r_125__100_, s_r_125__99_, s_r_125__98_, s_r_125__97_, s_r_125__96_, s_r_125__95_, s_r_125__94_, s_r_125__93_, s_r_125__92_, s_r_125__91_, s_r_125__90_, s_r_125__89_, s_r_125__88_, s_r_125__87_, s_r_125__86_, s_r_125__85_, s_r_125__84_, s_r_125__83_, s_r_125__82_, s_r_125__81_, s_r_125__80_, s_r_125__79_, s_r_125__78_, s_r_125__77_, s_r_125__76_, s_r_125__75_, s_r_125__74_, s_r_125__73_, s_r_125__72_, s_r_125__71_, s_r_125__70_, s_r_125__69_, s_r_125__68_, s_r_125__67_, s_r_125__66_, s_r_125__65_, s_r_125__64_, s_r_125__63_, s_r_125__62_, s_r_125__61_, s_r_125__60_, s_r_125__59_, s_r_125__58_, s_r_125__57_, s_r_125__56_, s_r_125__55_, s_r_125__54_, s_r_125__53_, s_r_125__52_, s_r_125__51_, s_r_125__50_, s_r_125__49_, s_r_125__48_, s_r_125__47_, s_r_125__46_, s_r_125__45_, s_r_125__44_, s_r_125__43_, s_r_125__42_, s_r_125__41_, s_r_125__40_, s_r_125__39_, s_r_125__38_, s_r_125__37_, s_r_125__36_, s_r_125__35_, s_r_125__34_, s_r_125__33_, s_r_125__32_, s_r_125__31_, s_r_125__30_, s_r_125__29_, s_r_125__28_, s_r_125__27_, s_r_125__26_, s_r_125__25_, s_r_125__24_, s_r_125__23_, s_r_125__22_, s_r_125__21_, s_r_125__20_, s_r_125__19_, s_r_125__18_, s_r_125__17_, s_r_125__16_, s_r_125__15_, s_r_125__14_, s_r_125__13_, s_r_125__12_, s_r_125__11_, s_r_125__10_, s_r_125__9_, s_r_125__8_, s_r_125__7_, s_r_125__6_, s_r_125__5_, s_r_125__4_, s_r_125__3_, s_r_125__2_, s_r_125__1_, s_r_125__0_ }),
    .c_i(c_r[125]),
    .prod_accum_i({ prod_accum_125__126_, prod_accum_125__125_, prod_accum_125__124_, prod_accum_125__123_, prod_accum_125__122_, prod_accum_125__121_, prod_accum_125__120_, prod_accum_125__119_, prod_accum_125__118_, prod_accum_125__117_, prod_accum_125__116_, prod_accum_125__115_, prod_accum_125__114_, prod_accum_125__113_, prod_accum_125__112_, prod_accum_125__111_, prod_accum_125__110_, prod_accum_125__109_, prod_accum_125__108_, prod_accum_125__107_, prod_accum_125__106_, prod_accum_125__105_, prod_accum_125__104_, prod_accum_125__103_, prod_accum_125__102_, prod_accum_125__101_, prod_accum_125__100_, prod_accum_125__99_, prod_accum_125__98_, prod_accum_125__97_, prod_accum_125__96_, prod_accum_125__95_, prod_accum_125__94_, prod_accum_125__93_, prod_accum_125__92_, prod_accum_125__91_, prod_accum_125__90_, prod_accum_125__89_, prod_accum_125__88_, prod_accum_125__87_, prod_accum_125__86_, prod_accum_125__85_, prod_accum_125__84_, prod_accum_125__83_, prod_accum_125__82_, prod_accum_125__81_, prod_accum_125__80_, prod_accum_125__79_, prod_accum_125__78_, prod_accum_125__77_, prod_accum_125__76_, prod_accum_125__75_, prod_accum_125__74_, prod_accum_125__73_, prod_accum_125__72_, prod_accum_125__71_, prod_accum_125__70_, prod_accum_125__69_, prod_accum_125__68_, prod_accum_125__67_, prod_accum_125__66_, prod_accum_125__65_, prod_accum_125__64_, prod_accum_125__63_, prod_accum_125__62_, prod_accum_125__61_, prod_accum_125__60_, prod_accum_125__59_, prod_accum_125__58_, prod_accum_125__57_, prod_accum_125__56_, prod_accum_125__55_, prod_accum_125__54_, prod_accum_125__53_, prod_accum_125__52_, prod_accum_125__51_, prod_accum_125__50_, prod_accum_125__49_, prod_accum_125__48_, prod_accum_125__47_, prod_accum_125__46_, prod_accum_125__45_, prod_accum_125__44_, prod_accum_125__43_, prod_accum_125__42_, prod_accum_125__41_, prod_accum_125__40_, prod_accum_125__39_, prod_accum_125__38_, prod_accum_125__37_, prod_accum_125__36_, prod_accum_125__35_, prod_accum_125__34_, prod_accum_125__33_, prod_accum_125__32_, prod_accum_125__31_, prod_accum_125__30_, prod_accum_125__29_, prod_accum_125__28_, prod_accum_125__27_, prod_accum_125__26_, prod_accum_125__25_, prod_accum_125__24_, prod_accum_125__23_, prod_accum_125__22_, prod_accum_125__21_, prod_accum_125__20_, prod_accum_125__19_, prod_accum_125__18_, prod_accum_125__17_, prod_accum_125__16_, prod_accum_125__15_, prod_accum_125__14_, prod_accum_125__13_, prod_accum_125__12_, prod_accum_125__11_, prod_accum_125__10_, prod_accum_125__9_, prod_accum_125__8_, prod_accum_125__7_, prod_accum_125__6_, prod_accum_125__5_, prod_accum_125__4_, prod_accum_125__3_, prod_accum_125__2_, prod_accum_125__1_, prod_accum_125__0_ }),
    .a_o({ SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128 }),
    .b_o({ SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256 }),
    .s_o(o[254:127]),
    .c_o(o[255]),
    .prod_accum_o({ prod_accum_126__127_, o[126:0] })
  );


endmodule

