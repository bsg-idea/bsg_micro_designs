

module top
(
  i,
  o
);

  input [127:0] i;
  output [65535:0] o;

  bsg_expand_bitmask
  wrapper
  (
    .i(i),
    .o(o)
  );


endmodule



module bsg_expand_bitmask
(
  i,
  o
);

  input [127:0] i;
  output [65535:0] o;
  wire [65535:0] o;
  assign o[65024] = i[127];
  assign o[65025] = i[127];
  assign o[65026] = i[127];
  assign o[65027] = i[127];
  assign o[65028] = i[127];
  assign o[65029] = i[127];
  assign o[65030] = i[127];
  assign o[65031] = i[127];
  assign o[65032] = i[127];
  assign o[65033] = i[127];
  assign o[65034] = i[127];
  assign o[65035] = i[127];
  assign o[65036] = i[127];
  assign o[65037] = i[127];
  assign o[65038] = i[127];
  assign o[65039] = i[127];
  assign o[65040] = i[127];
  assign o[65041] = i[127];
  assign o[65042] = i[127];
  assign o[65043] = i[127];
  assign o[65044] = i[127];
  assign o[65045] = i[127];
  assign o[65046] = i[127];
  assign o[65047] = i[127];
  assign o[65048] = i[127];
  assign o[65049] = i[127];
  assign o[65050] = i[127];
  assign o[65051] = i[127];
  assign o[65052] = i[127];
  assign o[65053] = i[127];
  assign o[65054] = i[127];
  assign o[65055] = i[127];
  assign o[65056] = i[127];
  assign o[65057] = i[127];
  assign o[65058] = i[127];
  assign o[65059] = i[127];
  assign o[65060] = i[127];
  assign o[65061] = i[127];
  assign o[65062] = i[127];
  assign o[65063] = i[127];
  assign o[65064] = i[127];
  assign o[65065] = i[127];
  assign o[65066] = i[127];
  assign o[65067] = i[127];
  assign o[65068] = i[127];
  assign o[65069] = i[127];
  assign o[65070] = i[127];
  assign o[65071] = i[127];
  assign o[65072] = i[127];
  assign o[65073] = i[127];
  assign o[65074] = i[127];
  assign o[65075] = i[127];
  assign o[65076] = i[127];
  assign o[65077] = i[127];
  assign o[65078] = i[127];
  assign o[65079] = i[127];
  assign o[65080] = i[127];
  assign o[65081] = i[127];
  assign o[65082] = i[127];
  assign o[65083] = i[127];
  assign o[65084] = i[127];
  assign o[65085] = i[127];
  assign o[65086] = i[127];
  assign o[65087] = i[127];
  assign o[65088] = i[127];
  assign o[65089] = i[127];
  assign o[65090] = i[127];
  assign o[65091] = i[127];
  assign o[65092] = i[127];
  assign o[65093] = i[127];
  assign o[65094] = i[127];
  assign o[65095] = i[127];
  assign o[65096] = i[127];
  assign o[65097] = i[127];
  assign o[65098] = i[127];
  assign o[65099] = i[127];
  assign o[65100] = i[127];
  assign o[65101] = i[127];
  assign o[65102] = i[127];
  assign o[65103] = i[127];
  assign o[65104] = i[127];
  assign o[65105] = i[127];
  assign o[65106] = i[127];
  assign o[65107] = i[127];
  assign o[65108] = i[127];
  assign o[65109] = i[127];
  assign o[65110] = i[127];
  assign o[65111] = i[127];
  assign o[65112] = i[127];
  assign o[65113] = i[127];
  assign o[65114] = i[127];
  assign o[65115] = i[127];
  assign o[65116] = i[127];
  assign o[65117] = i[127];
  assign o[65118] = i[127];
  assign o[65119] = i[127];
  assign o[65120] = i[127];
  assign o[65121] = i[127];
  assign o[65122] = i[127];
  assign o[65123] = i[127];
  assign o[65124] = i[127];
  assign o[65125] = i[127];
  assign o[65126] = i[127];
  assign o[65127] = i[127];
  assign o[65128] = i[127];
  assign o[65129] = i[127];
  assign o[65130] = i[127];
  assign o[65131] = i[127];
  assign o[65132] = i[127];
  assign o[65133] = i[127];
  assign o[65134] = i[127];
  assign o[65135] = i[127];
  assign o[65136] = i[127];
  assign o[65137] = i[127];
  assign o[65138] = i[127];
  assign o[65139] = i[127];
  assign o[65140] = i[127];
  assign o[65141] = i[127];
  assign o[65142] = i[127];
  assign o[65143] = i[127];
  assign o[65144] = i[127];
  assign o[65145] = i[127];
  assign o[65146] = i[127];
  assign o[65147] = i[127];
  assign o[65148] = i[127];
  assign o[65149] = i[127];
  assign o[65150] = i[127];
  assign o[65151] = i[127];
  assign o[65152] = i[127];
  assign o[65153] = i[127];
  assign o[65154] = i[127];
  assign o[65155] = i[127];
  assign o[65156] = i[127];
  assign o[65157] = i[127];
  assign o[65158] = i[127];
  assign o[65159] = i[127];
  assign o[65160] = i[127];
  assign o[65161] = i[127];
  assign o[65162] = i[127];
  assign o[65163] = i[127];
  assign o[65164] = i[127];
  assign o[65165] = i[127];
  assign o[65166] = i[127];
  assign o[65167] = i[127];
  assign o[65168] = i[127];
  assign o[65169] = i[127];
  assign o[65170] = i[127];
  assign o[65171] = i[127];
  assign o[65172] = i[127];
  assign o[65173] = i[127];
  assign o[65174] = i[127];
  assign o[65175] = i[127];
  assign o[65176] = i[127];
  assign o[65177] = i[127];
  assign o[65178] = i[127];
  assign o[65179] = i[127];
  assign o[65180] = i[127];
  assign o[65181] = i[127];
  assign o[65182] = i[127];
  assign o[65183] = i[127];
  assign o[65184] = i[127];
  assign o[65185] = i[127];
  assign o[65186] = i[127];
  assign o[65187] = i[127];
  assign o[65188] = i[127];
  assign o[65189] = i[127];
  assign o[65190] = i[127];
  assign o[65191] = i[127];
  assign o[65192] = i[127];
  assign o[65193] = i[127];
  assign o[65194] = i[127];
  assign o[65195] = i[127];
  assign o[65196] = i[127];
  assign o[65197] = i[127];
  assign o[65198] = i[127];
  assign o[65199] = i[127];
  assign o[65200] = i[127];
  assign o[65201] = i[127];
  assign o[65202] = i[127];
  assign o[65203] = i[127];
  assign o[65204] = i[127];
  assign o[65205] = i[127];
  assign o[65206] = i[127];
  assign o[65207] = i[127];
  assign o[65208] = i[127];
  assign o[65209] = i[127];
  assign o[65210] = i[127];
  assign o[65211] = i[127];
  assign o[65212] = i[127];
  assign o[65213] = i[127];
  assign o[65214] = i[127];
  assign o[65215] = i[127];
  assign o[65216] = i[127];
  assign o[65217] = i[127];
  assign o[65218] = i[127];
  assign o[65219] = i[127];
  assign o[65220] = i[127];
  assign o[65221] = i[127];
  assign o[65222] = i[127];
  assign o[65223] = i[127];
  assign o[65224] = i[127];
  assign o[65225] = i[127];
  assign o[65226] = i[127];
  assign o[65227] = i[127];
  assign o[65228] = i[127];
  assign o[65229] = i[127];
  assign o[65230] = i[127];
  assign o[65231] = i[127];
  assign o[65232] = i[127];
  assign o[65233] = i[127];
  assign o[65234] = i[127];
  assign o[65235] = i[127];
  assign o[65236] = i[127];
  assign o[65237] = i[127];
  assign o[65238] = i[127];
  assign o[65239] = i[127];
  assign o[65240] = i[127];
  assign o[65241] = i[127];
  assign o[65242] = i[127];
  assign o[65243] = i[127];
  assign o[65244] = i[127];
  assign o[65245] = i[127];
  assign o[65246] = i[127];
  assign o[65247] = i[127];
  assign o[65248] = i[127];
  assign o[65249] = i[127];
  assign o[65250] = i[127];
  assign o[65251] = i[127];
  assign o[65252] = i[127];
  assign o[65253] = i[127];
  assign o[65254] = i[127];
  assign o[65255] = i[127];
  assign o[65256] = i[127];
  assign o[65257] = i[127];
  assign o[65258] = i[127];
  assign o[65259] = i[127];
  assign o[65260] = i[127];
  assign o[65261] = i[127];
  assign o[65262] = i[127];
  assign o[65263] = i[127];
  assign o[65264] = i[127];
  assign o[65265] = i[127];
  assign o[65266] = i[127];
  assign o[65267] = i[127];
  assign o[65268] = i[127];
  assign o[65269] = i[127];
  assign o[65270] = i[127];
  assign o[65271] = i[127];
  assign o[65272] = i[127];
  assign o[65273] = i[127];
  assign o[65274] = i[127];
  assign o[65275] = i[127];
  assign o[65276] = i[127];
  assign o[65277] = i[127];
  assign o[65278] = i[127];
  assign o[65279] = i[127];
  assign o[65280] = i[127];
  assign o[65281] = i[127];
  assign o[65282] = i[127];
  assign o[65283] = i[127];
  assign o[65284] = i[127];
  assign o[65285] = i[127];
  assign o[65286] = i[127];
  assign o[65287] = i[127];
  assign o[65288] = i[127];
  assign o[65289] = i[127];
  assign o[65290] = i[127];
  assign o[65291] = i[127];
  assign o[65292] = i[127];
  assign o[65293] = i[127];
  assign o[65294] = i[127];
  assign o[65295] = i[127];
  assign o[65296] = i[127];
  assign o[65297] = i[127];
  assign o[65298] = i[127];
  assign o[65299] = i[127];
  assign o[65300] = i[127];
  assign o[65301] = i[127];
  assign o[65302] = i[127];
  assign o[65303] = i[127];
  assign o[65304] = i[127];
  assign o[65305] = i[127];
  assign o[65306] = i[127];
  assign o[65307] = i[127];
  assign o[65308] = i[127];
  assign o[65309] = i[127];
  assign o[65310] = i[127];
  assign o[65311] = i[127];
  assign o[65312] = i[127];
  assign o[65313] = i[127];
  assign o[65314] = i[127];
  assign o[65315] = i[127];
  assign o[65316] = i[127];
  assign o[65317] = i[127];
  assign o[65318] = i[127];
  assign o[65319] = i[127];
  assign o[65320] = i[127];
  assign o[65321] = i[127];
  assign o[65322] = i[127];
  assign o[65323] = i[127];
  assign o[65324] = i[127];
  assign o[65325] = i[127];
  assign o[65326] = i[127];
  assign o[65327] = i[127];
  assign o[65328] = i[127];
  assign o[65329] = i[127];
  assign o[65330] = i[127];
  assign o[65331] = i[127];
  assign o[65332] = i[127];
  assign o[65333] = i[127];
  assign o[65334] = i[127];
  assign o[65335] = i[127];
  assign o[65336] = i[127];
  assign o[65337] = i[127];
  assign o[65338] = i[127];
  assign o[65339] = i[127];
  assign o[65340] = i[127];
  assign o[65341] = i[127];
  assign o[65342] = i[127];
  assign o[65343] = i[127];
  assign o[65344] = i[127];
  assign o[65345] = i[127];
  assign o[65346] = i[127];
  assign o[65347] = i[127];
  assign o[65348] = i[127];
  assign o[65349] = i[127];
  assign o[65350] = i[127];
  assign o[65351] = i[127];
  assign o[65352] = i[127];
  assign o[65353] = i[127];
  assign o[65354] = i[127];
  assign o[65355] = i[127];
  assign o[65356] = i[127];
  assign o[65357] = i[127];
  assign o[65358] = i[127];
  assign o[65359] = i[127];
  assign o[65360] = i[127];
  assign o[65361] = i[127];
  assign o[65362] = i[127];
  assign o[65363] = i[127];
  assign o[65364] = i[127];
  assign o[65365] = i[127];
  assign o[65366] = i[127];
  assign o[65367] = i[127];
  assign o[65368] = i[127];
  assign o[65369] = i[127];
  assign o[65370] = i[127];
  assign o[65371] = i[127];
  assign o[65372] = i[127];
  assign o[65373] = i[127];
  assign o[65374] = i[127];
  assign o[65375] = i[127];
  assign o[65376] = i[127];
  assign o[65377] = i[127];
  assign o[65378] = i[127];
  assign o[65379] = i[127];
  assign o[65380] = i[127];
  assign o[65381] = i[127];
  assign o[65382] = i[127];
  assign o[65383] = i[127];
  assign o[65384] = i[127];
  assign o[65385] = i[127];
  assign o[65386] = i[127];
  assign o[65387] = i[127];
  assign o[65388] = i[127];
  assign o[65389] = i[127];
  assign o[65390] = i[127];
  assign o[65391] = i[127];
  assign o[65392] = i[127];
  assign o[65393] = i[127];
  assign o[65394] = i[127];
  assign o[65395] = i[127];
  assign o[65396] = i[127];
  assign o[65397] = i[127];
  assign o[65398] = i[127];
  assign o[65399] = i[127];
  assign o[65400] = i[127];
  assign o[65401] = i[127];
  assign o[65402] = i[127];
  assign o[65403] = i[127];
  assign o[65404] = i[127];
  assign o[65405] = i[127];
  assign o[65406] = i[127];
  assign o[65407] = i[127];
  assign o[65408] = i[127];
  assign o[65409] = i[127];
  assign o[65410] = i[127];
  assign o[65411] = i[127];
  assign o[65412] = i[127];
  assign o[65413] = i[127];
  assign o[65414] = i[127];
  assign o[65415] = i[127];
  assign o[65416] = i[127];
  assign o[65417] = i[127];
  assign o[65418] = i[127];
  assign o[65419] = i[127];
  assign o[65420] = i[127];
  assign o[65421] = i[127];
  assign o[65422] = i[127];
  assign o[65423] = i[127];
  assign o[65424] = i[127];
  assign o[65425] = i[127];
  assign o[65426] = i[127];
  assign o[65427] = i[127];
  assign o[65428] = i[127];
  assign o[65429] = i[127];
  assign o[65430] = i[127];
  assign o[65431] = i[127];
  assign o[65432] = i[127];
  assign o[65433] = i[127];
  assign o[65434] = i[127];
  assign o[65435] = i[127];
  assign o[65436] = i[127];
  assign o[65437] = i[127];
  assign o[65438] = i[127];
  assign o[65439] = i[127];
  assign o[65440] = i[127];
  assign o[65441] = i[127];
  assign o[65442] = i[127];
  assign o[65443] = i[127];
  assign o[65444] = i[127];
  assign o[65445] = i[127];
  assign o[65446] = i[127];
  assign o[65447] = i[127];
  assign o[65448] = i[127];
  assign o[65449] = i[127];
  assign o[65450] = i[127];
  assign o[65451] = i[127];
  assign o[65452] = i[127];
  assign o[65453] = i[127];
  assign o[65454] = i[127];
  assign o[65455] = i[127];
  assign o[65456] = i[127];
  assign o[65457] = i[127];
  assign o[65458] = i[127];
  assign o[65459] = i[127];
  assign o[65460] = i[127];
  assign o[65461] = i[127];
  assign o[65462] = i[127];
  assign o[65463] = i[127];
  assign o[65464] = i[127];
  assign o[65465] = i[127];
  assign o[65466] = i[127];
  assign o[65467] = i[127];
  assign o[65468] = i[127];
  assign o[65469] = i[127];
  assign o[65470] = i[127];
  assign o[65471] = i[127];
  assign o[65472] = i[127];
  assign o[65473] = i[127];
  assign o[65474] = i[127];
  assign o[65475] = i[127];
  assign o[65476] = i[127];
  assign o[65477] = i[127];
  assign o[65478] = i[127];
  assign o[65479] = i[127];
  assign o[65480] = i[127];
  assign o[65481] = i[127];
  assign o[65482] = i[127];
  assign o[65483] = i[127];
  assign o[65484] = i[127];
  assign o[65485] = i[127];
  assign o[65486] = i[127];
  assign o[65487] = i[127];
  assign o[65488] = i[127];
  assign o[65489] = i[127];
  assign o[65490] = i[127];
  assign o[65491] = i[127];
  assign o[65492] = i[127];
  assign o[65493] = i[127];
  assign o[65494] = i[127];
  assign o[65495] = i[127];
  assign o[65496] = i[127];
  assign o[65497] = i[127];
  assign o[65498] = i[127];
  assign o[65499] = i[127];
  assign o[65500] = i[127];
  assign o[65501] = i[127];
  assign o[65502] = i[127];
  assign o[65503] = i[127];
  assign o[65504] = i[127];
  assign o[65505] = i[127];
  assign o[65506] = i[127];
  assign o[65507] = i[127];
  assign o[65508] = i[127];
  assign o[65509] = i[127];
  assign o[65510] = i[127];
  assign o[65511] = i[127];
  assign o[65512] = i[127];
  assign o[65513] = i[127];
  assign o[65514] = i[127];
  assign o[65515] = i[127];
  assign o[65516] = i[127];
  assign o[65517] = i[127];
  assign o[65518] = i[127];
  assign o[65519] = i[127];
  assign o[65520] = i[127];
  assign o[65521] = i[127];
  assign o[65522] = i[127];
  assign o[65523] = i[127];
  assign o[65524] = i[127];
  assign o[65525] = i[127];
  assign o[65526] = i[127];
  assign o[65527] = i[127];
  assign o[65528] = i[127];
  assign o[65529] = i[127];
  assign o[65530] = i[127];
  assign o[65531] = i[127];
  assign o[65532] = i[127];
  assign o[65533] = i[127];
  assign o[65534] = i[127];
  assign o[65535] = i[127];
  assign o[64512] = i[126];
  assign o[64513] = i[126];
  assign o[64514] = i[126];
  assign o[64515] = i[126];
  assign o[64516] = i[126];
  assign o[64517] = i[126];
  assign o[64518] = i[126];
  assign o[64519] = i[126];
  assign o[64520] = i[126];
  assign o[64521] = i[126];
  assign o[64522] = i[126];
  assign o[64523] = i[126];
  assign o[64524] = i[126];
  assign o[64525] = i[126];
  assign o[64526] = i[126];
  assign o[64527] = i[126];
  assign o[64528] = i[126];
  assign o[64529] = i[126];
  assign o[64530] = i[126];
  assign o[64531] = i[126];
  assign o[64532] = i[126];
  assign o[64533] = i[126];
  assign o[64534] = i[126];
  assign o[64535] = i[126];
  assign o[64536] = i[126];
  assign o[64537] = i[126];
  assign o[64538] = i[126];
  assign o[64539] = i[126];
  assign o[64540] = i[126];
  assign o[64541] = i[126];
  assign o[64542] = i[126];
  assign o[64543] = i[126];
  assign o[64544] = i[126];
  assign o[64545] = i[126];
  assign o[64546] = i[126];
  assign o[64547] = i[126];
  assign o[64548] = i[126];
  assign o[64549] = i[126];
  assign o[64550] = i[126];
  assign o[64551] = i[126];
  assign o[64552] = i[126];
  assign o[64553] = i[126];
  assign o[64554] = i[126];
  assign o[64555] = i[126];
  assign o[64556] = i[126];
  assign o[64557] = i[126];
  assign o[64558] = i[126];
  assign o[64559] = i[126];
  assign o[64560] = i[126];
  assign o[64561] = i[126];
  assign o[64562] = i[126];
  assign o[64563] = i[126];
  assign o[64564] = i[126];
  assign o[64565] = i[126];
  assign o[64566] = i[126];
  assign o[64567] = i[126];
  assign o[64568] = i[126];
  assign o[64569] = i[126];
  assign o[64570] = i[126];
  assign o[64571] = i[126];
  assign o[64572] = i[126];
  assign o[64573] = i[126];
  assign o[64574] = i[126];
  assign o[64575] = i[126];
  assign o[64576] = i[126];
  assign o[64577] = i[126];
  assign o[64578] = i[126];
  assign o[64579] = i[126];
  assign o[64580] = i[126];
  assign o[64581] = i[126];
  assign o[64582] = i[126];
  assign o[64583] = i[126];
  assign o[64584] = i[126];
  assign o[64585] = i[126];
  assign o[64586] = i[126];
  assign o[64587] = i[126];
  assign o[64588] = i[126];
  assign o[64589] = i[126];
  assign o[64590] = i[126];
  assign o[64591] = i[126];
  assign o[64592] = i[126];
  assign o[64593] = i[126];
  assign o[64594] = i[126];
  assign o[64595] = i[126];
  assign o[64596] = i[126];
  assign o[64597] = i[126];
  assign o[64598] = i[126];
  assign o[64599] = i[126];
  assign o[64600] = i[126];
  assign o[64601] = i[126];
  assign o[64602] = i[126];
  assign o[64603] = i[126];
  assign o[64604] = i[126];
  assign o[64605] = i[126];
  assign o[64606] = i[126];
  assign o[64607] = i[126];
  assign o[64608] = i[126];
  assign o[64609] = i[126];
  assign o[64610] = i[126];
  assign o[64611] = i[126];
  assign o[64612] = i[126];
  assign o[64613] = i[126];
  assign o[64614] = i[126];
  assign o[64615] = i[126];
  assign o[64616] = i[126];
  assign o[64617] = i[126];
  assign o[64618] = i[126];
  assign o[64619] = i[126];
  assign o[64620] = i[126];
  assign o[64621] = i[126];
  assign o[64622] = i[126];
  assign o[64623] = i[126];
  assign o[64624] = i[126];
  assign o[64625] = i[126];
  assign o[64626] = i[126];
  assign o[64627] = i[126];
  assign o[64628] = i[126];
  assign o[64629] = i[126];
  assign o[64630] = i[126];
  assign o[64631] = i[126];
  assign o[64632] = i[126];
  assign o[64633] = i[126];
  assign o[64634] = i[126];
  assign o[64635] = i[126];
  assign o[64636] = i[126];
  assign o[64637] = i[126];
  assign o[64638] = i[126];
  assign o[64639] = i[126];
  assign o[64640] = i[126];
  assign o[64641] = i[126];
  assign o[64642] = i[126];
  assign o[64643] = i[126];
  assign o[64644] = i[126];
  assign o[64645] = i[126];
  assign o[64646] = i[126];
  assign o[64647] = i[126];
  assign o[64648] = i[126];
  assign o[64649] = i[126];
  assign o[64650] = i[126];
  assign o[64651] = i[126];
  assign o[64652] = i[126];
  assign o[64653] = i[126];
  assign o[64654] = i[126];
  assign o[64655] = i[126];
  assign o[64656] = i[126];
  assign o[64657] = i[126];
  assign o[64658] = i[126];
  assign o[64659] = i[126];
  assign o[64660] = i[126];
  assign o[64661] = i[126];
  assign o[64662] = i[126];
  assign o[64663] = i[126];
  assign o[64664] = i[126];
  assign o[64665] = i[126];
  assign o[64666] = i[126];
  assign o[64667] = i[126];
  assign o[64668] = i[126];
  assign o[64669] = i[126];
  assign o[64670] = i[126];
  assign o[64671] = i[126];
  assign o[64672] = i[126];
  assign o[64673] = i[126];
  assign o[64674] = i[126];
  assign o[64675] = i[126];
  assign o[64676] = i[126];
  assign o[64677] = i[126];
  assign o[64678] = i[126];
  assign o[64679] = i[126];
  assign o[64680] = i[126];
  assign o[64681] = i[126];
  assign o[64682] = i[126];
  assign o[64683] = i[126];
  assign o[64684] = i[126];
  assign o[64685] = i[126];
  assign o[64686] = i[126];
  assign o[64687] = i[126];
  assign o[64688] = i[126];
  assign o[64689] = i[126];
  assign o[64690] = i[126];
  assign o[64691] = i[126];
  assign o[64692] = i[126];
  assign o[64693] = i[126];
  assign o[64694] = i[126];
  assign o[64695] = i[126];
  assign o[64696] = i[126];
  assign o[64697] = i[126];
  assign o[64698] = i[126];
  assign o[64699] = i[126];
  assign o[64700] = i[126];
  assign o[64701] = i[126];
  assign o[64702] = i[126];
  assign o[64703] = i[126];
  assign o[64704] = i[126];
  assign o[64705] = i[126];
  assign o[64706] = i[126];
  assign o[64707] = i[126];
  assign o[64708] = i[126];
  assign o[64709] = i[126];
  assign o[64710] = i[126];
  assign o[64711] = i[126];
  assign o[64712] = i[126];
  assign o[64713] = i[126];
  assign o[64714] = i[126];
  assign o[64715] = i[126];
  assign o[64716] = i[126];
  assign o[64717] = i[126];
  assign o[64718] = i[126];
  assign o[64719] = i[126];
  assign o[64720] = i[126];
  assign o[64721] = i[126];
  assign o[64722] = i[126];
  assign o[64723] = i[126];
  assign o[64724] = i[126];
  assign o[64725] = i[126];
  assign o[64726] = i[126];
  assign o[64727] = i[126];
  assign o[64728] = i[126];
  assign o[64729] = i[126];
  assign o[64730] = i[126];
  assign o[64731] = i[126];
  assign o[64732] = i[126];
  assign o[64733] = i[126];
  assign o[64734] = i[126];
  assign o[64735] = i[126];
  assign o[64736] = i[126];
  assign o[64737] = i[126];
  assign o[64738] = i[126];
  assign o[64739] = i[126];
  assign o[64740] = i[126];
  assign o[64741] = i[126];
  assign o[64742] = i[126];
  assign o[64743] = i[126];
  assign o[64744] = i[126];
  assign o[64745] = i[126];
  assign o[64746] = i[126];
  assign o[64747] = i[126];
  assign o[64748] = i[126];
  assign o[64749] = i[126];
  assign o[64750] = i[126];
  assign o[64751] = i[126];
  assign o[64752] = i[126];
  assign o[64753] = i[126];
  assign o[64754] = i[126];
  assign o[64755] = i[126];
  assign o[64756] = i[126];
  assign o[64757] = i[126];
  assign o[64758] = i[126];
  assign o[64759] = i[126];
  assign o[64760] = i[126];
  assign o[64761] = i[126];
  assign o[64762] = i[126];
  assign o[64763] = i[126];
  assign o[64764] = i[126];
  assign o[64765] = i[126];
  assign o[64766] = i[126];
  assign o[64767] = i[126];
  assign o[64768] = i[126];
  assign o[64769] = i[126];
  assign o[64770] = i[126];
  assign o[64771] = i[126];
  assign o[64772] = i[126];
  assign o[64773] = i[126];
  assign o[64774] = i[126];
  assign o[64775] = i[126];
  assign o[64776] = i[126];
  assign o[64777] = i[126];
  assign o[64778] = i[126];
  assign o[64779] = i[126];
  assign o[64780] = i[126];
  assign o[64781] = i[126];
  assign o[64782] = i[126];
  assign o[64783] = i[126];
  assign o[64784] = i[126];
  assign o[64785] = i[126];
  assign o[64786] = i[126];
  assign o[64787] = i[126];
  assign o[64788] = i[126];
  assign o[64789] = i[126];
  assign o[64790] = i[126];
  assign o[64791] = i[126];
  assign o[64792] = i[126];
  assign o[64793] = i[126];
  assign o[64794] = i[126];
  assign o[64795] = i[126];
  assign o[64796] = i[126];
  assign o[64797] = i[126];
  assign o[64798] = i[126];
  assign o[64799] = i[126];
  assign o[64800] = i[126];
  assign o[64801] = i[126];
  assign o[64802] = i[126];
  assign o[64803] = i[126];
  assign o[64804] = i[126];
  assign o[64805] = i[126];
  assign o[64806] = i[126];
  assign o[64807] = i[126];
  assign o[64808] = i[126];
  assign o[64809] = i[126];
  assign o[64810] = i[126];
  assign o[64811] = i[126];
  assign o[64812] = i[126];
  assign o[64813] = i[126];
  assign o[64814] = i[126];
  assign o[64815] = i[126];
  assign o[64816] = i[126];
  assign o[64817] = i[126];
  assign o[64818] = i[126];
  assign o[64819] = i[126];
  assign o[64820] = i[126];
  assign o[64821] = i[126];
  assign o[64822] = i[126];
  assign o[64823] = i[126];
  assign o[64824] = i[126];
  assign o[64825] = i[126];
  assign o[64826] = i[126];
  assign o[64827] = i[126];
  assign o[64828] = i[126];
  assign o[64829] = i[126];
  assign o[64830] = i[126];
  assign o[64831] = i[126];
  assign o[64832] = i[126];
  assign o[64833] = i[126];
  assign o[64834] = i[126];
  assign o[64835] = i[126];
  assign o[64836] = i[126];
  assign o[64837] = i[126];
  assign o[64838] = i[126];
  assign o[64839] = i[126];
  assign o[64840] = i[126];
  assign o[64841] = i[126];
  assign o[64842] = i[126];
  assign o[64843] = i[126];
  assign o[64844] = i[126];
  assign o[64845] = i[126];
  assign o[64846] = i[126];
  assign o[64847] = i[126];
  assign o[64848] = i[126];
  assign o[64849] = i[126];
  assign o[64850] = i[126];
  assign o[64851] = i[126];
  assign o[64852] = i[126];
  assign o[64853] = i[126];
  assign o[64854] = i[126];
  assign o[64855] = i[126];
  assign o[64856] = i[126];
  assign o[64857] = i[126];
  assign o[64858] = i[126];
  assign o[64859] = i[126];
  assign o[64860] = i[126];
  assign o[64861] = i[126];
  assign o[64862] = i[126];
  assign o[64863] = i[126];
  assign o[64864] = i[126];
  assign o[64865] = i[126];
  assign o[64866] = i[126];
  assign o[64867] = i[126];
  assign o[64868] = i[126];
  assign o[64869] = i[126];
  assign o[64870] = i[126];
  assign o[64871] = i[126];
  assign o[64872] = i[126];
  assign o[64873] = i[126];
  assign o[64874] = i[126];
  assign o[64875] = i[126];
  assign o[64876] = i[126];
  assign o[64877] = i[126];
  assign o[64878] = i[126];
  assign o[64879] = i[126];
  assign o[64880] = i[126];
  assign o[64881] = i[126];
  assign o[64882] = i[126];
  assign o[64883] = i[126];
  assign o[64884] = i[126];
  assign o[64885] = i[126];
  assign o[64886] = i[126];
  assign o[64887] = i[126];
  assign o[64888] = i[126];
  assign o[64889] = i[126];
  assign o[64890] = i[126];
  assign o[64891] = i[126];
  assign o[64892] = i[126];
  assign o[64893] = i[126];
  assign o[64894] = i[126];
  assign o[64895] = i[126];
  assign o[64896] = i[126];
  assign o[64897] = i[126];
  assign o[64898] = i[126];
  assign o[64899] = i[126];
  assign o[64900] = i[126];
  assign o[64901] = i[126];
  assign o[64902] = i[126];
  assign o[64903] = i[126];
  assign o[64904] = i[126];
  assign o[64905] = i[126];
  assign o[64906] = i[126];
  assign o[64907] = i[126];
  assign o[64908] = i[126];
  assign o[64909] = i[126];
  assign o[64910] = i[126];
  assign o[64911] = i[126];
  assign o[64912] = i[126];
  assign o[64913] = i[126];
  assign o[64914] = i[126];
  assign o[64915] = i[126];
  assign o[64916] = i[126];
  assign o[64917] = i[126];
  assign o[64918] = i[126];
  assign o[64919] = i[126];
  assign o[64920] = i[126];
  assign o[64921] = i[126];
  assign o[64922] = i[126];
  assign o[64923] = i[126];
  assign o[64924] = i[126];
  assign o[64925] = i[126];
  assign o[64926] = i[126];
  assign o[64927] = i[126];
  assign o[64928] = i[126];
  assign o[64929] = i[126];
  assign o[64930] = i[126];
  assign o[64931] = i[126];
  assign o[64932] = i[126];
  assign o[64933] = i[126];
  assign o[64934] = i[126];
  assign o[64935] = i[126];
  assign o[64936] = i[126];
  assign o[64937] = i[126];
  assign o[64938] = i[126];
  assign o[64939] = i[126];
  assign o[64940] = i[126];
  assign o[64941] = i[126];
  assign o[64942] = i[126];
  assign o[64943] = i[126];
  assign o[64944] = i[126];
  assign o[64945] = i[126];
  assign o[64946] = i[126];
  assign o[64947] = i[126];
  assign o[64948] = i[126];
  assign o[64949] = i[126];
  assign o[64950] = i[126];
  assign o[64951] = i[126];
  assign o[64952] = i[126];
  assign o[64953] = i[126];
  assign o[64954] = i[126];
  assign o[64955] = i[126];
  assign o[64956] = i[126];
  assign o[64957] = i[126];
  assign o[64958] = i[126];
  assign o[64959] = i[126];
  assign o[64960] = i[126];
  assign o[64961] = i[126];
  assign o[64962] = i[126];
  assign o[64963] = i[126];
  assign o[64964] = i[126];
  assign o[64965] = i[126];
  assign o[64966] = i[126];
  assign o[64967] = i[126];
  assign o[64968] = i[126];
  assign o[64969] = i[126];
  assign o[64970] = i[126];
  assign o[64971] = i[126];
  assign o[64972] = i[126];
  assign o[64973] = i[126];
  assign o[64974] = i[126];
  assign o[64975] = i[126];
  assign o[64976] = i[126];
  assign o[64977] = i[126];
  assign o[64978] = i[126];
  assign o[64979] = i[126];
  assign o[64980] = i[126];
  assign o[64981] = i[126];
  assign o[64982] = i[126];
  assign o[64983] = i[126];
  assign o[64984] = i[126];
  assign o[64985] = i[126];
  assign o[64986] = i[126];
  assign o[64987] = i[126];
  assign o[64988] = i[126];
  assign o[64989] = i[126];
  assign o[64990] = i[126];
  assign o[64991] = i[126];
  assign o[64992] = i[126];
  assign o[64993] = i[126];
  assign o[64994] = i[126];
  assign o[64995] = i[126];
  assign o[64996] = i[126];
  assign o[64997] = i[126];
  assign o[64998] = i[126];
  assign o[64999] = i[126];
  assign o[65000] = i[126];
  assign o[65001] = i[126];
  assign o[65002] = i[126];
  assign o[65003] = i[126];
  assign o[65004] = i[126];
  assign o[65005] = i[126];
  assign o[65006] = i[126];
  assign o[65007] = i[126];
  assign o[65008] = i[126];
  assign o[65009] = i[126];
  assign o[65010] = i[126];
  assign o[65011] = i[126];
  assign o[65012] = i[126];
  assign o[65013] = i[126];
  assign o[65014] = i[126];
  assign o[65015] = i[126];
  assign o[65016] = i[126];
  assign o[65017] = i[126];
  assign o[65018] = i[126];
  assign o[65019] = i[126];
  assign o[65020] = i[126];
  assign o[65021] = i[126];
  assign o[65022] = i[126];
  assign o[65023] = i[126];
  assign o[64000] = i[125];
  assign o[64001] = i[125];
  assign o[64002] = i[125];
  assign o[64003] = i[125];
  assign o[64004] = i[125];
  assign o[64005] = i[125];
  assign o[64006] = i[125];
  assign o[64007] = i[125];
  assign o[64008] = i[125];
  assign o[64009] = i[125];
  assign o[64010] = i[125];
  assign o[64011] = i[125];
  assign o[64012] = i[125];
  assign o[64013] = i[125];
  assign o[64014] = i[125];
  assign o[64015] = i[125];
  assign o[64016] = i[125];
  assign o[64017] = i[125];
  assign o[64018] = i[125];
  assign o[64019] = i[125];
  assign o[64020] = i[125];
  assign o[64021] = i[125];
  assign o[64022] = i[125];
  assign o[64023] = i[125];
  assign o[64024] = i[125];
  assign o[64025] = i[125];
  assign o[64026] = i[125];
  assign o[64027] = i[125];
  assign o[64028] = i[125];
  assign o[64029] = i[125];
  assign o[64030] = i[125];
  assign o[64031] = i[125];
  assign o[64032] = i[125];
  assign o[64033] = i[125];
  assign o[64034] = i[125];
  assign o[64035] = i[125];
  assign o[64036] = i[125];
  assign o[64037] = i[125];
  assign o[64038] = i[125];
  assign o[64039] = i[125];
  assign o[64040] = i[125];
  assign o[64041] = i[125];
  assign o[64042] = i[125];
  assign o[64043] = i[125];
  assign o[64044] = i[125];
  assign o[64045] = i[125];
  assign o[64046] = i[125];
  assign o[64047] = i[125];
  assign o[64048] = i[125];
  assign o[64049] = i[125];
  assign o[64050] = i[125];
  assign o[64051] = i[125];
  assign o[64052] = i[125];
  assign o[64053] = i[125];
  assign o[64054] = i[125];
  assign o[64055] = i[125];
  assign o[64056] = i[125];
  assign o[64057] = i[125];
  assign o[64058] = i[125];
  assign o[64059] = i[125];
  assign o[64060] = i[125];
  assign o[64061] = i[125];
  assign o[64062] = i[125];
  assign o[64063] = i[125];
  assign o[64064] = i[125];
  assign o[64065] = i[125];
  assign o[64066] = i[125];
  assign o[64067] = i[125];
  assign o[64068] = i[125];
  assign o[64069] = i[125];
  assign o[64070] = i[125];
  assign o[64071] = i[125];
  assign o[64072] = i[125];
  assign o[64073] = i[125];
  assign o[64074] = i[125];
  assign o[64075] = i[125];
  assign o[64076] = i[125];
  assign o[64077] = i[125];
  assign o[64078] = i[125];
  assign o[64079] = i[125];
  assign o[64080] = i[125];
  assign o[64081] = i[125];
  assign o[64082] = i[125];
  assign o[64083] = i[125];
  assign o[64084] = i[125];
  assign o[64085] = i[125];
  assign o[64086] = i[125];
  assign o[64087] = i[125];
  assign o[64088] = i[125];
  assign o[64089] = i[125];
  assign o[64090] = i[125];
  assign o[64091] = i[125];
  assign o[64092] = i[125];
  assign o[64093] = i[125];
  assign o[64094] = i[125];
  assign o[64095] = i[125];
  assign o[64096] = i[125];
  assign o[64097] = i[125];
  assign o[64098] = i[125];
  assign o[64099] = i[125];
  assign o[64100] = i[125];
  assign o[64101] = i[125];
  assign o[64102] = i[125];
  assign o[64103] = i[125];
  assign o[64104] = i[125];
  assign o[64105] = i[125];
  assign o[64106] = i[125];
  assign o[64107] = i[125];
  assign o[64108] = i[125];
  assign o[64109] = i[125];
  assign o[64110] = i[125];
  assign o[64111] = i[125];
  assign o[64112] = i[125];
  assign o[64113] = i[125];
  assign o[64114] = i[125];
  assign o[64115] = i[125];
  assign o[64116] = i[125];
  assign o[64117] = i[125];
  assign o[64118] = i[125];
  assign o[64119] = i[125];
  assign o[64120] = i[125];
  assign o[64121] = i[125];
  assign o[64122] = i[125];
  assign o[64123] = i[125];
  assign o[64124] = i[125];
  assign o[64125] = i[125];
  assign o[64126] = i[125];
  assign o[64127] = i[125];
  assign o[64128] = i[125];
  assign o[64129] = i[125];
  assign o[64130] = i[125];
  assign o[64131] = i[125];
  assign o[64132] = i[125];
  assign o[64133] = i[125];
  assign o[64134] = i[125];
  assign o[64135] = i[125];
  assign o[64136] = i[125];
  assign o[64137] = i[125];
  assign o[64138] = i[125];
  assign o[64139] = i[125];
  assign o[64140] = i[125];
  assign o[64141] = i[125];
  assign o[64142] = i[125];
  assign o[64143] = i[125];
  assign o[64144] = i[125];
  assign o[64145] = i[125];
  assign o[64146] = i[125];
  assign o[64147] = i[125];
  assign o[64148] = i[125];
  assign o[64149] = i[125];
  assign o[64150] = i[125];
  assign o[64151] = i[125];
  assign o[64152] = i[125];
  assign o[64153] = i[125];
  assign o[64154] = i[125];
  assign o[64155] = i[125];
  assign o[64156] = i[125];
  assign o[64157] = i[125];
  assign o[64158] = i[125];
  assign o[64159] = i[125];
  assign o[64160] = i[125];
  assign o[64161] = i[125];
  assign o[64162] = i[125];
  assign o[64163] = i[125];
  assign o[64164] = i[125];
  assign o[64165] = i[125];
  assign o[64166] = i[125];
  assign o[64167] = i[125];
  assign o[64168] = i[125];
  assign o[64169] = i[125];
  assign o[64170] = i[125];
  assign o[64171] = i[125];
  assign o[64172] = i[125];
  assign o[64173] = i[125];
  assign o[64174] = i[125];
  assign o[64175] = i[125];
  assign o[64176] = i[125];
  assign o[64177] = i[125];
  assign o[64178] = i[125];
  assign o[64179] = i[125];
  assign o[64180] = i[125];
  assign o[64181] = i[125];
  assign o[64182] = i[125];
  assign o[64183] = i[125];
  assign o[64184] = i[125];
  assign o[64185] = i[125];
  assign o[64186] = i[125];
  assign o[64187] = i[125];
  assign o[64188] = i[125];
  assign o[64189] = i[125];
  assign o[64190] = i[125];
  assign o[64191] = i[125];
  assign o[64192] = i[125];
  assign o[64193] = i[125];
  assign o[64194] = i[125];
  assign o[64195] = i[125];
  assign o[64196] = i[125];
  assign o[64197] = i[125];
  assign o[64198] = i[125];
  assign o[64199] = i[125];
  assign o[64200] = i[125];
  assign o[64201] = i[125];
  assign o[64202] = i[125];
  assign o[64203] = i[125];
  assign o[64204] = i[125];
  assign o[64205] = i[125];
  assign o[64206] = i[125];
  assign o[64207] = i[125];
  assign o[64208] = i[125];
  assign o[64209] = i[125];
  assign o[64210] = i[125];
  assign o[64211] = i[125];
  assign o[64212] = i[125];
  assign o[64213] = i[125];
  assign o[64214] = i[125];
  assign o[64215] = i[125];
  assign o[64216] = i[125];
  assign o[64217] = i[125];
  assign o[64218] = i[125];
  assign o[64219] = i[125];
  assign o[64220] = i[125];
  assign o[64221] = i[125];
  assign o[64222] = i[125];
  assign o[64223] = i[125];
  assign o[64224] = i[125];
  assign o[64225] = i[125];
  assign o[64226] = i[125];
  assign o[64227] = i[125];
  assign o[64228] = i[125];
  assign o[64229] = i[125];
  assign o[64230] = i[125];
  assign o[64231] = i[125];
  assign o[64232] = i[125];
  assign o[64233] = i[125];
  assign o[64234] = i[125];
  assign o[64235] = i[125];
  assign o[64236] = i[125];
  assign o[64237] = i[125];
  assign o[64238] = i[125];
  assign o[64239] = i[125];
  assign o[64240] = i[125];
  assign o[64241] = i[125];
  assign o[64242] = i[125];
  assign o[64243] = i[125];
  assign o[64244] = i[125];
  assign o[64245] = i[125];
  assign o[64246] = i[125];
  assign o[64247] = i[125];
  assign o[64248] = i[125];
  assign o[64249] = i[125];
  assign o[64250] = i[125];
  assign o[64251] = i[125];
  assign o[64252] = i[125];
  assign o[64253] = i[125];
  assign o[64254] = i[125];
  assign o[64255] = i[125];
  assign o[64256] = i[125];
  assign o[64257] = i[125];
  assign o[64258] = i[125];
  assign o[64259] = i[125];
  assign o[64260] = i[125];
  assign o[64261] = i[125];
  assign o[64262] = i[125];
  assign o[64263] = i[125];
  assign o[64264] = i[125];
  assign o[64265] = i[125];
  assign o[64266] = i[125];
  assign o[64267] = i[125];
  assign o[64268] = i[125];
  assign o[64269] = i[125];
  assign o[64270] = i[125];
  assign o[64271] = i[125];
  assign o[64272] = i[125];
  assign o[64273] = i[125];
  assign o[64274] = i[125];
  assign o[64275] = i[125];
  assign o[64276] = i[125];
  assign o[64277] = i[125];
  assign o[64278] = i[125];
  assign o[64279] = i[125];
  assign o[64280] = i[125];
  assign o[64281] = i[125];
  assign o[64282] = i[125];
  assign o[64283] = i[125];
  assign o[64284] = i[125];
  assign o[64285] = i[125];
  assign o[64286] = i[125];
  assign o[64287] = i[125];
  assign o[64288] = i[125];
  assign o[64289] = i[125];
  assign o[64290] = i[125];
  assign o[64291] = i[125];
  assign o[64292] = i[125];
  assign o[64293] = i[125];
  assign o[64294] = i[125];
  assign o[64295] = i[125];
  assign o[64296] = i[125];
  assign o[64297] = i[125];
  assign o[64298] = i[125];
  assign o[64299] = i[125];
  assign o[64300] = i[125];
  assign o[64301] = i[125];
  assign o[64302] = i[125];
  assign o[64303] = i[125];
  assign o[64304] = i[125];
  assign o[64305] = i[125];
  assign o[64306] = i[125];
  assign o[64307] = i[125];
  assign o[64308] = i[125];
  assign o[64309] = i[125];
  assign o[64310] = i[125];
  assign o[64311] = i[125];
  assign o[64312] = i[125];
  assign o[64313] = i[125];
  assign o[64314] = i[125];
  assign o[64315] = i[125];
  assign o[64316] = i[125];
  assign o[64317] = i[125];
  assign o[64318] = i[125];
  assign o[64319] = i[125];
  assign o[64320] = i[125];
  assign o[64321] = i[125];
  assign o[64322] = i[125];
  assign o[64323] = i[125];
  assign o[64324] = i[125];
  assign o[64325] = i[125];
  assign o[64326] = i[125];
  assign o[64327] = i[125];
  assign o[64328] = i[125];
  assign o[64329] = i[125];
  assign o[64330] = i[125];
  assign o[64331] = i[125];
  assign o[64332] = i[125];
  assign o[64333] = i[125];
  assign o[64334] = i[125];
  assign o[64335] = i[125];
  assign o[64336] = i[125];
  assign o[64337] = i[125];
  assign o[64338] = i[125];
  assign o[64339] = i[125];
  assign o[64340] = i[125];
  assign o[64341] = i[125];
  assign o[64342] = i[125];
  assign o[64343] = i[125];
  assign o[64344] = i[125];
  assign o[64345] = i[125];
  assign o[64346] = i[125];
  assign o[64347] = i[125];
  assign o[64348] = i[125];
  assign o[64349] = i[125];
  assign o[64350] = i[125];
  assign o[64351] = i[125];
  assign o[64352] = i[125];
  assign o[64353] = i[125];
  assign o[64354] = i[125];
  assign o[64355] = i[125];
  assign o[64356] = i[125];
  assign o[64357] = i[125];
  assign o[64358] = i[125];
  assign o[64359] = i[125];
  assign o[64360] = i[125];
  assign o[64361] = i[125];
  assign o[64362] = i[125];
  assign o[64363] = i[125];
  assign o[64364] = i[125];
  assign o[64365] = i[125];
  assign o[64366] = i[125];
  assign o[64367] = i[125];
  assign o[64368] = i[125];
  assign o[64369] = i[125];
  assign o[64370] = i[125];
  assign o[64371] = i[125];
  assign o[64372] = i[125];
  assign o[64373] = i[125];
  assign o[64374] = i[125];
  assign o[64375] = i[125];
  assign o[64376] = i[125];
  assign o[64377] = i[125];
  assign o[64378] = i[125];
  assign o[64379] = i[125];
  assign o[64380] = i[125];
  assign o[64381] = i[125];
  assign o[64382] = i[125];
  assign o[64383] = i[125];
  assign o[64384] = i[125];
  assign o[64385] = i[125];
  assign o[64386] = i[125];
  assign o[64387] = i[125];
  assign o[64388] = i[125];
  assign o[64389] = i[125];
  assign o[64390] = i[125];
  assign o[64391] = i[125];
  assign o[64392] = i[125];
  assign o[64393] = i[125];
  assign o[64394] = i[125];
  assign o[64395] = i[125];
  assign o[64396] = i[125];
  assign o[64397] = i[125];
  assign o[64398] = i[125];
  assign o[64399] = i[125];
  assign o[64400] = i[125];
  assign o[64401] = i[125];
  assign o[64402] = i[125];
  assign o[64403] = i[125];
  assign o[64404] = i[125];
  assign o[64405] = i[125];
  assign o[64406] = i[125];
  assign o[64407] = i[125];
  assign o[64408] = i[125];
  assign o[64409] = i[125];
  assign o[64410] = i[125];
  assign o[64411] = i[125];
  assign o[64412] = i[125];
  assign o[64413] = i[125];
  assign o[64414] = i[125];
  assign o[64415] = i[125];
  assign o[64416] = i[125];
  assign o[64417] = i[125];
  assign o[64418] = i[125];
  assign o[64419] = i[125];
  assign o[64420] = i[125];
  assign o[64421] = i[125];
  assign o[64422] = i[125];
  assign o[64423] = i[125];
  assign o[64424] = i[125];
  assign o[64425] = i[125];
  assign o[64426] = i[125];
  assign o[64427] = i[125];
  assign o[64428] = i[125];
  assign o[64429] = i[125];
  assign o[64430] = i[125];
  assign o[64431] = i[125];
  assign o[64432] = i[125];
  assign o[64433] = i[125];
  assign o[64434] = i[125];
  assign o[64435] = i[125];
  assign o[64436] = i[125];
  assign o[64437] = i[125];
  assign o[64438] = i[125];
  assign o[64439] = i[125];
  assign o[64440] = i[125];
  assign o[64441] = i[125];
  assign o[64442] = i[125];
  assign o[64443] = i[125];
  assign o[64444] = i[125];
  assign o[64445] = i[125];
  assign o[64446] = i[125];
  assign o[64447] = i[125];
  assign o[64448] = i[125];
  assign o[64449] = i[125];
  assign o[64450] = i[125];
  assign o[64451] = i[125];
  assign o[64452] = i[125];
  assign o[64453] = i[125];
  assign o[64454] = i[125];
  assign o[64455] = i[125];
  assign o[64456] = i[125];
  assign o[64457] = i[125];
  assign o[64458] = i[125];
  assign o[64459] = i[125];
  assign o[64460] = i[125];
  assign o[64461] = i[125];
  assign o[64462] = i[125];
  assign o[64463] = i[125];
  assign o[64464] = i[125];
  assign o[64465] = i[125];
  assign o[64466] = i[125];
  assign o[64467] = i[125];
  assign o[64468] = i[125];
  assign o[64469] = i[125];
  assign o[64470] = i[125];
  assign o[64471] = i[125];
  assign o[64472] = i[125];
  assign o[64473] = i[125];
  assign o[64474] = i[125];
  assign o[64475] = i[125];
  assign o[64476] = i[125];
  assign o[64477] = i[125];
  assign o[64478] = i[125];
  assign o[64479] = i[125];
  assign o[64480] = i[125];
  assign o[64481] = i[125];
  assign o[64482] = i[125];
  assign o[64483] = i[125];
  assign o[64484] = i[125];
  assign o[64485] = i[125];
  assign o[64486] = i[125];
  assign o[64487] = i[125];
  assign o[64488] = i[125];
  assign o[64489] = i[125];
  assign o[64490] = i[125];
  assign o[64491] = i[125];
  assign o[64492] = i[125];
  assign o[64493] = i[125];
  assign o[64494] = i[125];
  assign o[64495] = i[125];
  assign o[64496] = i[125];
  assign o[64497] = i[125];
  assign o[64498] = i[125];
  assign o[64499] = i[125];
  assign o[64500] = i[125];
  assign o[64501] = i[125];
  assign o[64502] = i[125];
  assign o[64503] = i[125];
  assign o[64504] = i[125];
  assign o[64505] = i[125];
  assign o[64506] = i[125];
  assign o[64507] = i[125];
  assign o[64508] = i[125];
  assign o[64509] = i[125];
  assign o[64510] = i[125];
  assign o[64511] = i[125];
  assign o[63488] = i[124];
  assign o[63489] = i[124];
  assign o[63490] = i[124];
  assign o[63491] = i[124];
  assign o[63492] = i[124];
  assign o[63493] = i[124];
  assign o[63494] = i[124];
  assign o[63495] = i[124];
  assign o[63496] = i[124];
  assign o[63497] = i[124];
  assign o[63498] = i[124];
  assign o[63499] = i[124];
  assign o[63500] = i[124];
  assign o[63501] = i[124];
  assign o[63502] = i[124];
  assign o[63503] = i[124];
  assign o[63504] = i[124];
  assign o[63505] = i[124];
  assign o[63506] = i[124];
  assign o[63507] = i[124];
  assign o[63508] = i[124];
  assign o[63509] = i[124];
  assign o[63510] = i[124];
  assign o[63511] = i[124];
  assign o[63512] = i[124];
  assign o[63513] = i[124];
  assign o[63514] = i[124];
  assign o[63515] = i[124];
  assign o[63516] = i[124];
  assign o[63517] = i[124];
  assign o[63518] = i[124];
  assign o[63519] = i[124];
  assign o[63520] = i[124];
  assign o[63521] = i[124];
  assign o[63522] = i[124];
  assign o[63523] = i[124];
  assign o[63524] = i[124];
  assign o[63525] = i[124];
  assign o[63526] = i[124];
  assign o[63527] = i[124];
  assign o[63528] = i[124];
  assign o[63529] = i[124];
  assign o[63530] = i[124];
  assign o[63531] = i[124];
  assign o[63532] = i[124];
  assign o[63533] = i[124];
  assign o[63534] = i[124];
  assign o[63535] = i[124];
  assign o[63536] = i[124];
  assign o[63537] = i[124];
  assign o[63538] = i[124];
  assign o[63539] = i[124];
  assign o[63540] = i[124];
  assign o[63541] = i[124];
  assign o[63542] = i[124];
  assign o[63543] = i[124];
  assign o[63544] = i[124];
  assign o[63545] = i[124];
  assign o[63546] = i[124];
  assign o[63547] = i[124];
  assign o[63548] = i[124];
  assign o[63549] = i[124];
  assign o[63550] = i[124];
  assign o[63551] = i[124];
  assign o[63552] = i[124];
  assign o[63553] = i[124];
  assign o[63554] = i[124];
  assign o[63555] = i[124];
  assign o[63556] = i[124];
  assign o[63557] = i[124];
  assign o[63558] = i[124];
  assign o[63559] = i[124];
  assign o[63560] = i[124];
  assign o[63561] = i[124];
  assign o[63562] = i[124];
  assign o[63563] = i[124];
  assign o[63564] = i[124];
  assign o[63565] = i[124];
  assign o[63566] = i[124];
  assign o[63567] = i[124];
  assign o[63568] = i[124];
  assign o[63569] = i[124];
  assign o[63570] = i[124];
  assign o[63571] = i[124];
  assign o[63572] = i[124];
  assign o[63573] = i[124];
  assign o[63574] = i[124];
  assign o[63575] = i[124];
  assign o[63576] = i[124];
  assign o[63577] = i[124];
  assign o[63578] = i[124];
  assign o[63579] = i[124];
  assign o[63580] = i[124];
  assign o[63581] = i[124];
  assign o[63582] = i[124];
  assign o[63583] = i[124];
  assign o[63584] = i[124];
  assign o[63585] = i[124];
  assign o[63586] = i[124];
  assign o[63587] = i[124];
  assign o[63588] = i[124];
  assign o[63589] = i[124];
  assign o[63590] = i[124];
  assign o[63591] = i[124];
  assign o[63592] = i[124];
  assign o[63593] = i[124];
  assign o[63594] = i[124];
  assign o[63595] = i[124];
  assign o[63596] = i[124];
  assign o[63597] = i[124];
  assign o[63598] = i[124];
  assign o[63599] = i[124];
  assign o[63600] = i[124];
  assign o[63601] = i[124];
  assign o[63602] = i[124];
  assign o[63603] = i[124];
  assign o[63604] = i[124];
  assign o[63605] = i[124];
  assign o[63606] = i[124];
  assign o[63607] = i[124];
  assign o[63608] = i[124];
  assign o[63609] = i[124];
  assign o[63610] = i[124];
  assign o[63611] = i[124];
  assign o[63612] = i[124];
  assign o[63613] = i[124];
  assign o[63614] = i[124];
  assign o[63615] = i[124];
  assign o[63616] = i[124];
  assign o[63617] = i[124];
  assign o[63618] = i[124];
  assign o[63619] = i[124];
  assign o[63620] = i[124];
  assign o[63621] = i[124];
  assign o[63622] = i[124];
  assign o[63623] = i[124];
  assign o[63624] = i[124];
  assign o[63625] = i[124];
  assign o[63626] = i[124];
  assign o[63627] = i[124];
  assign o[63628] = i[124];
  assign o[63629] = i[124];
  assign o[63630] = i[124];
  assign o[63631] = i[124];
  assign o[63632] = i[124];
  assign o[63633] = i[124];
  assign o[63634] = i[124];
  assign o[63635] = i[124];
  assign o[63636] = i[124];
  assign o[63637] = i[124];
  assign o[63638] = i[124];
  assign o[63639] = i[124];
  assign o[63640] = i[124];
  assign o[63641] = i[124];
  assign o[63642] = i[124];
  assign o[63643] = i[124];
  assign o[63644] = i[124];
  assign o[63645] = i[124];
  assign o[63646] = i[124];
  assign o[63647] = i[124];
  assign o[63648] = i[124];
  assign o[63649] = i[124];
  assign o[63650] = i[124];
  assign o[63651] = i[124];
  assign o[63652] = i[124];
  assign o[63653] = i[124];
  assign o[63654] = i[124];
  assign o[63655] = i[124];
  assign o[63656] = i[124];
  assign o[63657] = i[124];
  assign o[63658] = i[124];
  assign o[63659] = i[124];
  assign o[63660] = i[124];
  assign o[63661] = i[124];
  assign o[63662] = i[124];
  assign o[63663] = i[124];
  assign o[63664] = i[124];
  assign o[63665] = i[124];
  assign o[63666] = i[124];
  assign o[63667] = i[124];
  assign o[63668] = i[124];
  assign o[63669] = i[124];
  assign o[63670] = i[124];
  assign o[63671] = i[124];
  assign o[63672] = i[124];
  assign o[63673] = i[124];
  assign o[63674] = i[124];
  assign o[63675] = i[124];
  assign o[63676] = i[124];
  assign o[63677] = i[124];
  assign o[63678] = i[124];
  assign o[63679] = i[124];
  assign o[63680] = i[124];
  assign o[63681] = i[124];
  assign o[63682] = i[124];
  assign o[63683] = i[124];
  assign o[63684] = i[124];
  assign o[63685] = i[124];
  assign o[63686] = i[124];
  assign o[63687] = i[124];
  assign o[63688] = i[124];
  assign o[63689] = i[124];
  assign o[63690] = i[124];
  assign o[63691] = i[124];
  assign o[63692] = i[124];
  assign o[63693] = i[124];
  assign o[63694] = i[124];
  assign o[63695] = i[124];
  assign o[63696] = i[124];
  assign o[63697] = i[124];
  assign o[63698] = i[124];
  assign o[63699] = i[124];
  assign o[63700] = i[124];
  assign o[63701] = i[124];
  assign o[63702] = i[124];
  assign o[63703] = i[124];
  assign o[63704] = i[124];
  assign o[63705] = i[124];
  assign o[63706] = i[124];
  assign o[63707] = i[124];
  assign o[63708] = i[124];
  assign o[63709] = i[124];
  assign o[63710] = i[124];
  assign o[63711] = i[124];
  assign o[63712] = i[124];
  assign o[63713] = i[124];
  assign o[63714] = i[124];
  assign o[63715] = i[124];
  assign o[63716] = i[124];
  assign o[63717] = i[124];
  assign o[63718] = i[124];
  assign o[63719] = i[124];
  assign o[63720] = i[124];
  assign o[63721] = i[124];
  assign o[63722] = i[124];
  assign o[63723] = i[124];
  assign o[63724] = i[124];
  assign o[63725] = i[124];
  assign o[63726] = i[124];
  assign o[63727] = i[124];
  assign o[63728] = i[124];
  assign o[63729] = i[124];
  assign o[63730] = i[124];
  assign o[63731] = i[124];
  assign o[63732] = i[124];
  assign o[63733] = i[124];
  assign o[63734] = i[124];
  assign o[63735] = i[124];
  assign o[63736] = i[124];
  assign o[63737] = i[124];
  assign o[63738] = i[124];
  assign o[63739] = i[124];
  assign o[63740] = i[124];
  assign o[63741] = i[124];
  assign o[63742] = i[124];
  assign o[63743] = i[124];
  assign o[63744] = i[124];
  assign o[63745] = i[124];
  assign o[63746] = i[124];
  assign o[63747] = i[124];
  assign o[63748] = i[124];
  assign o[63749] = i[124];
  assign o[63750] = i[124];
  assign o[63751] = i[124];
  assign o[63752] = i[124];
  assign o[63753] = i[124];
  assign o[63754] = i[124];
  assign o[63755] = i[124];
  assign o[63756] = i[124];
  assign o[63757] = i[124];
  assign o[63758] = i[124];
  assign o[63759] = i[124];
  assign o[63760] = i[124];
  assign o[63761] = i[124];
  assign o[63762] = i[124];
  assign o[63763] = i[124];
  assign o[63764] = i[124];
  assign o[63765] = i[124];
  assign o[63766] = i[124];
  assign o[63767] = i[124];
  assign o[63768] = i[124];
  assign o[63769] = i[124];
  assign o[63770] = i[124];
  assign o[63771] = i[124];
  assign o[63772] = i[124];
  assign o[63773] = i[124];
  assign o[63774] = i[124];
  assign o[63775] = i[124];
  assign o[63776] = i[124];
  assign o[63777] = i[124];
  assign o[63778] = i[124];
  assign o[63779] = i[124];
  assign o[63780] = i[124];
  assign o[63781] = i[124];
  assign o[63782] = i[124];
  assign o[63783] = i[124];
  assign o[63784] = i[124];
  assign o[63785] = i[124];
  assign o[63786] = i[124];
  assign o[63787] = i[124];
  assign o[63788] = i[124];
  assign o[63789] = i[124];
  assign o[63790] = i[124];
  assign o[63791] = i[124];
  assign o[63792] = i[124];
  assign o[63793] = i[124];
  assign o[63794] = i[124];
  assign o[63795] = i[124];
  assign o[63796] = i[124];
  assign o[63797] = i[124];
  assign o[63798] = i[124];
  assign o[63799] = i[124];
  assign o[63800] = i[124];
  assign o[63801] = i[124];
  assign o[63802] = i[124];
  assign o[63803] = i[124];
  assign o[63804] = i[124];
  assign o[63805] = i[124];
  assign o[63806] = i[124];
  assign o[63807] = i[124];
  assign o[63808] = i[124];
  assign o[63809] = i[124];
  assign o[63810] = i[124];
  assign o[63811] = i[124];
  assign o[63812] = i[124];
  assign o[63813] = i[124];
  assign o[63814] = i[124];
  assign o[63815] = i[124];
  assign o[63816] = i[124];
  assign o[63817] = i[124];
  assign o[63818] = i[124];
  assign o[63819] = i[124];
  assign o[63820] = i[124];
  assign o[63821] = i[124];
  assign o[63822] = i[124];
  assign o[63823] = i[124];
  assign o[63824] = i[124];
  assign o[63825] = i[124];
  assign o[63826] = i[124];
  assign o[63827] = i[124];
  assign o[63828] = i[124];
  assign o[63829] = i[124];
  assign o[63830] = i[124];
  assign o[63831] = i[124];
  assign o[63832] = i[124];
  assign o[63833] = i[124];
  assign o[63834] = i[124];
  assign o[63835] = i[124];
  assign o[63836] = i[124];
  assign o[63837] = i[124];
  assign o[63838] = i[124];
  assign o[63839] = i[124];
  assign o[63840] = i[124];
  assign o[63841] = i[124];
  assign o[63842] = i[124];
  assign o[63843] = i[124];
  assign o[63844] = i[124];
  assign o[63845] = i[124];
  assign o[63846] = i[124];
  assign o[63847] = i[124];
  assign o[63848] = i[124];
  assign o[63849] = i[124];
  assign o[63850] = i[124];
  assign o[63851] = i[124];
  assign o[63852] = i[124];
  assign o[63853] = i[124];
  assign o[63854] = i[124];
  assign o[63855] = i[124];
  assign o[63856] = i[124];
  assign o[63857] = i[124];
  assign o[63858] = i[124];
  assign o[63859] = i[124];
  assign o[63860] = i[124];
  assign o[63861] = i[124];
  assign o[63862] = i[124];
  assign o[63863] = i[124];
  assign o[63864] = i[124];
  assign o[63865] = i[124];
  assign o[63866] = i[124];
  assign o[63867] = i[124];
  assign o[63868] = i[124];
  assign o[63869] = i[124];
  assign o[63870] = i[124];
  assign o[63871] = i[124];
  assign o[63872] = i[124];
  assign o[63873] = i[124];
  assign o[63874] = i[124];
  assign o[63875] = i[124];
  assign o[63876] = i[124];
  assign o[63877] = i[124];
  assign o[63878] = i[124];
  assign o[63879] = i[124];
  assign o[63880] = i[124];
  assign o[63881] = i[124];
  assign o[63882] = i[124];
  assign o[63883] = i[124];
  assign o[63884] = i[124];
  assign o[63885] = i[124];
  assign o[63886] = i[124];
  assign o[63887] = i[124];
  assign o[63888] = i[124];
  assign o[63889] = i[124];
  assign o[63890] = i[124];
  assign o[63891] = i[124];
  assign o[63892] = i[124];
  assign o[63893] = i[124];
  assign o[63894] = i[124];
  assign o[63895] = i[124];
  assign o[63896] = i[124];
  assign o[63897] = i[124];
  assign o[63898] = i[124];
  assign o[63899] = i[124];
  assign o[63900] = i[124];
  assign o[63901] = i[124];
  assign o[63902] = i[124];
  assign o[63903] = i[124];
  assign o[63904] = i[124];
  assign o[63905] = i[124];
  assign o[63906] = i[124];
  assign o[63907] = i[124];
  assign o[63908] = i[124];
  assign o[63909] = i[124];
  assign o[63910] = i[124];
  assign o[63911] = i[124];
  assign o[63912] = i[124];
  assign o[63913] = i[124];
  assign o[63914] = i[124];
  assign o[63915] = i[124];
  assign o[63916] = i[124];
  assign o[63917] = i[124];
  assign o[63918] = i[124];
  assign o[63919] = i[124];
  assign o[63920] = i[124];
  assign o[63921] = i[124];
  assign o[63922] = i[124];
  assign o[63923] = i[124];
  assign o[63924] = i[124];
  assign o[63925] = i[124];
  assign o[63926] = i[124];
  assign o[63927] = i[124];
  assign o[63928] = i[124];
  assign o[63929] = i[124];
  assign o[63930] = i[124];
  assign o[63931] = i[124];
  assign o[63932] = i[124];
  assign o[63933] = i[124];
  assign o[63934] = i[124];
  assign o[63935] = i[124];
  assign o[63936] = i[124];
  assign o[63937] = i[124];
  assign o[63938] = i[124];
  assign o[63939] = i[124];
  assign o[63940] = i[124];
  assign o[63941] = i[124];
  assign o[63942] = i[124];
  assign o[63943] = i[124];
  assign o[63944] = i[124];
  assign o[63945] = i[124];
  assign o[63946] = i[124];
  assign o[63947] = i[124];
  assign o[63948] = i[124];
  assign o[63949] = i[124];
  assign o[63950] = i[124];
  assign o[63951] = i[124];
  assign o[63952] = i[124];
  assign o[63953] = i[124];
  assign o[63954] = i[124];
  assign o[63955] = i[124];
  assign o[63956] = i[124];
  assign o[63957] = i[124];
  assign o[63958] = i[124];
  assign o[63959] = i[124];
  assign o[63960] = i[124];
  assign o[63961] = i[124];
  assign o[63962] = i[124];
  assign o[63963] = i[124];
  assign o[63964] = i[124];
  assign o[63965] = i[124];
  assign o[63966] = i[124];
  assign o[63967] = i[124];
  assign o[63968] = i[124];
  assign o[63969] = i[124];
  assign o[63970] = i[124];
  assign o[63971] = i[124];
  assign o[63972] = i[124];
  assign o[63973] = i[124];
  assign o[63974] = i[124];
  assign o[63975] = i[124];
  assign o[63976] = i[124];
  assign o[63977] = i[124];
  assign o[63978] = i[124];
  assign o[63979] = i[124];
  assign o[63980] = i[124];
  assign o[63981] = i[124];
  assign o[63982] = i[124];
  assign o[63983] = i[124];
  assign o[63984] = i[124];
  assign o[63985] = i[124];
  assign o[63986] = i[124];
  assign o[63987] = i[124];
  assign o[63988] = i[124];
  assign o[63989] = i[124];
  assign o[63990] = i[124];
  assign o[63991] = i[124];
  assign o[63992] = i[124];
  assign o[63993] = i[124];
  assign o[63994] = i[124];
  assign o[63995] = i[124];
  assign o[63996] = i[124];
  assign o[63997] = i[124];
  assign o[63998] = i[124];
  assign o[63999] = i[124];
  assign o[62976] = i[123];
  assign o[62977] = i[123];
  assign o[62978] = i[123];
  assign o[62979] = i[123];
  assign o[62980] = i[123];
  assign o[62981] = i[123];
  assign o[62982] = i[123];
  assign o[62983] = i[123];
  assign o[62984] = i[123];
  assign o[62985] = i[123];
  assign o[62986] = i[123];
  assign o[62987] = i[123];
  assign o[62988] = i[123];
  assign o[62989] = i[123];
  assign o[62990] = i[123];
  assign o[62991] = i[123];
  assign o[62992] = i[123];
  assign o[62993] = i[123];
  assign o[62994] = i[123];
  assign o[62995] = i[123];
  assign o[62996] = i[123];
  assign o[62997] = i[123];
  assign o[62998] = i[123];
  assign o[62999] = i[123];
  assign o[63000] = i[123];
  assign o[63001] = i[123];
  assign o[63002] = i[123];
  assign o[63003] = i[123];
  assign o[63004] = i[123];
  assign o[63005] = i[123];
  assign o[63006] = i[123];
  assign o[63007] = i[123];
  assign o[63008] = i[123];
  assign o[63009] = i[123];
  assign o[63010] = i[123];
  assign o[63011] = i[123];
  assign o[63012] = i[123];
  assign o[63013] = i[123];
  assign o[63014] = i[123];
  assign o[63015] = i[123];
  assign o[63016] = i[123];
  assign o[63017] = i[123];
  assign o[63018] = i[123];
  assign o[63019] = i[123];
  assign o[63020] = i[123];
  assign o[63021] = i[123];
  assign o[63022] = i[123];
  assign o[63023] = i[123];
  assign o[63024] = i[123];
  assign o[63025] = i[123];
  assign o[63026] = i[123];
  assign o[63027] = i[123];
  assign o[63028] = i[123];
  assign o[63029] = i[123];
  assign o[63030] = i[123];
  assign o[63031] = i[123];
  assign o[63032] = i[123];
  assign o[63033] = i[123];
  assign o[63034] = i[123];
  assign o[63035] = i[123];
  assign o[63036] = i[123];
  assign o[63037] = i[123];
  assign o[63038] = i[123];
  assign o[63039] = i[123];
  assign o[63040] = i[123];
  assign o[63041] = i[123];
  assign o[63042] = i[123];
  assign o[63043] = i[123];
  assign o[63044] = i[123];
  assign o[63045] = i[123];
  assign o[63046] = i[123];
  assign o[63047] = i[123];
  assign o[63048] = i[123];
  assign o[63049] = i[123];
  assign o[63050] = i[123];
  assign o[63051] = i[123];
  assign o[63052] = i[123];
  assign o[63053] = i[123];
  assign o[63054] = i[123];
  assign o[63055] = i[123];
  assign o[63056] = i[123];
  assign o[63057] = i[123];
  assign o[63058] = i[123];
  assign o[63059] = i[123];
  assign o[63060] = i[123];
  assign o[63061] = i[123];
  assign o[63062] = i[123];
  assign o[63063] = i[123];
  assign o[63064] = i[123];
  assign o[63065] = i[123];
  assign o[63066] = i[123];
  assign o[63067] = i[123];
  assign o[63068] = i[123];
  assign o[63069] = i[123];
  assign o[63070] = i[123];
  assign o[63071] = i[123];
  assign o[63072] = i[123];
  assign o[63073] = i[123];
  assign o[63074] = i[123];
  assign o[63075] = i[123];
  assign o[63076] = i[123];
  assign o[63077] = i[123];
  assign o[63078] = i[123];
  assign o[63079] = i[123];
  assign o[63080] = i[123];
  assign o[63081] = i[123];
  assign o[63082] = i[123];
  assign o[63083] = i[123];
  assign o[63084] = i[123];
  assign o[63085] = i[123];
  assign o[63086] = i[123];
  assign o[63087] = i[123];
  assign o[63088] = i[123];
  assign o[63089] = i[123];
  assign o[63090] = i[123];
  assign o[63091] = i[123];
  assign o[63092] = i[123];
  assign o[63093] = i[123];
  assign o[63094] = i[123];
  assign o[63095] = i[123];
  assign o[63096] = i[123];
  assign o[63097] = i[123];
  assign o[63098] = i[123];
  assign o[63099] = i[123];
  assign o[63100] = i[123];
  assign o[63101] = i[123];
  assign o[63102] = i[123];
  assign o[63103] = i[123];
  assign o[63104] = i[123];
  assign o[63105] = i[123];
  assign o[63106] = i[123];
  assign o[63107] = i[123];
  assign o[63108] = i[123];
  assign o[63109] = i[123];
  assign o[63110] = i[123];
  assign o[63111] = i[123];
  assign o[63112] = i[123];
  assign o[63113] = i[123];
  assign o[63114] = i[123];
  assign o[63115] = i[123];
  assign o[63116] = i[123];
  assign o[63117] = i[123];
  assign o[63118] = i[123];
  assign o[63119] = i[123];
  assign o[63120] = i[123];
  assign o[63121] = i[123];
  assign o[63122] = i[123];
  assign o[63123] = i[123];
  assign o[63124] = i[123];
  assign o[63125] = i[123];
  assign o[63126] = i[123];
  assign o[63127] = i[123];
  assign o[63128] = i[123];
  assign o[63129] = i[123];
  assign o[63130] = i[123];
  assign o[63131] = i[123];
  assign o[63132] = i[123];
  assign o[63133] = i[123];
  assign o[63134] = i[123];
  assign o[63135] = i[123];
  assign o[63136] = i[123];
  assign o[63137] = i[123];
  assign o[63138] = i[123];
  assign o[63139] = i[123];
  assign o[63140] = i[123];
  assign o[63141] = i[123];
  assign o[63142] = i[123];
  assign o[63143] = i[123];
  assign o[63144] = i[123];
  assign o[63145] = i[123];
  assign o[63146] = i[123];
  assign o[63147] = i[123];
  assign o[63148] = i[123];
  assign o[63149] = i[123];
  assign o[63150] = i[123];
  assign o[63151] = i[123];
  assign o[63152] = i[123];
  assign o[63153] = i[123];
  assign o[63154] = i[123];
  assign o[63155] = i[123];
  assign o[63156] = i[123];
  assign o[63157] = i[123];
  assign o[63158] = i[123];
  assign o[63159] = i[123];
  assign o[63160] = i[123];
  assign o[63161] = i[123];
  assign o[63162] = i[123];
  assign o[63163] = i[123];
  assign o[63164] = i[123];
  assign o[63165] = i[123];
  assign o[63166] = i[123];
  assign o[63167] = i[123];
  assign o[63168] = i[123];
  assign o[63169] = i[123];
  assign o[63170] = i[123];
  assign o[63171] = i[123];
  assign o[63172] = i[123];
  assign o[63173] = i[123];
  assign o[63174] = i[123];
  assign o[63175] = i[123];
  assign o[63176] = i[123];
  assign o[63177] = i[123];
  assign o[63178] = i[123];
  assign o[63179] = i[123];
  assign o[63180] = i[123];
  assign o[63181] = i[123];
  assign o[63182] = i[123];
  assign o[63183] = i[123];
  assign o[63184] = i[123];
  assign o[63185] = i[123];
  assign o[63186] = i[123];
  assign o[63187] = i[123];
  assign o[63188] = i[123];
  assign o[63189] = i[123];
  assign o[63190] = i[123];
  assign o[63191] = i[123];
  assign o[63192] = i[123];
  assign o[63193] = i[123];
  assign o[63194] = i[123];
  assign o[63195] = i[123];
  assign o[63196] = i[123];
  assign o[63197] = i[123];
  assign o[63198] = i[123];
  assign o[63199] = i[123];
  assign o[63200] = i[123];
  assign o[63201] = i[123];
  assign o[63202] = i[123];
  assign o[63203] = i[123];
  assign o[63204] = i[123];
  assign o[63205] = i[123];
  assign o[63206] = i[123];
  assign o[63207] = i[123];
  assign o[63208] = i[123];
  assign o[63209] = i[123];
  assign o[63210] = i[123];
  assign o[63211] = i[123];
  assign o[63212] = i[123];
  assign o[63213] = i[123];
  assign o[63214] = i[123];
  assign o[63215] = i[123];
  assign o[63216] = i[123];
  assign o[63217] = i[123];
  assign o[63218] = i[123];
  assign o[63219] = i[123];
  assign o[63220] = i[123];
  assign o[63221] = i[123];
  assign o[63222] = i[123];
  assign o[63223] = i[123];
  assign o[63224] = i[123];
  assign o[63225] = i[123];
  assign o[63226] = i[123];
  assign o[63227] = i[123];
  assign o[63228] = i[123];
  assign o[63229] = i[123];
  assign o[63230] = i[123];
  assign o[63231] = i[123];
  assign o[63232] = i[123];
  assign o[63233] = i[123];
  assign o[63234] = i[123];
  assign o[63235] = i[123];
  assign o[63236] = i[123];
  assign o[63237] = i[123];
  assign o[63238] = i[123];
  assign o[63239] = i[123];
  assign o[63240] = i[123];
  assign o[63241] = i[123];
  assign o[63242] = i[123];
  assign o[63243] = i[123];
  assign o[63244] = i[123];
  assign o[63245] = i[123];
  assign o[63246] = i[123];
  assign o[63247] = i[123];
  assign o[63248] = i[123];
  assign o[63249] = i[123];
  assign o[63250] = i[123];
  assign o[63251] = i[123];
  assign o[63252] = i[123];
  assign o[63253] = i[123];
  assign o[63254] = i[123];
  assign o[63255] = i[123];
  assign o[63256] = i[123];
  assign o[63257] = i[123];
  assign o[63258] = i[123];
  assign o[63259] = i[123];
  assign o[63260] = i[123];
  assign o[63261] = i[123];
  assign o[63262] = i[123];
  assign o[63263] = i[123];
  assign o[63264] = i[123];
  assign o[63265] = i[123];
  assign o[63266] = i[123];
  assign o[63267] = i[123];
  assign o[63268] = i[123];
  assign o[63269] = i[123];
  assign o[63270] = i[123];
  assign o[63271] = i[123];
  assign o[63272] = i[123];
  assign o[63273] = i[123];
  assign o[63274] = i[123];
  assign o[63275] = i[123];
  assign o[63276] = i[123];
  assign o[63277] = i[123];
  assign o[63278] = i[123];
  assign o[63279] = i[123];
  assign o[63280] = i[123];
  assign o[63281] = i[123];
  assign o[63282] = i[123];
  assign o[63283] = i[123];
  assign o[63284] = i[123];
  assign o[63285] = i[123];
  assign o[63286] = i[123];
  assign o[63287] = i[123];
  assign o[63288] = i[123];
  assign o[63289] = i[123];
  assign o[63290] = i[123];
  assign o[63291] = i[123];
  assign o[63292] = i[123];
  assign o[63293] = i[123];
  assign o[63294] = i[123];
  assign o[63295] = i[123];
  assign o[63296] = i[123];
  assign o[63297] = i[123];
  assign o[63298] = i[123];
  assign o[63299] = i[123];
  assign o[63300] = i[123];
  assign o[63301] = i[123];
  assign o[63302] = i[123];
  assign o[63303] = i[123];
  assign o[63304] = i[123];
  assign o[63305] = i[123];
  assign o[63306] = i[123];
  assign o[63307] = i[123];
  assign o[63308] = i[123];
  assign o[63309] = i[123];
  assign o[63310] = i[123];
  assign o[63311] = i[123];
  assign o[63312] = i[123];
  assign o[63313] = i[123];
  assign o[63314] = i[123];
  assign o[63315] = i[123];
  assign o[63316] = i[123];
  assign o[63317] = i[123];
  assign o[63318] = i[123];
  assign o[63319] = i[123];
  assign o[63320] = i[123];
  assign o[63321] = i[123];
  assign o[63322] = i[123];
  assign o[63323] = i[123];
  assign o[63324] = i[123];
  assign o[63325] = i[123];
  assign o[63326] = i[123];
  assign o[63327] = i[123];
  assign o[63328] = i[123];
  assign o[63329] = i[123];
  assign o[63330] = i[123];
  assign o[63331] = i[123];
  assign o[63332] = i[123];
  assign o[63333] = i[123];
  assign o[63334] = i[123];
  assign o[63335] = i[123];
  assign o[63336] = i[123];
  assign o[63337] = i[123];
  assign o[63338] = i[123];
  assign o[63339] = i[123];
  assign o[63340] = i[123];
  assign o[63341] = i[123];
  assign o[63342] = i[123];
  assign o[63343] = i[123];
  assign o[63344] = i[123];
  assign o[63345] = i[123];
  assign o[63346] = i[123];
  assign o[63347] = i[123];
  assign o[63348] = i[123];
  assign o[63349] = i[123];
  assign o[63350] = i[123];
  assign o[63351] = i[123];
  assign o[63352] = i[123];
  assign o[63353] = i[123];
  assign o[63354] = i[123];
  assign o[63355] = i[123];
  assign o[63356] = i[123];
  assign o[63357] = i[123];
  assign o[63358] = i[123];
  assign o[63359] = i[123];
  assign o[63360] = i[123];
  assign o[63361] = i[123];
  assign o[63362] = i[123];
  assign o[63363] = i[123];
  assign o[63364] = i[123];
  assign o[63365] = i[123];
  assign o[63366] = i[123];
  assign o[63367] = i[123];
  assign o[63368] = i[123];
  assign o[63369] = i[123];
  assign o[63370] = i[123];
  assign o[63371] = i[123];
  assign o[63372] = i[123];
  assign o[63373] = i[123];
  assign o[63374] = i[123];
  assign o[63375] = i[123];
  assign o[63376] = i[123];
  assign o[63377] = i[123];
  assign o[63378] = i[123];
  assign o[63379] = i[123];
  assign o[63380] = i[123];
  assign o[63381] = i[123];
  assign o[63382] = i[123];
  assign o[63383] = i[123];
  assign o[63384] = i[123];
  assign o[63385] = i[123];
  assign o[63386] = i[123];
  assign o[63387] = i[123];
  assign o[63388] = i[123];
  assign o[63389] = i[123];
  assign o[63390] = i[123];
  assign o[63391] = i[123];
  assign o[63392] = i[123];
  assign o[63393] = i[123];
  assign o[63394] = i[123];
  assign o[63395] = i[123];
  assign o[63396] = i[123];
  assign o[63397] = i[123];
  assign o[63398] = i[123];
  assign o[63399] = i[123];
  assign o[63400] = i[123];
  assign o[63401] = i[123];
  assign o[63402] = i[123];
  assign o[63403] = i[123];
  assign o[63404] = i[123];
  assign o[63405] = i[123];
  assign o[63406] = i[123];
  assign o[63407] = i[123];
  assign o[63408] = i[123];
  assign o[63409] = i[123];
  assign o[63410] = i[123];
  assign o[63411] = i[123];
  assign o[63412] = i[123];
  assign o[63413] = i[123];
  assign o[63414] = i[123];
  assign o[63415] = i[123];
  assign o[63416] = i[123];
  assign o[63417] = i[123];
  assign o[63418] = i[123];
  assign o[63419] = i[123];
  assign o[63420] = i[123];
  assign o[63421] = i[123];
  assign o[63422] = i[123];
  assign o[63423] = i[123];
  assign o[63424] = i[123];
  assign o[63425] = i[123];
  assign o[63426] = i[123];
  assign o[63427] = i[123];
  assign o[63428] = i[123];
  assign o[63429] = i[123];
  assign o[63430] = i[123];
  assign o[63431] = i[123];
  assign o[63432] = i[123];
  assign o[63433] = i[123];
  assign o[63434] = i[123];
  assign o[63435] = i[123];
  assign o[63436] = i[123];
  assign o[63437] = i[123];
  assign o[63438] = i[123];
  assign o[63439] = i[123];
  assign o[63440] = i[123];
  assign o[63441] = i[123];
  assign o[63442] = i[123];
  assign o[63443] = i[123];
  assign o[63444] = i[123];
  assign o[63445] = i[123];
  assign o[63446] = i[123];
  assign o[63447] = i[123];
  assign o[63448] = i[123];
  assign o[63449] = i[123];
  assign o[63450] = i[123];
  assign o[63451] = i[123];
  assign o[63452] = i[123];
  assign o[63453] = i[123];
  assign o[63454] = i[123];
  assign o[63455] = i[123];
  assign o[63456] = i[123];
  assign o[63457] = i[123];
  assign o[63458] = i[123];
  assign o[63459] = i[123];
  assign o[63460] = i[123];
  assign o[63461] = i[123];
  assign o[63462] = i[123];
  assign o[63463] = i[123];
  assign o[63464] = i[123];
  assign o[63465] = i[123];
  assign o[63466] = i[123];
  assign o[63467] = i[123];
  assign o[63468] = i[123];
  assign o[63469] = i[123];
  assign o[63470] = i[123];
  assign o[63471] = i[123];
  assign o[63472] = i[123];
  assign o[63473] = i[123];
  assign o[63474] = i[123];
  assign o[63475] = i[123];
  assign o[63476] = i[123];
  assign o[63477] = i[123];
  assign o[63478] = i[123];
  assign o[63479] = i[123];
  assign o[63480] = i[123];
  assign o[63481] = i[123];
  assign o[63482] = i[123];
  assign o[63483] = i[123];
  assign o[63484] = i[123];
  assign o[63485] = i[123];
  assign o[63486] = i[123];
  assign o[63487] = i[123];
  assign o[62464] = i[122];
  assign o[62465] = i[122];
  assign o[62466] = i[122];
  assign o[62467] = i[122];
  assign o[62468] = i[122];
  assign o[62469] = i[122];
  assign o[62470] = i[122];
  assign o[62471] = i[122];
  assign o[62472] = i[122];
  assign o[62473] = i[122];
  assign o[62474] = i[122];
  assign o[62475] = i[122];
  assign o[62476] = i[122];
  assign o[62477] = i[122];
  assign o[62478] = i[122];
  assign o[62479] = i[122];
  assign o[62480] = i[122];
  assign o[62481] = i[122];
  assign o[62482] = i[122];
  assign o[62483] = i[122];
  assign o[62484] = i[122];
  assign o[62485] = i[122];
  assign o[62486] = i[122];
  assign o[62487] = i[122];
  assign o[62488] = i[122];
  assign o[62489] = i[122];
  assign o[62490] = i[122];
  assign o[62491] = i[122];
  assign o[62492] = i[122];
  assign o[62493] = i[122];
  assign o[62494] = i[122];
  assign o[62495] = i[122];
  assign o[62496] = i[122];
  assign o[62497] = i[122];
  assign o[62498] = i[122];
  assign o[62499] = i[122];
  assign o[62500] = i[122];
  assign o[62501] = i[122];
  assign o[62502] = i[122];
  assign o[62503] = i[122];
  assign o[62504] = i[122];
  assign o[62505] = i[122];
  assign o[62506] = i[122];
  assign o[62507] = i[122];
  assign o[62508] = i[122];
  assign o[62509] = i[122];
  assign o[62510] = i[122];
  assign o[62511] = i[122];
  assign o[62512] = i[122];
  assign o[62513] = i[122];
  assign o[62514] = i[122];
  assign o[62515] = i[122];
  assign o[62516] = i[122];
  assign o[62517] = i[122];
  assign o[62518] = i[122];
  assign o[62519] = i[122];
  assign o[62520] = i[122];
  assign o[62521] = i[122];
  assign o[62522] = i[122];
  assign o[62523] = i[122];
  assign o[62524] = i[122];
  assign o[62525] = i[122];
  assign o[62526] = i[122];
  assign o[62527] = i[122];
  assign o[62528] = i[122];
  assign o[62529] = i[122];
  assign o[62530] = i[122];
  assign o[62531] = i[122];
  assign o[62532] = i[122];
  assign o[62533] = i[122];
  assign o[62534] = i[122];
  assign o[62535] = i[122];
  assign o[62536] = i[122];
  assign o[62537] = i[122];
  assign o[62538] = i[122];
  assign o[62539] = i[122];
  assign o[62540] = i[122];
  assign o[62541] = i[122];
  assign o[62542] = i[122];
  assign o[62543] = i[122];
  assign o[62544] = i[122];
  assign o[62545] = i[122];
  assign o[62546] = i[122];
  assign o[62547] = i[122];
  assign o[62548] = i[122];
  assign o[62549] = i[122];
  assign o[62550] = i[122];
  assign o[62551] = i[122];
  assign o[62552] = i[122];
  assign o[62553] = i[122];
  assign o[62554] = i[122];
  assign o[62555] = i[122];
  assign o[62556] = i[122];
  assign o[62557] = i[122];
  assign o[62558] = i[122];
  assign o[62559] = i[122];
  assign o[62560] = i[122];
  assign o[62561] = i[122];
  assign o[62562] = i[122];
  assign o[62563] = i[122];
  assign o[62564] = i[122];
  assign o[62565] = i[122];
  assign o[62566] = i[122];
  assign o[62567] = i[122];
  assign o[62568] = i[122];
  assign o[62569] = i[122];
  assign o[62570] = i[122];
  assign o[62571] = i[122];
  assign o[62572] = i[122];
  assign o[62573] = i[122];
  assign o[62574] = i[122];
  assign o[62575] = i[122];
  assign o[62576] = i[122];
  assign o[62577] = i[122];
  assign o[62578] = i[122];
  assign o[62579] = i[122];
  assign o[62580] = i[122];
  assign o[62581] = i[122];
  assign o[62582] = i[122];
  assign o[62583] = i[122];
  assign o[62584] = i[122];
  assign o[62585] = i[122];
  assign o[62586] = i[122];
  assign o[62587] = i[122];
  assign o[62588] = i[122];
  assign o[62589] = i[122];
  assign o[62590] = i[122];
  assign o[62591] = i[122];
  assign o[62592] = i[122];
  assign o[62593] = i[122];
  assign o[62594] = i[122];
  assign o[62595] = i[122];
  assign o[62596] = i[122];
  assign o[62597] = i[122];
  assign o[62598] = i[122];
  assign o[62599] = i[122];
  assign o[62600] = i[122];
  assign o[62601] = i[122];
  assign o[62602] = i[122];
  assign o[62603] = i[122];
  assign o[62604] = i[122];
  assign o[62605] = i[122];
  assign o[62606] = i[122];
  assign o[62607] = i[122];
  assign o[62608] = i[122];
  assign o[62609] = i[122];
  assign o[62610] = i[122];
  assign o[62611] = i[122];
  assign o[62612] = i[122];
  assign o[62613] = i[122];
  assign o[62614] = i[122];
  assign o[62615] = i[122];
  assign o[62616] = i[122];
  assign o[62617] = i[122];
  assign o[62618] = i[122];
  assign o[62619] = i[122];
  assign o[62620] = i[122];
  assign o[62621] = i[122];
  assign o[62622] = i[122];
  assign o[62623] = i[122];
  assign o[62624] = i[122];
  assign o[62625] = i[122];
  assign o[62626] = i[122];
  assign o[62627] = i[122];
  assign o[62628] = i[122];
  assign o[62629] = i[122];
  assign o[62630] = i[122];
  assign o[62631] = i[122];
  assign o[62632] = i[122];
  assign o[62633] = i[122];
  assign o[62634] = i[122];
  assign o[62635] = i[122];
  assign o[62636] = i[122];
  assign o[62637] = i[122];
  assign o[62638] = i[122];
  assign o[62639] = i[122];
  assign o[62640] = i[122];
  assign o[62641] = i[122];
  assign o[62642] = i[122];
  assign o[62643] = i[122];
  assign o[62644] = i[122];
  assign o[62645] = i[122];
  assign o[62646] = i[122];
  assign o[62647] = i[122];
  assign o[62648] = i[122];
  assign o[62649] = i[122];
  assign o[62650] = i[122];
  assign o[62651] = i[122];
  assign o[62652] = i[122];
  assign o[62653] = i[122];
  assign o[62654] = i[122];
  assign o[62655] = i[122];
  assign o[62656] = i[122];
  assign o[62657] = i[122];
  assign o[62658] = i[122];
  assign o[62659] = i[122];
  assign o[62660] = i[122];
  assign o[62661] = i[122];
  assign o[62662] = i[122];
  assign o[62663] = i[122];
  assign o[62664] = i[122];
  assign o[62665] = i[122];
  assign o[62666] = i[122];
  assign o[62667] = i[122];
  assign o[62668] = i[122];
  assign o[62669] = i[122];
  assign o[62670] = i[122];
  assign o[62671] = i[122];
  assign o[62672] = i[122];
  assign o[62673] = i[122];
  assign o[62674] = i[122];
  assign o[62675] = i[122];
  assign o[62676] = i[122];
  assign o[62677] = i[122];
  assign o[62678] = i[122];
  assign o[62679] = i[122];
  assign o[62680] = i[122];
  assign o[62681] = i[122];
  assign o[62682] = i[122];
  assign o[62683] = i[122];
  assign o[62684] = i[122];
  assign o[62685] = i[122];
  assign o[62686] = i[122];
  assign o[62687] = i[122];
  assign o[62688] = i[122];
  assign o[62689] = i[122];
  assign o[62690] = i[122];
  assign o[62691] = i[122];
  assign o[62692] = i[122];
  assign o[62693] = i[122];
  assign o[62694] = i[122];
  assign o[62695] = i[122];
  assign o[62696] = i[122];
  assign o[62697] = i[122];
  assign o[62698] = i[122];
  assign o[62699] = i[122];
  assign o[62700] = i[122];
  assign o[62701] = i[122];
  assign o[62702] = i[122];
  assign o[62703] = i[122];
  assign o[62704] = i[122];
  assign o[62705] = i[122];
  assign o[62706] = i[122];
  assign o[62707] = i[122];
  assign o[62708] = i[122];
  assign o[62709] = i[122];
  assign o[62710] = i[122];
  assign o[62711] = i[122];
  assign o[62712] = i[122];
  assign o[62713] = i[122];
  assign o[62714] = i[122];
  assign o[62715] = i[122];
  assign o[62716] = i[122];
  assign o[62717] = i[122];
  assign o[62718] = i[122];
  assign o[62719] = i[122];
  assign o[62720] = i[122];
  assign o[62721] = i[122];
  assign o[62722] = i[122];
  assign o[62723] = i[122];
  assign o[62724] = i[122];
  assign o[62725] = i[122];
  assign o[62726] = i[122];
  assign o[62727] = i[122];
  assign o[62728] = i[122];
  assign o[62729] = i[122];
  assign o[62730] = i[122];
  assign o[62731] = i[122];
  assign o[62732] = i[122];
  assign o[62733] = i[122];
  assign o[62734] = i[122];
  assign o[62735] = i[122];
  assign o[62736] = i[122];
  assign o[62737] = i[122];
  assign o[62738] = i[122];
  assign o[62739] = i[122];
  assign o[62740] = i[122];
  assign o[62741] = i[122];
  assign o[62742] = i[122];
  assign o[62743] = i[122];
  assign o[62744] = i[122];
  assign o[62745] = i[122];
  assign o[62746] = i[122];
  assign o[62747] = i[122];
  assign o[62748] = i[122];
  assign o[62749] = i[122];
  assign o[62750] = i[122];
  assign o[62751] = i[122];
  assign o[62752] = i[122];
  assign o[62753] = i[122];
  assign o[62754] = i[122];
  assign o[62755] = i[122];
  assign o[62756] = i[122];
  assign o[62757] = i[122];
  assign o[62758] = i[122];
  assign o[62759] = i[122];
  assign o[62760] = i[122];
  assign o[62761] = i[122];
  assign o[62762] = i[122];
  assign o[62763] = i[122];
  assign o[62764] = i[122];
  assign o[62765] = i[122];
  assign o[62766] = i[122];
  assign o[62767] = i[122];
  assign o[62768] = i[122];
  assign o[62769] = i[122];
  assign o[62770] = i[122];
  assign o[62771] = i[122];
  assign o[62772] = i[122];
  assign o[62773] = i[122];
  assign o[62774] = i[122];
  assign o[62775] = i[122];
  assign o[62776] = i[122];
  assign o[62777] = i[122];
  assign o[62778] = i[122];
  assign o[62779] = i[122];
  assign o[62780] = i[122];
  assign o[62781] = i[122];
  assign o[62782] = i[122];
  assign o[62783] = i[122];
  assign o[62784] = i[122];
  assign o[62785] = i[122];
  assign o[62786] = i[122];
  assign o[62787] = i[122];
  assign o[62788] = i[122];
  assign o[62789] = i[122];
  assign o[62790] = i[122];
  assign o[62791] = i[122];
  assign o[62792] = i[122];
  assign o[62793] = i[122];
  assign o[62794] = i[122];
  assign o[62795] = i[122];
  assign o[62796] = i[122];
  assign o[62797] = i[122];
  assign o[62798] = i[122];
  assign o[62799] = i[122];
  assign o[62800] = i[122];
  assign o[62801] = i[122];
  assign o[62802] = i[122];
  assign o[62803] = i[122];
  assign o[62804] = i[122];
  assign o[62805] = i[122];
  assign o[62806] = i[122];
  assign o[62807] = i[122];
  assign o[62808] = i[122];
  assign o[62809] = i[122];
  assign o[62810] = i[122];
  assign o[62811] = i[122];
  assign o[62812] = i[122];
  assign o[62813] = i[122];
  assign o[62814] = i[122];
  assign o[62815] = i[122];
  assign o[62816] = i[122];
  assign o[62817] = i[122];
  assign o[62818] = i[122];
  assign o[62819] = i[122];
  assign o[62820] = i[122];
  assign o[62821] = i[122];
  assign o[62822] = i[122];
  assign o[62823] = i[122];
  assign o[62824] = i[122];
  assign o[62825] = i[122];
  assign o[62826] = i[122];
  assign o[62827] = i[122];
  assign o[62828] = i[122];
  assign o[62829] = i[122];
  assign o[62830] = i[122];
  assign o[62831] = i[122];
  assign o[62832] = i[122];
  assign o[62833] = i[122];
  assign o[62834] = i[122];
  assign o[62835] = i[122];
  assign o[62836] = i[122];
  assign o[62837] = i[122];
  assign o[62838] = i[122];
  assign o[62839] = i[122];
  assign o[62840] = i[122];
  assign o[62841] = i[122];
  assign o[62842] = i[122];
  assign o[62843] = i[122];
  assign o[62844] = i[122];
  assign o[62845] = i[122];
  assign o[62846] = i[122];
  assign o[62847] = i[122];
  assign o[62848] = i[122];
  assign o[62849] = i[122];
  assign o[62850] = i[122];
  assign o[62851] = i[122];
  assign o[62852] = i[122];
  assign o[62853] = i[122];
  assign o[62854] = i[122];
  assign o[62855] = i[122];
  assign o[62856] = i[122];
  assign o[62857] = i[122];
  assign o[62858] = i[122];
  assign o[62859] = i[122];
  assign o[62860] = i[122];
  assign o[62861] = i[122];
  assign o[62862] = i[122];
  assign o[62863] = i[122];
  assign o[62864] = i[122];
  assign o[62865] = i[122];
  assign o[62866] = i[122];
  assign o[62867] = i[122];
  assign o[62868] = i[122];
  assign o[62869] = i[122];
  assign o[62870] = i[122];
  assign o[62871] = i[122];
  assign o[62872] = i[122];
  assign o[62873] = i[122];
  assign o[62874] = i[122];
  assign o[62875] = i[122];
  assign o[62876] = i[122];
  assign o[62877] = i[122];
  assign o[62878] = i[122];
  assign o[62879] = i[122];
  assign o[62880] = i[122];
  assign o[62881] = i[122];
  assign o[62882] = i[122];
  assign o[62883] = i[122];
  assign o[62884] = i[122];
  assign o[62885] = i[122];
  assign o[62886] = i[122];
  assign o[62887] = i[122];
  assign o[62888] = i[122];
  assign o[62889] = i[122];
  assign o[62890] = i[122];
  assign o[62891] = i[122];
  assign o[62892] = i[122];
  assign o[62893] = i[122];
  assign o[62894] = i[122];
  assign o[62895] = i[122];
  assign o[62896] = i[122];
  assign o[62897] = i[122];
  assign o[62898] = i[122];
  assign o[62899] = i[122];
  assign o[62900] = i[122];
  assign o[62901] = i[122];
  assign o[62902] = i[122];
  assign o[62903] = i[122];
  assign o[62904] = i[122];
  assign o[62905] = i[122];
  assign o[62906] = i[122];
  assign o[62907] = i[122];
  assign o[62908] = i[122];
  assign o[62909] = i[122];
  assign o[62910] = i[122];
  assign o[62911] = i[122];
  assign o[62912] = i[122];
  assign o[62913] = i[122];
  assign o[62914] = i[122];
  assign o[62915] = i[122];
  assign o[62916] = i[122];
  assign o[62917] = i[122];
  assign o[62918] = i[122];
  assign o[62919] = i[122];
  assign o[62920] = i[122];
  assign o[62921] = i[122];
  assign o[62922] = i[122];
  assign o[62923] = i[122];
  assign o[62924] = i[122];
  assign o[62925] = i[122];
  assign o[62926] = i[122];
  assign o[62927] = i[122];
  assign o[62928] = i[122];
  assign o[62929] = i[122];
  assign o[62930] = i[122];
  assign o[62931] = i[122];
  assign o[62932] = i[122];
  assign o[62933] = i[122];
  assign o[62934] = i[122];
  assign o[62935] = i[122];
  assign o[62936] = i[122];
  assign o[62937] = i[122];
  assign o[62938] = i[122];
  assign o[62939] = i[122];
  assign o[62940] = i[122];
  assign o[62941] = i[122];
  assign o[62942] = i[122];
  assign o[62943] = i[122];
  assign o[62944] = i[122];
  assign o[62945] = i[122];
  assign o[62946] = i[122];
  assign o[62947] = i[122];
  assign o[62948] = i[122];
  assign o[62949] = i[122];
  assign o[62950] = i[122];
  assign o[62951] = i[122];
  assign o[62952] = i[122];
  assign o[62953] = i[122];
  assign o[62954] = i[122];
  assign o[62955] = i[122];
  assign o[62956] = i[122];
  assign o[62957] = i[122];
  assign o[62958] = i[122];
  assign o[62959] = i[122];
  assign o[62960] = i[122];
  assign o[62961] = i[122];
  assign o[62962] = i[122];
  assign o[62963] = i[122];
  assign o[62964] = i[122];
  assign o[62965] = i[122];
  assign o[62966] = i[122];
  assign o[62967] = i[122];
  assign o[62968] = i[122];
  assign o[62969] = i[122];
  assign o[62970] = i[122];
  assign o[62971] = i[122];
  assign o[62972] = i[122];
  assign o[62973] = i[122];
  assign o[62974] = i[122];
  assign o[62975] = i[122];
  assign o[61952] = i[121];
  assign o[61953] = i[121];
  assign o[61954] = i[121];
  assign o[61955] = i[121];
  assign o[61956] = i[121];
  assign o[61957] = i[121];
  assign o[61958] = i[121];
  assign o[61959] = i[121];
  assign o[61960] = i[121];
  assign o[61961] = i[121];
  assign o[61962] = i[121];
  assign o[61963] = i[121];
  assign o[61964] = i[121];
  assign o[61965] = i[121];
  assign o[61966] = i[121];
  assign o[61967] = i[121];
  assign o[61968] = i[121];
  assign o[61969] = i[121];
  assign o[61970] = i[121];
  assign o[61971] = i[121];
  assign o[61972] = i[121];
  assign o[61973] = i[121];
  assign o[61974] = i[121];
  assign o[61975] = i[121];
  assign o[61976] = i[121];
  assign o[61977] = i[121];
  assign o[61978] = i[121];
  assign o[61979] = i[121];
  assign o[61980] = i[121];
  assign o[61981] = i[121];
  assign o[61982] = i[121];
  assign o[61983] = i[121];
  assign o[61984] = i[121];
  assign o[61985] = i[121];
  assign o[61986] = i[121];
  assign o[61987] = i[121];
  assign o[61988] = i[121];
  assign o[61989] = i[121];
  assign o[61990] = i[121];
  assign o[61991] = i[121];
  assign o[61992] = i[121];
  assign o[61993] = i[121];
  assign o[61994] = i[121];
  assign o[61995] = i[121];
  assign o[61996] = i[121];
  assign o[61997] = i[121];
  assign o[61998] = i[121];
  assign o[61999] = i[121];
  assign o[62000] = i[121];
  assign o[62001] = i[121];
  assign o[62002] = i[121];
  assign o[62003] = i[121];
  assign o[62004] = i[121];
  assign o[62005] = i[121];
  assign o[62006] = i[121];
  assign o[62007] = i[121];
  assign o[62008] = i[121];
  assign o[62009] = i[121];
  assign o[62010] = i[121];
  assign o[62011] = i[121];
  assign o[62012] = i[121];
  assign o[62013] = i[121];
  assign o[62014] = i[121];
  assign o[62015] = i[121];
  assign o[62016] = i[121];
  assign o[62017] = i[121];
  assign o[62018] = i[121];
  assign o[62019] = i[121];
  assign o[62020] = i[121];
  assign o[62021] = i[121];
  assign o[62022] = i[121];
  assign o[62023] = i[121];
  assign o[62024] = i[121];
  assign o[62025] = i[121];
  assign o[62026] = i[121];
  assign o[62027] = i[121];
  assign o[62028] = i[121];
  assign o[62029] = i[121];
  assign o[62030] = i[121];
  assign o[62031] = i[121];
  assign o[62032] = i[121];
  assign o[62033] = i[121];
  assign o[62034] = i[121];
  assign o[62035] = i[121];
  assign o[62036] = i[121];
  assign o[62037] = i[121];
  assign o[62038] = i[121];
  assign o[62039] = i[121];
  assign o[62040] = i[121];
  assign o[62041] = i[121];
  assign o[62042] = i[121];
  assign o[62043] = i[121];
  assign o[62044] = i[121];
  assign o[62045] = i[121];
  assign o[62046] = i[121];
  assign o[62047] = i[121];
  assign o[62048] = i[121];
  assign o[62049] = i[121];
  assign o[62050] = i[121];
  assign o[62051] = i[121];
  assign o[62052] = i[121];
  assign o[62053] = i[121];
  assign o[62054] = i[121];
  assign o[62055] = i[121];
  assign o[62056] = i[121];
  assign o[62057] = i[121];
  assign o[62058] = i[121];
  assign o[62059] = i[121];
  assign o[62060] = i[121];
  assign o[62061] = i[121];
  assign o[62062] = i[121];
  assign o[62063] = i[121];
  assign o[62064] = i[121];
  assign o[62065] = i[121];
  assign o[62066] = i[121];
  assign o[62067] = i[121];
  assign o[62068] = i[121];
  assign o[62069] = i[121];
  assign o[62070] = i[121];
  assign o[62071] = i[121];
  assign o[62072] = i[121];
  assign o[62073] = i[121];
  assign o[62074] = i[121];
  assign o[62075] = i[121];
  assign o[62076] = i[121];
  assign o[62077] = i[121];
  assign o[62078] = i[121];
  assign o[62079] = i[121];
  assign o[62080] = i[121];
  assign o[62081] = i[121];
  assign o[62082] = i[121];
  assign o[62083] = i[121];
  assign o[62084] = i[121];
  assign o[62085] = i[121];
  assign o[62086] = i[121];
  assign o[62087] = i[121];
  assign o[62088] = i[121];
  assign o[62089] = i[121];
  assign o[62090] = i[121];
  assign o[62091] = i[121];
  assign o[62092] = i[121];
  assign o[62093] = i[121];
  assign o[62094] = i[121];
  assign o[62095] = i[121];
  assign o[62096] = i[121];
  assign o[62097] = i[121];
  assign o[62098] = i[121];
  assign o[62099] = i[121];
  assign o[62100] = i[121];
  assign o[62101] = i[121];
  assign o[62102] = i[121];
  assign o[62103] = i[121];
  assign o[62104] = i[121];
  assign o[62105] = i[121];
  assign o[62106] = i[121];
  assign o[62107] = i[121];
  assign o[62108] = i[121];
  assign o[62109] = i[121];
  assign o[62110] = i[121];
  assign o[62111] = i[121];
  assign o[62112] = i[121];
  assign o[62113] = i[121];
  assign o[62114] = i[121];
  assign o[62115] = i[121];
  assign o[62116] = i[121];
  assign o[62117] = i[121];
  assign o[62118] = i[121];
  assign o[62119] = i[121];
  assign o[62120] = i[121];
  assign o[62121] = i[121];
  assign o[62122] = i[121];
  assign o[62123] = i[121];
  assign o[62124] = i[121];
  assign o[62125] = i[121];
  assign o[62126] = i[121];
  assign o[62127] = i[121];
  assign o[62128] = i[121];
  assign o[62129] = i[121];
  assign o[62130] = i[121];
  assign o[62131] = i[121];
  assign o[62132] = i[121];
  assign o[62133] = i[121];
  assign o[62134] = i[121];
  assign o[62135] = i[121];
  assign o[62136] = i[121];
  assign o[62137] = i[121];
  assign o[62138] = i[121];
  assign o[62139] = i[121];
  assign o[62140] = i[121];
  assign o[62141] = i[121];
  assign o[62142] = i[121];
  assign o[62143] = i[121];
  assign o[62144] = i[121];
  assign o[62145] = i[121];
  assign o[62146] = i[121];
  assign o[62147] = i[121];
  assign o[62148] = i[121];
  assign o[62149] = i[121];
  assign o[62150] = i[121];
  assign o[62151] = i[121];
  assign o[62152] = i[121];
  assign o[62153] = i[121];
  assign o[62154] = i[121];
  assign o[62155] = i[121];
  assign o[62156] = i[121];
  assign o[62157] = i[121];
  assign o[62158] = i[121];
  assign o[62159] = i[121];
  assign o[62160] = i[121];
  assign o[62161] = i[121];
  assign o[62162] = i[121];
  assign o[62163] = i[121];
  assign o[62164] = i[121];
  assign o[62165] = i[121];
  assign o[62166] = i[121];
  assign o[62167] = i[121];
  assign o[62168] = i[121];
  assign o[62169] = i[121];
  assign o[62170] = i[121];
  assign o[62171] = i[121];
  assign o[62172] = i[121];
  assign o[62173] = i[121];
  assign o[62174] = i[121];
  assign o[62175] = i[121];
  assign o[62176] = i[121];
  assign o[62177] = i[121];
  assign o[62178] = i[121];
  assign o[62179] = i[121];
  assign o[62180] = i[121];
  assign o[62181] = i[121];
  assign o[62182] = i[121];
  assign o[62183] = i[121];
  assign o[62184] = i[121];
  assign o[62185] = i[121];
  assign o[62186] = i[121];
  assign o[62187] = i[121];
  assign o[62188] = i[121];
  assign o[62189] = i[121];
  assign o[62190] = i[121];
  assign o[62191] = i[121];
  assign o[62192] = i[121];
  assign o[62193] = i[121];
  assign o[62194] = i[121];
  assign o[62195] = i[121];
  assign o[62196] = i[121];
  assign o[62197] = i[121];
  assign o[62198] = i[121];
  assign o[62199] = i[121];
  assign o[62200] = i[121];
  assign o[62201] = i[121];
  assign o[62202] = i[121];
  assign o[62203] = i[121];
  assign o[62204] = i[121];
  assign o[62205] = i[121];
  assign o[62206] = i[121];
  assign o[62207] = i[121];
  assign o[62208] = i[121];
  assign o[62209] = i[121];
  assign o[62210] = i[121];
  assign o[62211] = i[121];
  assign o[62212] = i[121];
  assign o[62213] = i[121];
  assign o[62214] = i[121];
  assign o[62215] = i[121];
  assign o[62216] = i[121];
  assign o[62217] = i[121];
  assign o[62218] = i[121];
  assign o[62219] = i[121];
  assign o[62220] = i[121];
  assign o[62221] = i[121];
  assign o[62222] = i[121];
  assign o[62223] = i[121];
  assign o[62224] = i[121];
  assign o[62225] = i[121];
  assign o[62226] = i[121];
  assign o[62227] = i[121];
  assign o[62228] = i[121];
  assign o[62229] = i[121];
  assign o[62230] = i[121];
  assign o[62231] = i[121];
  assign o[62232] = i[121];
  assign o[62233] = i[121];
  assign o[62234] = i[121];
  assign o[62235] = i[121];
  assign o[62236] = i[121];
  assign o[62237] = i[121];
  assign o[62238] = i[121];
  assign o[62239] = i[121];
  assign o[62240] = i[121];
  assign o[62241] = i[121];
  assign o[62242] = i[121];
  assign o[62243] = i[121];
  assign o[62244] = i[121];
  assign o[62245] = i[121];
  assign o[62246] = i[121];
  assign o[62247] = i[121];
  assign o[62248] = i[121];
  assign o[62249] = i[121];
  assign o[62250] = i[121];
  assign o[62251] = i[121];
  assign o[62252] = i[121];
  assign o[62253] = i[121];
  assign o[62254] = i[121];
  assign o[62255] = i[121];
  assign o[62256] = i[121];
  assign o[62257] = i[121];
  assign o[62258] = i[121];
  assign o[62259] = i[121];
  assign o[62260] = i[121];
  assign o[62261] = i[121];
  assign o[62262] = i[121];
  assign o[62263] = i[121];
  assign o[62264] = i[121];
  assign o[62265] = i[121];
  assign o[62266] = i[121];
  assign o[62267] = i[121];
  assign o[62268] = i[121];
  assign o[62269] = i[121];
  assign o[62270] = i[121];
  assign o[62271] = i[121];
  assign o[62272] = i[121];
  assign o[62273] = i[121];
  assign o[62274] = i[121];
  assign o[62275] = i[121];
  assign o[62276] = i[121];
  assign o[62277] = i[121];
  assign o[62278] = i[121];
  assign o[62279] = i[121];
  assign o[62280] = i[121];
  assign o[62281] = i[121];
  assign o[62282] = i[121];
  assign o[62283] = i[121];
  assign o[62284] = i[121];
  assign o[62285] = i[121];
  assign o[62286] = i[121];
  assign o[62287] = i[121];
  assign o[62288] = i[121];
  assign o[62289] = i[121];
  assign o[62290] = i[121];
  assign o[62291] = i[121];
  assign o[62292] = i[121];
  assign o[62293] = i[121];
  assign o[62294] = i[121];
  assign o[62295] = i[121];
  assign o[62296] = i[121];
  assign o[62297] = i[121];
  assign o[62298] = i[121];
  assign o[62299] = i[121];
  assign o[62300] = i[121];
  assign o[62301] = i[121];
  assign o[62302] = i[121];
  assign o[62303] = i[121];
  assign o[62304] = i[121];
  assign o[62305] = i[121];
  assign o[62306] = i[121];
  assign o[62307] = i[121];
  assign o[62308] = i[121];
  assign o[62309] = i[121];
  assign o[62310] = i[121];
  assign o[62311] = i[121];
  assign o[62312] = i[121];
  assign o[62313] = i[121];
  assign o[62314] = i[121];
  assign o[62315] = i[121];
  assign o[62316] = i[121];
  assign o[62317] = i[121];
  assign o[62318] = i[121];
  assign o[62319] = i[121];
  assign o[62320] = i[121];
  assign o[62321] = i[121];
  assign o[62322] = i[121];
  assign o[62323] = i[121];
  assign o[62324] = i[121];
  assign o[62325] = i[121];
  assign o[62326] = i[121];
  assign o[62327] = i[121];
  assign o[62328] = i[121];
  assign o[62329] = i[121];
  assign o[62330] = i[121];
  assign o[62331] = i[121];
  assign o[62332] = i[121];
  assign o[62333] = i[121];
  assign o[62334] = i[121];
  assign o[62335] = i[121];
  assign o[62336] = i[121];
  assign o[62337] = i[121];
  assign o[62338] = i[121];
  assign o[62339] = i[121];
  assign o[62340] = i[121];
  assign o[62341] = i[121];
  assign o[62342] = i[121];
  assign o[62343] = i[121];
  assign o[62344] = i[121];
  assign o[62345] = i[121];
  assign o[62346] = i[121];
  assign o[62347] = i[121];
  assign o[62348] = i[121];
  assign o[62349] = i[121];
  assign o[62350] = i[121];
  assign o[62351] = i[121];
  assign o[62352] = i[121];
  assign o[62353] = i[121];
  assign o[62354] = i[121];
  assign o[62355] = i[121];
  assign o[62356] = i[121];
  assign o[62357] = i[121];
  assign o[62358] = i[121];
  assign o[62359] = i[121];
  assign o[62360] = i[121];
  assign o[62361] = i[121];
  assign o[62362] = i[121];
  assign o[62363] = i[121];
  assign o[62364] = i[121];
  assign o[62365] = i[121];
  assign o[62366] = i[121];
  assign o[62367] = i[121];
  assign o[62368] = i[121];
  assign o[62369] = i[121];
  assign o[62370] = i[121];
  assign o[62371] = i[121];
  assign o[62372] = i[121];
  assign o[62373] = i[121];
  assign o[62374] = i[121];
  assign o[62375] = i[121];
  assign o[62376] = i[121];
  assign o[62377] = i[121];
  assign o[62378] = i[121];
  assign o[62379] = i[121];
  assign o[62380] = i[121];
  assign o[62381] = i[121];
  assign o[62382] = i[121];
  assign o[62383] = i[121];
  assign o[62384] = i[121];
  assign o[62385] = i[121];
  assign o[62386] = i[121];
  assign o[62387] = i[121];
  assign o[62388] = i[121];
  assign o[62389] = i[121];
  assign o[62390] = i[121];
  assign o[62391] = i[121];
  assign o[62392] = i[121];
  assign o[62393] = i[121];
  assign o[62394] = i[121];
  assign o[62395] = i[121];
  assign o[62396] = i[121];
  assign o[62397] = i[121];
  assign o[62398] = i[121];
  assign o[62399] = i[121];
  assign o[62400] = i[121];
  assign o[62401] = i[121];
  assign o[62402] = i[121];
  assign o[62403] = i[121];
  assign o[62404] = i[121];
  assign o[62405] = i[121];
  assign o[62406] = i[121];
  assign o[62407] = i[121];
  assign o[62408] = i[121];
  assign o[62409] = i[121];
  assign o[62410] = i[121];
  assign o[62411] = i[121];
  assign o[62412] = i[121];
  assign o[62413] = i[121];
  assign o[62414] = i[121];
  assign o[62415] = i[121];
  assign o[62416] = i[121];
  assign o[62417] = i[121];
  assign o[62418] = i[121];
  assign o[62419] = i[121];
  assign o[62420] = i[121];
  assign o[62421] = i[121];
  assign o[62422] = i[121];
  assign o[62423] = i[121];
  assign o[62424] = i[121];
  assign o[62425] = i[121];
  assign o[62426] = i[121];
  assign o[62427] = i[121];
  assign o[62428] = i[121];
  assign o[62429] = i[121];
  assign o[62430] = i[121];
  assign o[62431] = i[121];
  assign o[62432] = i[121];
  assign o[62433] = i[121];
  assign o[62434] = i[121];
  assign o[62435] = i[121];
  assign o[62436] = i[121];
  assign o[62437] = i[121];
  assign o[62438] = i[121];
  assign o[62439] = i[121];
  assign o[62440] = i[121];
  assign o[62441] = i[121];
  assign o[62442] = i[121];
  assign o[62443] = i[121];
  assign o[62444] = i[121];
  assign o[62445] = i[121];
  assign o[62446] = i[121];
  assign o[62447] = i[121];
  assign o[62448] = i[121];
  assign o[62449] = i[121];
  assign o[62450] = i[121];
  assign o[62451] = i[121];
  assign o[62452] = i[121];
  assign o[62453] = i[121];
  assign o[62454] = i[121];
  assign o[62455] = i[121];
  assign o[62456] = i[121];
  assign o[62457] = i[121];
  assign o[62458] = i[121];
  assign o[62459] = i[121];
  assign o[62460] = i[121];
  assign o[62461] = i[121];
  assign o[62462] = i[121];
  assign o[62463] = i[121];
  assign o[61440] = i[120];
  assign o[61441] = i[120];
  assign o[61442] = i[120];
  assign o[61443] = i[120];
  assign o[61444] = i[120];
  assign o[61445] = i[120];
  assign o[61446] = i[120];
  assign o[61447] = i[120];
  assign o[61448] = i[120];
  assign o[61449] = i[120];
  assign o[61450] = i[120];
  assign o[61451] = i[120];
  assign o[61452] = i[120];
  assign o[61453] = i[120];
  assign o[61454] = i[120];
  assign o[61455] = i[120];
  assign o[61456] = i[120];
  assign o[61457] = i[120];
  assign o[61458] = i[120];
  assign o[61459] = i[120];
  assign o[61460] = i[120];
  assign o[61461] = i[120];
  assign o[61462] = i[120];
  assign o[61463] = i[120];
  assign o[61464] = i[120];
  assign o[61465] = i[120];
  assign o[61466] = i[120];
  assign o[61467] = i[120];
  assign o[61468] = i[120];
  assign o[61469] = i[120];
  assign o[61470] = i[120];
  assign o[61471] = i[120];
  assign o[61472] = i[120];
  assign o[61473] = i[120];
  assign o[61474] = i[120];
  assign o[61475] = i[120];
  assign o[61476] = i[120];
  assign o[61477] = i[120];
  assign o[61478] = i[120];
  assign o[61479] = i[120];
  assign o[61480] = i[120];
  assign o[61481] = i[120];
  assign o[61482] = i[120];
  assign o[61483] = i[120];
  assign o[61484] = i[120];
  assign o[61485] = i[120];
  assign o[61486] = i[120];
  assign o[61487] = i[120];
  assign o[61488] = i[120];
  assign o[61489] = i[120];
  assign o[61490] = i[120];
  assign o[61491] = i[120];
  assign o[61492] = i[120];
  assign o[61493] = i[120];
  assign o[61494] = i[120];
  assign o[61495] = i[120];
  assign o[61496] = i[120];
  assign o[61497] = i[120];
  assign o[61498] = i[120];
  assign o[61499] = i[120];
  assign o[61500] = i[120];
  assign o[61501] = i[120];
  assign o[61502] = i[120];
  assign o[61503] = i[120];
  assign o[61504] = i[120];
  assign o[61505] = i[120];
  assign o[61506] = i[120];
  assign o[61507] = i[120];
  assign o[61508] = i[120];
  assign o[61509] = i[120];
  assign o[61510] = i[120];
  assign o[61511] = i[120];
  assign o[61512] = i[120];
  assign o[61513] = i[120];
  assign o[61514] = i[120];
  assign o[61515] = i[120];
  assign o[61516] = i[120];
  assign o[61517] = i[120];
  assign o[61518] = i[120];
  assign o[61519] = i[120];
  assign o[61520] = i[120];
  assign o[61521] = i[120];
  assign o[61522] = i[120];
  assign o[61523] = i[120];
  assign o[61524] = i[120];
  assign o[61525] = i[120];
  assign o[61526] = i[120];
  assign o[61527] = i[120];
  assign o[61528] = i[120];
  assign o[61529] = i[120];
  assign o[61530] = i[120];
  assign o[61531] = i[120];
  assign o[61532] = i[120];
  assign o[61533] = i[120];
  assign o[61534] = i[120];
  assign o[61535] = i[120];
  assign o[61536] = i[120];
  assign o[61537] = i[120];
  assign o[61538] = i[120];
  assign o[61539] = i[120];
  assign o[61540] = i[120];
  assign o[61541] = i[120];
  assign o[61542] = i[120];
  assign o[61543] = i[120];
  assign o[61544] = i[120];
  assign o[61545] = i[120];
  assign o[61546] = i[120];
  assign o[61547] = i[120];
  assign o[61548] = i[120];
  assign o[61549] = i[120];
  assign o[61550] = i[120];
  assign o[61551] = i[120];
  assign o[61552] = i[120];
  assign o[61553] = i[120];
  assign o[61554] = i[120];
  assign o[61555] = i[120];
  assign o[61556] = i[120];
  assign o[61557] = i[120];
  assign o[61558] = i[120];
  assign o[61559] = i[120];
  assign o[61560] = i[120];
  assign o[61561] = i[120];
  assign o[61562] = i[120];
  assign o[61563] = i[120];
  assign o[61564] = i[120];
  assign o[61565] = i[120];
  assign o[61566] = i[120];
  assign o[61567] = i[120];
  assign o[61568] = i[120];
  assign o[61569] = i[120];
  assign o[61570] = i[120];
  assign o[61571] = i[120];
  assign o[61572] = i[120];
  assign o[61573] = i[120];
  assign o[61574] = i[120];
  assign o[61575] = i[120];
  assign o[61576] = i[120];
  assign o[61577] = i[120];
  assign o[61578] = i[120];
  assign o[61579] = i[120];
  assign o[61580] = i[120];
  assign o[61581] = i[120];
  assign o[61582] = i[120];
  assign o[61583] = i[120];
  assign o[61584] = i[120];
  assign o[61585] = i[120];
  assign o[61586] = i[120];
  assign o[61587] = i[120];
  assign o[61588] = i[120];
  assign o[61589] = i[120];
  assign o[61590] = i[120];
  assign o[61591] = i[120];
  assign o[61592] = i[120];
  assign o[61593] = i[120];
  assign o[61594] = i[120];
  assign o[61595] = i[120];
  assign o[61596] = i[120];
  assign o[61597] = i[120];
  assign o[61598] = i[120];
  assign o[61599] = i[120];
  assign o[61600] = i[120];
  assign o[61601] = i[120];
  assign o[61602] = i[120];
  assign o[61603] = i[120];
  assign o[61604] = i[120];
  assign o[61605] = i[120];
  assign o[61606] = i[120];
  assign o[61607] = i[120];
  assign o[61608] = i[120];
  assign o[61609] = i[120];
  assign o[61610] = i[120];
  assign o[61611] = i[120];
  assign o[61612] = i[120];
  assign o[61613] = i[120];
  assign o[61614] = i[120];
  assign o[61615] = i[120];
  assign o[61616] = i[120];
  assign o[61617] = i[120];
  assign o[61618] = i[120];
  assign o[61619] = i[120];
  assign o[61620] = i[120];
  assign o[61621] = i[120];
  assign o[61622] = i[120];
  assign o[61623] = i[120];
  assign o[61624] = i[120];
  assign o[61625] = i[120];
  assign o[61626] = i[120];
  assign o[61627] = i[120];
  assign o[61628] = i[120];
  assign o[61629] = i[120];
  assign o[61630] = i[120];
  assign o[61631] = i[120];
  assign o[61632] = i[120];
  assign o[61633] = i[120];
  assign o[61634] = i[120];
  assign o[61635] = i[120];
  assign o[61636] = i[120];
  assign o[61637] = i[120];
  assign o[61638] = i[120];
  assign o[61639] = i[120];
  assign o[61640] = i[120];
  assign o[61641] = i[120];
  assign o[61642] = i[120];
  assign o[61643] = i[120];
  assign o[61644] = i[120];
  assign o[61645] = i[120];
  assign o[61646] = i[120];
  assign o[61647] = i[120];
  assign o[61648] = i[120];
  assign o[61649] = i[120];
  assign o[61650] = i[120];
  assign o[61651] = i[120];
  assign o[61652] = i[120];
  assign o[61653] = i[120];
  assign o[61654] = i[120];
  assign o[61655] = i[120];
  assign o[61656] = i[120];
  assign o[61657] = i[120];
  assign o[61658] = i[120];
  assign o[61659] = i[120];
  assign o[61660] = i[120];
  assign o[61661] = i[120];
  assign o[61662] = i[120];
  assign o[61663] = i[120];
  assign o[61664] = i[120];
  assign o[61665] = i[120];
  assign o[61666] = i[120];
  assign o[61667] = i[120];
  assign o[61668] = i[120];
  assign o[61669] = i[120];
  assign o[61670] = i[120];
  assign o[61671] = i[120];
  assign o[61672] = i[120];
  assign o[61673] = i[120];
  assign o[61674] = i[120];
  assign o[61675] = i[120];
  assign o[61676] = i[120];
  assign o[61677] = i[120];
  assign o[61678] = i[120];
  assign o[61679] = i[120];
  assign o[61680] = i[120];
  assign o[61681] = i[120];
  assign o[61682] = i[120];
  assign o[61683] = i[120];
  assign o[61684] = i[120];
  assign o[61685] = i[120];
  assign o[61686] = i[120];
  assign o[61687] = i[120];
  assign o[61688] = i[120];
  assign o[61689] = i[120];
  assign o[61690] = i[120];
  assign o[61691] = i[120];
  assign o[61692] = i[120];
  assign o[61693] = i[120];
  assign o[61694] = i[120];
  assign o[61695] = i[120];
  assign o[61696] = i[120];
  assign o[61697] = i[120];
  assign o[61698] = i[120];
  assign o[61699] = i[120];
  assign o[61700] = i[120];
  assign o[61701] = i[120];
  assign o[61702] = i[120];
  assign o[61703] = i[120];
  assign o[61704] = i[120];
  assign o[61705] = i[120];
  assign o[61706] = i[120];
  assign o[61707] = i[120];
  assign o[61708] = i[120];
  assign o[61709] = i[120];
  assign o[61710] = i[120];
  assign o[61711] = i[120];
  assign o[61712] = i[120];
  assign o[61713] = i[120];
  assign o[61714] = i[120];
  assign o[61715] = i[120];
  assign o[61716] = i[120];
  assign o[61717] = i[120];
  assign o[61718] = i[120];
  assign o[61719] = i[120];
  assign o[61720] = i[120];
  assign o[61721] = i[120];
  assign o[61722] = i[120];
  assign o[61723] = i[120];
  assign o[61724] = i[120];
  assign o[61725] = i[120];
  assign o[61726] = i[120];
  assign o[61727] = i[120];
  assign o[61728] = i[120];
  assign o[61729] = i[120];
  assign o[61730] = i[120];
  assign o[61731] = i[120];
  assign o[61732] = i[120];
  assign o[61733] = i[120];
  assign o[61734] = i[120];
  assign o[61735] = i[120];
  assign o[61736] = i[120];
  assign o[61737] = i[120];
  assign o[61738] = i[120];
  assign o[61739] = i[120];
  assign o[61740] = i[120];
  assign o[61741] = i[120];
  assign o[61742] = i[120];
  assign o[61743] = i[120];
  assign o[61744] = i[120];
  assign o[61745] = i[120];
  assign o[61746] = i[120];
  assign o[61747] = i[120];
  assign o[61748] = i[120];
  assign o[61749] = i[120];
  assign o[61750] = i[120];
  assign o[61751] = i[120];
  assign o[61752] = i[120];
  assign o[61753] = i[120];
  assign o[61754] = i[120];
  assign o[61755] = i[120];
  assign o[61756] = i[120];
  assign o[61757] = i[120];
  assign o[61758] = i[120];
  assign o[61759] = i[120];
  assign o[61760] = i[120];
  assign o[61761] = i[120];
  assign o[61762] = i[120];
  assign o[61763] = i[120];
  assign o[61764] = i[120];
  assign o[61765] = i[120];
  assign o[61766] = i[120];
  assign o[61767] = i[120];
  assign o[61768] = i[120];
  assign o[61769] = i[120];
  assign o[61770] = i[120];
  assign o[61771] = i[120];
  assign o[61772] = i[120];
  assign o[61773] = i[120];
  assign o[61774] = i[120];
  assign o[61775] = i[120];
  assign o[61776] = i[120];
  assign o[61777] = i[120];
  assign o[61778] = i[120];
  assign o[61779] = i[120];
  assign o[61780] = i[120];
  assign o[61781] = i[120];
  assign o[61782] = i[120];
  assign o[61783] = i[120];
  assign o[61784] = i[120];
  assign o[61785] = i[120];
  assign o[61786] = i[120];
  assign o[61787] = i[120];
  assign o[61788] = i[120];
  assign o[61789] = i[120];
  assign o[61790] = i[120];
  assign o[61791] = i[120];
  assign o[61792] = i[120];
  assign o[61793] = i[120];
  assign o[61794] = i[120];
  assign o[61795] = i[120];
  assign o[61796] = i[120];
  assign o[61797] = i[120];
  assign o[61798] = i[120];
  assign o[61799] = i[120];
  assign o[61800] = i[120];
  assign o[61801] = i[120];
  assign o[61802] = i[120];
  assign o[61803] = i[120];
  assign o[61804] = i[120];
  assign o[61805] = i[120];
  assign o[61806] = i[120];
  assign o[61807] = i[120];
  assign o[61808] = i[120];
  assign o[61809] = i[120];
  assign o[61810] = i[120];
  assign o[61811] = i[120];
  assign o[61812] = i[120];
  assign o[61813] = i[120];
  assign o[61814] = i[120];
  assign o[61815] = i[120];
  assign o[61816] = i[120];
  assign o[61817] = i[120];
  assign o[61818] = i[120];
  assign o[61819] = i[120];
  assign o[61820] = i[120];
  assign o[61821] = i[120];
  assign o[61822] = i[120];
  assign o[61823] = i[120];
  assign o[61824] = i[120];
  assign o[61825] = i[120];
  assign o[61826] = i[120];
  assign o[61827] = i[120];
  assign o[61828] = i[120];
  assign o[61829] = i[120];
  assign o[61830] = i[120];
  assign o[61831] = i[120];
  assign o[61832] = i[120];
  assign o[61833] = i[120];
  assign o[61834] = i[120];
  assign o[61835] = i[120];
  assign o[61836] = i[120];
  assign o[61837] = i[120];
  assign o[61838] = i[120];
  assign o[61839] = i[120];
  assign o[61840] = i[120];
  assign o[61841] = i[120];
  assign o[61842] = i[120];
  assign o[61843] = i[120];
  assign o[61844] = i[120];
  assign o[61845] = i[120];
  assign o[61846] = i[120];
  assign o[61847] = i[120];
  assign o[61848] = i[120];
  assign o[61849] = i[120];
  assign o[61850] = i[120];
  assign o[61851] = i[120];
  assign o[61852] = i[120];
  assign o[61853] = i[120];
  assign o[61854] = i[120];
  assign o[61855] = i[120];
  assign o[61856] = i[120];
  assign o[61857] = i[120];
  assign o[61858] = i[120];
  assign o[61859] = i[120];
  assign o[61860] = i[120];
  assign o[61861] = i[120];
  assign o[61862] = i[120];
  assign o[61863] = i[120];
  assign o[61864] = i[120];
  assign o[61865] = i[120];
  assign o[61866] = i[120];
  assign o[61867] = i[120];
  assign o[61868] = i[120];
  assign o[61869] = i[120];
  assign o[61870] = i[120];
  assign o[61871] = i[120];
  assign o[61872] = i[120];
  assign o[61873] = i[120];
  assign o[61874] = i[120];
  assign o[61875] = i[120];
  assign o[61876] = i[120];
  assign o[61877] = i[120];
  assign o[61878] = i[120];
  assign o[61879] = i[120];
  assign o[61880] = i[120];
  assign o[61881] = i[120];
  assign o[61882] = i[120];
  assign o[61883] = i[120];
  assign o[61884] = i[120];
  assign o[61885] = i[120];
  assign o[61886] = i[120];
  assign o[61887] = i[120];
  assign o[61888] = i[120];
  assign o[61889] = i[120];
  assign o[61890] = i[120];
  assign o[61891] = i[120];
  assign o[61892] = i[120];
  assign o[61893] = i[120];
  assign o[61894] = i[120];
  assign o[61895] = i[120];
  assign o[61896] = i[120];
  assign o[61897] = i[120];
  assign o[61898] = i[120];
  assign o[61899] = i[120];
  assign o[61900] = i[120];
  assign o[61901] = i[120];
  assign o[61902] = i[120];
  assign o[61903] = i[120];
  assign o[61904] = i[120];
  assign o[61905] = i[120];
  assign o[61906] = i[120];
  assign o[61907] = i[120];
  assign o[61908] = i[120];
  assign o[61909] = i[120];
  assign o[61910] = i[120];
  assign o[61911] = i[120];
  assign o[61912] = i[120];
  assign o[61913] = i[120];
  assign o[61914] = i[120];
  assign o[61915] = i[120];
  assign o[61916] = i[120];
  assign o[61917] = i[120];
  assign o[61918] = i[120];
  assign o[61919] = i[120];
  assign o[61920] = i[120];
  assign o[61921] = i[120];
  assign o[61922] = i[120];
  assign o[61923] = i[120];
  assign o[61924] = i[120];
  assign o[61925] = i[120];
  assign o[61926] = i[120];
  assign o[61927] = i[120];
  assign o[61928] = i[120];
  assign o[61929] = i[120];
  assign o[61930] = i[120];
  assign o[61931] = i[120];
  assign o[61932] = i[120];
  assign o[61933] = i[120];
  assign o[61934] = i[120];
  assign o[61935] = i[120];
  assign o[61936] = i[120];
  assign o[61937] = i[120];
  assign o[61938] = i[120];
  assign o[61939] = i[120];
  assign o[61940] = i[120];
  assign o[61941] = i[120];
  assign o[61942] = i[120];
  assign o[61943] = i[120];
  assign o[61944] = i[120];
  assign o[61945] = i[120];
  assign o[61946] = i[120];
  assign o[61947] = i[120];
  assign o[61948] = i[120];
  assign o[61949] = i[120];
  assign o[61950] = i[120];
  assign o[61951] = i[120];
  assign o[60928] = i[119];
  assign o[60929] = i[119];
  assign o[60930] = i[119];
  assign o[60931] = i[119];
  assign o[60932] = i[119];
  assign o[60933] = i[119];
  assign o[60934] = i[119];
  assign o[60935] = i[119];
  assign o[60936] = i[119];
  assign o[60937] = i[119];
  assign o[60938] = i[119];
  assign o[60939] = i[119];
  assign o[60940] = i[119];
  assign o[60941] = i[119];
  assign o[60942] = i[119];
  assign o[60943] = i[119];
  assign o[60944] = i[119];
  assign o[60945] = i[119];
  assign o[60946] = i[119];
  assign o[60947] = i[119];
  assign o[60948] = i[119];
  assign o[60949] = i[119];
  assign o[60950] = i[119];
  assign o[60951] = i[119];
  assign o[60952] = i[119];
  assign o[60953] = i[119];
  assign o[60954] = i[119];
  assign o[60955] = i[119];
  assign o[60956] = i[119];
  assign o[60957] = i[119];
  assign o[60958] = i[119];
  assign o[60959] = i[119];
  assign o[60960] = i[119];
  assign o[60961] = i[119];
  assign o[60962] = i[119];
  assign o[60963] = i[119];
  assign o[60964] = i[119];
  assign o[60965] = i[119];
  assign o[60966] = i[119];
  assign o[60967] = i[119];
  assign o[60968] = i[119];
  assign o[60969] = i[119];
  assign o[60970] = i[119];
  assign o[60971] = i[119];
  assign o[60972] = i[119];
  assign o[60973] = i[119];
  assign o[60974] = i[119];
  assign o[60975] = i[119];
  assign o[60976] = i[119];
  assign o[60977] = i[119];
  assign o[60978] = i[119];
  assign o[60979] = i[119];
  assign o[60980] = i[119];
  assign o[60981] = i[119];
  assign o[60982] = i[119];
  assign o[60983] = i[119];
  assign o[60984] = i[119];
  assign o[60985] = i[119];
  assign o[60986] = i[119];
  assign o[60987] = i[119];
  assign o[60988] = i[119];
  assign o[60989] = i[119];
  assign o[60990] = i[119];
  assign o[60991] = i[119];
  assign o[60992] = i[119];
  assign o[60993] = i[119];
  assign o[60994] = i[119];
  assign o[60995] = i[119];
  assign o[60996] = i[119];
  assign o[60997] = i[119];
  assign o[60998] = i[119];
  assign o[60999] = i[119];
  assign o[61000] = i[119];
  assign o[61001] = i[119];
  assign o[61002] = i[119];
  assign o[61003] = i[119];
  assign o[61004] = i[119];
  assign o[61005] = i[119];
  assign o[61006] = i[119];
  assign o[61007] = i[119];
  assign o[61008] = i[119];
  assign o[61009] = i[119];
  assign o[61010] = i[119];
  assign o[61011] = i[119];
  assign o[61012] = i[119];
  assign o[61013] = i[119];
  assign o[61014] = i[119];
  assign o[61015] = i[119];
  assign o[61016] = i[119];
  assign o[61017] = i[119];
  assign o[61018] = i[119];
  assign o[61019] = i[119];
  assign o[61020] = i[119];
  assign o[61021] = i[119];
  assign o[61022] = i[119];
  assign o[61023] = i[119];
  assign o[61024] = i[119];
  assign o[61025] = i[119];
  assign o[61026] = i[119];
  assign o[61027] = i[119];
  assign o[61028] = i[119];
  assign o[61029] = i[119];
  assign o[61030] = i[119];
  assign o[61031] = i[119];
  assign o[61032] = i[119];
  assign o[61033] = i[119];
  assign o[61034] = i[119];
  assign o[61035] = i[119];
  assign o[61036] = i[119];
  assign o[61037] = i[119];
  assign o[61038] = i[119];
  assign o[61039] = i[119];
  assign o[61040] = i[119];
  assign o[61041] = i[119];
  assign o[61042] = i[119];
  assign o[61043] = i[119];
  assign o[61044] = i[119];
  assign o[61045] = i[119];
  assign o[61046] = i[119];
  assign o[61047] = i[119];
  assign o[61048] = i[119];
  assign o[61049] = i[119];
  assign o[61050] = i[119];
  assign o[61051] = i[119];
  assign o[61052] = i[119];
  assign o[61053] = i[119];
  assign o[61054] = i[119];
  assign o[61055] = i[119];
  assign o[61056] = i[119];
  assign o[61057] = i[119];
  assign o[61058] = i[119];
  assign o[61059] = i[119];
  assign o[61060] = i[119];
  assign o[61061] = i[119];
  assign o[61062] = i[119];
  assign o[61063] = i[119];
  assign o[61064] = i[119];
  assign o[61065] = i[119];
  assign o[61066] = i[119];
  assign o[61067] = i[119];
  assign o[61068] = i[119];
  assign o[61069] = i[119];
  assign o[61070] = i[119];
  assign o[61071] = i[119];
  assign o[61072] = i[119];
  assign o[61073] = i[119];
  assign o[61074] = i[119];
  assign o[61075] = i[119];
  assign o[61076] = i[119];
  assign o[61077] = i[119];
  assign o[61078] = i[119];
  assign o[61079] = i[119];
  assign o[61080] = i[119];
  assign o[61081] = i[119];
  assign o[61082] = i[119];
  assign o[61083] = i[119];
  assign o[61084] = i[119];
  assign o[61085] = i[119];
  assign o[61086] = i[119];
  assign o[61087] = i[119];
  assign o[61088] = i[119];
  assign o[61089] = i[119];
  assign o[61090] = i[119];
  assign o[61091] = i[119];
  assign o[61092] = i[119];
  assign o[61093] = i[119];
  assign o[61094] = i[119];
  assign o[61095] = i[119];
  assign o[61096] = i[119];
  assign o[61097] = i[119];
  assign o[61098] = i[119];
  assign o[61099] = i[119];
  assign o[61100] = i[119];
  assign o[61101] = i[119];
  assign o[61102] = i[119];
  assign o[61103] = i[119];
  assign o[61104] = i[119];
  assign o[61105] = i[119];
  assign o[61106] = i[119];
  assign o[61107] = i[119];
  assign o[61108] = i[119];
  assign o[61109] = i[119];
  assign o[61110] = i[119];
  assign o[61111] = i[119];
  assign o[61112] = i[119];
  assign o[61113] = i[119];
  assign o[61114] = i[119];
  assign o[61115] = i[119];
  assign o[61116] = i[119];
  assign o[61117] = i[119];
  assign o[61118] = i[119];
  assign o[61119] = i[119];
  assign o[61120] = i[119];
  assign o[61121] = i[119];
  assign o[61122] = i[119];
  assign o[61123] = i[119];
  assign o[61124] = i[119];
  assign o[61125] = i[119];
  assign o[61126] = i[119];
  assign o[61127] = i[119];
  assign o[61128] = i[119];
  assign o[61129] = i[119];
  assign o[61130] = i[119];
  assign o[61131] = i[119];
  assign o[61132] = i[119];
  assign o[61133] = i[119];
  assign o[61134] = i[119];
  assign o[61135] = i[119];
  assign o[61136] = i[119];
  assign o[61137] = i[119];
  assign o[61138] = i[119];
  assign o[61139] = i[119];
  assign o[61140] = i[119];
  assign o[61141] = i[119];
  assign o[61142] = i[119];
  assign o[61143] = i[119];
  assign o[61144] = i[119];
  assign o[61145] = i[119];
  assign o[61146] = i[119];
  assign o[61147] = i[119];
  assign o[61148] = i[119];
  assign o[61149] = i[119];
  assign o[61150] = i[119];
  assign o[61151] = i[119];
  assign o[61152] = i[119];
  assign o[61153] = i[119];
  assign o[61154] = i[119];
  assign o[61155] = i[119];
  assign o[61156] = i[119];
  assign o[61157] = i[119];
  assign o[61158] = i[119];
  assign o[61159] = i[119];
  assign o[61160] = i[119];
  assign o[61161] = i[119];
  assign o[61162] = i[119];
  assign o[61163] = i[119];
  assign o[61164] = i[119];
  assign o[61165] = i[119];
  assign o[61166] = i[119];
  assign o[61167] = i[119];
  assign o[61168] = i[119];
  assign o[61169] = i[119];
  assign o[61170] = i[119];
  assign o[61171] = i[119];
  assign o[61172] = i[119];
  assign o[61173] = i[119];
  assign o[61174] = i[119];
  assign o[61175] = i[119];
  assign o[61176] = i[119];
  assign o[61177] = i[119];
  assign o[61178] = i[119];
  assign o[61179] = i[119];
  assign o[61180] = i[119];
  assign o[61181] = i[119];
  assign o[61182] = i[119];
  assign o[61183] = i[119];
  assign o[61184] = i[119];
  assign o[61185] = i[119];
  assign o[61186] = i[119];
  assign o[61187] = i[119];
  assign o[61188] = i[119];
  assign o[61189] = i[119];
  assign o[61190] = i[119];
  assign o[61191] = i[119];
  assign o[61192] = i[119];
  assign o[61193] = i[119];
  assign o[61194] = i[119];
  assign o[61195] = i[119];
  assign o[61196] = i[119];
  assign o[61197] = i[119];
  assign o[61198] = i[119];
  assign o[61199] = i[119];
  assign o[61200] = i[119];
  assign o[61201] = i[119];
  assign o[61202] = i[119];
  assign o[61203] = i[119];
  assign o[61204] = i[119];
  assign o[61205] = i[119];
  assign o[61206] = i[119];
  assign o[61207] = i[119];
  assign o[61208] = i[119];
  assign o[61209] = i[119];
  assign o[61210] = i[119];
  assign o[61211] = i[119];
  assign o[61212] = i[119];
  assign o[61213] = i[119];
  assign o[61214] = i[119];
  assign o[61215] = i[119];
  assign o[61216] = i[119];
  assign o[61217] = i[119];
  assign o[61218] = i[119];
  assign o[61219] = i[119];
  assign o[61220] = i[119];
  assign o[61221] = i[119];
  assign o[61222] = i[119];
  assign o[61223] = i[119];
  assign o[61224] = i[119];
  assign o[61225] = i[119];
  assign o[61226] = i[119];
  assign o[61227] = i[119];
  assign o[61228] = i[119];
  assign o[61229] = i[119];
  assign o[61230] = i[119];
  assign o[61231] = i[119];
  assign o[61232] = i[119];
  assign o[61233] = i[119];
  assign o[61234] = i[119];
  assign o[61235] = i[119];
  assign o[61236] = i[119];
  assign o[61237] = i[119];
  assign o[61238] = i[119];
  assign o[61239] = i[119];
  assign o[61240] = i[119];
  assign o[61241] = i[119];
  assign o[61242] = i[119];
  assign o[61243] = i[119];
  assign o[61244] = i[119];
  assign o[61245] = i[119];
  assign o[61246] = i[119];
  assign o[61247] = i[119];
  assign o[61248] = i[119];
  assign o[61249] = i[119];
  assign o[61250] = i[119];
  assign o[61251] = i[119];
  assign o[61252] = i[119];
  assign o[61253] = i[119];
  assign o[61254] = i[119];
  assign o[61255] = i[119];
  assign o[61256] = i[119];
  assign o[61257] = i[119];
  assign o[61258] = i[119];
  assign o[61259] = i[119];
  assign o[61260] = i[119];
  assign o[61261] = i[119];
  assign o[61262] = i[119];
  assign o[61263] = i[119];
  assign o[61264] = i[119];
  assign o[61265] = i[119];
  assign o[61266] = i[119];
  assign o[61267] = i[119];
  assign o[61268] = i[119];
  assign o[61269] = i[119];
  assign o[61270] = i[119];
  assign o[61271] = i[119];
  assign o[61272] = i[119];
  assign o[61273] = i[119];
  assign o[61274] = i[119];
  assign o[61275] = i[119];
  assign o[61276] = i[119];
  assign o[61277] = i[119];
  assign o[61278] = i[119];
  assign o[61279] = i[119];
  assign o[61280] = i[119];
  assign o[61281] = i[119];
  assign o[61282] = i[119];
  assign o[61283] = i[119];
  assign o[61284] = i[119];
  assign o[61285] = i[119];
  assign o[61286] = i[119];
  assign o[61287] = i[119];
  assign o[61288] = i[119];
  assign o[61289] = i[119];
  assign o[61290] = i[119];
  assign o[61291] = i[119];
  assign o[61292] = i[119];
  assign o[61293] = i[119];
  assign o[61294] = i[119];
  assign o[61295] = i[119];
  assign o[61296] = i[119];
  assign o[61297] = i[119];
  assign o[61298] = i[119];
  assign o[61299] = i[119];
  assign o[61300] = i[119];
  assign o[61301] = i[119];
  assign o[61302] = i[119];
  assign o[61303] = i[119];
  assign o[61304] = i[119];
  assign o[61305] = i[119];
  assign o[61306] = i[119];
  assign o[61307] = i[119];
  assign o[61308] = i[119];
  assign o[61309] = i[119];
  assign o[61310] = i[119];
  assign o[61311] = i[119];
  assign o[61312] = i[119];
  assign o[61313] = i[119];
  assign o[61314] = i[119];
  assign o[61315] = i[119];
  assign o[61316] = i[119];
  assign o[61317] = i[119];
  assign o[61318] = i[119];
  assign o[61319] = i[119];
  assign o[61320] = i[119];
  assign o[61321] = i[119];
  assign o[61322] = i[119];
  assign o[61323] = i[119];
  assign o[61324] = i[119];
  assign o[61325] = i[119];
  assign o[61326] = i[119];
  assign o[61327] = i[119];
  assign o[61328] = i[119];
  assign o[61329] = i[119];
  assign o[61330] = i[119];
  assign o[61331] = i[119];
  assign o[61332] = i[119];
  assign o[61333] = i[119];
  assign o[61334] = i[119];
  assign o[61335] = i[119];
  assign o[61336] = i[119];
  assign o[61337] = i[119];
  assign o[61338] = i[119];
  assign o[61339] = i[119];
  assign o[61340] = i[119];
  assign o[61341] = i[119];
  assign o[61342] = i[119];
  assign o[61343] = i[119];
  assign o[61344] = i[119];
  assign o[61345] = i[119];
  assign o[61346] = i[119];
  assign o[61347] = i[119];
  assign o[61348] = i[119];
  assign o[61349] = i[119];
  assign o[61350] = i[119];
  assign o[61351] = i[119];
  assign o[61352] = i[119];
  assign o[61353] = i[119];
  assign o[61354] = i[119];
  assign o[61355] = i[119];
  assign o[61356] = i[119];
  assign o[61357] = i[119];
  assign o[61358] = i[119];
  assign o[61359] = i[119];
  assign o[61360] = i[119];
  assign o[61361] = i[119];
  assign o[61362] = i[119];
  assign o[61363] = i[119];
  assign o[61364] = i[119];
  assign o[61365] = i[119];
  assign o[61366] = i[119];
  assign o[61367] = i[119];
  assign o[61368] = i[119];
  assign o[61369] = i[119];
  assign o[61370] = i[119];
  assign o[61371] = i[119];
  assign o[61372] = i[119];
  assign o[61373] = i[119];
  assign o[61374] = i[119];
  assign o[61375] = i[119];
  assign o[61376] = i[119];
  assign o[61377] = i[119];
  assign o[61378] = i[119];
  assign o[61379] = i[119];
  assign o[61380] = i[119];
  assign o[61381] = i[119];
  assign o[61382] = i[119];
  assign o[61383] = i[119];
  assign o[61384] = i[119];
  assign o[61385] = i[119];
  assign o[61386] = i[119];
  assign o[61387] = i[119];
  assign o[61388] = i[119];
  assign o[61389] = i[119];
  assign o[61390] = i[119];
  assign o[61391] = i[119];
  assign o[61392] = i[119];
  assign o[61393] = i[119];
  assign o[61394] = i[119];
  assign o[61395] = i[119];
  assign o[61396] = i[119];
  assign o[61397] = i[119];
  assign o[61398] = i[119];
  assign o[61399] = i[119];
  assign o[61400] = i[119];
  assign o[61401] = i[119];
  assign o[61402] = i[119];
  assign o[61403] = i[119];
  assign o[61404] = i[119];
  assign o[61405] = i[119];
  assign o[61406] = i[119];
  assign o[61407] = i[119];
  assign o[61408] = i[119];
  assign o[61409] = i[119];
  assign o[61410] = i[119];
  assign o[61411] = i[119];
  assign o[61412] = i[119];
  assign o[61413] = i[119];
  assign o[61414] = i[119];
  assign o[61415] = i[119];
  assign o[61416] = i[119];
  assign o[61417] = i[119];
  assign o[61418] = i[119];
  assign o[61419] = i[119];
  assign o[61420] = i[119];
  assign o[61421] = i[119];
  assign o[61422] = i[119];
  assign o[61423] = i[119];
  assign o[61424] = i[119];
  assign o[61425] = i[119];
  assign o[61426] = i[119];
  assign o[61427] = i[119];
  assign o[61428] = i[119];
  assign o[61429] = i[119];
  assign o[61430] = i[119];
  assign o[61431] = i[119];
  assign o[61432] = i[119];
  assign o[61433] = i[119];
  assign o[61434] = i[119];
  assign o[61435] = i[119];
  assign o[61436] = i[119];
  assign o[61437] = i[119];
  assign o[61438] = i[119];
  assign o[61439] = i[119];
  assign o[60416] = i[118];
  assign o[60417] = i[118];
  assign o[60418] = i[118];
  assign o[60419] = i[118];
  assign o[60420] = i[118];
  assign o[60421] = i[118];
  assign o[60422] = i[118];
  assign o[60423] = i[118];
  assign o[60424] = i[118];
  assign o[60425] = i[118];
  assign o[60426] = i[118];
  assign o[60427] = i[118];
  assign o[60428] = i[118];
  assign o[60429] = i[118];
  assign o[60430] = i[118];
  assign o[60431] = i[118];
  assign o[60432] = i[118];
  assign o[60433] = i[118];
  assign o[60434] = i[118];
  assign o[60435] = i[118];
  assign o[60436] = i[118];
  assign o[60437] = i[118];
  assign o[60438] = i[118];
  assign o[60439] = i[118];
  assign o[60440] = i[118];
  assign o[60441] = i[118];
  assign o[60442] = i[118];
  assign o[60443] = i[118];
  assign o[60444] = i[118];
  assign o[60445] = i[118];
  assign o[60446] = i[118];
  assign o[60447] = i[118];
  assign o[60448] = i[118];
  assign o[60449] = i[118];
  assign o[60450] = i[118];
  assign o[60451] = i[118];
  assign o[60452] = i[118];
  assign o[60453] = i[118];
  assign o[60454] = i[118];
  assign o[60455] = i[118];
  assign o[60456] = i[118];
  assign o[60457] = i[118];
  assign o[60458] = i[118];
  assign o[60459] = i[118];
  assign o[60460] = i[118];
  assign o[60461] = i[118];
  assign o[60462] = i[118];
  assign o[60463] = i[118];
  assign o[60464] = i[118];
  assign o[60465] = i[118];
  assign o[60466] = i[118];
  assign o[60467] = i[118];
  assign o[60468] = i[118];
  assign o[60469] = i[118];
  assign o[60470] = i[118];
  assign o[60471] = i[118];
  assign o[60472] = i[118];
  assign o[60473] = i[118];
  assign o[60474] = i[118];
  assign o[60475] = i[118];
  assign o[60476] = i[118];
  assign o[60477] = i[118];
  assign o[60478] = i[118];
  assign o[60479] = i[118];
  assign o[60480] = i[118];
  assign o[60481] = i[118];
  assign o[60482] = i[118];
  assign o[60483] = i[118];
  assign o[60484] = i[118];
  assign o[60485] = i[118];
  assign o[60486] = i[118];
  assign o[60487] = i[118];
  assign o[60488] = i[118];
  assign o[60489] = i[118];
  assign o[60490] = i[118];
  assign o[60491] = i[118];
  assign o[60492] = i[118];
  assign o[60493] = i[118];
  assign o[60494] = i[118];
  assign o[60495] = i[118];
  assign o[60496] = i[118];
  assign o[60497] = i[118];
  assign o[60498] = i[118];
  assign o[60499] = i[118];
  assign o[60500] = i[118];
  assign o[60501] = i[118];
  assign o[60502] = i[118];
  assign o[60503] = i[118];
  assign o[60504] = i[118];
  assign o[60505] = i[118];
  assign o[60506] = i[118];
  assign o[60507] = i[118];
  assign o[60508] = i[118];
  assign o[60509] = i[118];
  assign o[60510] = i[118];
  assign o[60511] = i[118];
  assign o[60512] = i[118];
  assign o[60513] = i[118];
  assign o[60514] = i[118];
  assign o[60515] = i[118];
  assign o[60516] = i[118];
  assign o[60517] = i[118];
  assign o[60518] = i[118];
  assign o[60519] = i[118];
  assign o[60520] = i[118];
  assign o[60521] = i[118];
  assign o[60522] = i[118];
  assign o[60523] = i[118];
  assign o[60524] = i[118];
  assign o[60525] = i[118];
  assign o[60526] = i[118];
  assign o[60527] = i[118];
  assign o[60528] = i[118];
  assign o[60529] = i[118];
  assign o[60530] = i[118];
  assign o[60531] = i[118];
  assign o[60532] = i[118];
  assign o[60533] = i[118];
  assign o[60534] = i[118];
  assign o[60535] = i[118];
  assign o[60536] = i[118];
  assign o[60537] = i[118];
  assign o[60538] = i[118];
  assign o[60539] = i[118];
  assign o[60540] = i[118];
  assign o[60541] = i[118];
  assign o[60542] = i[118];
  assign o[60543] = i[118];
  assign o[60544] = i[118];
  assign o[60545] = i[118];
  assign o[60546] = i[118];
  assign o[60547] = i[118];
  assign o[60548] = i[118];
  assign o[60549] = i[118];
  assign o[60550] = i[118];
  assign o[60551] = i[118];
  assign o[60552] = i[118];
  assign o[60553] = i[118];
  assign o[60554] = i[118];
  assign o[60555] = i[118];
  assign o[60556] = i[118];
  assign o[60557] = i[118];
  assign o[60558] = i[118];
  assign o[60559] = i[118];
  assign o[60560] = i[118];
  assign o[60561] = i[118];
  assign o[60562] = i[118];
  assign o[60563] = i[118];
  assign o[60564] = i[118];
  assign o[60565] = i[118];
  assign o[60566] = i[118];
  assign o[60567] = i[118];
  assign o[60568] = i[118];
  assign o[60569] = i[118];
  assign o[60570] = i[118];
  assign o[60571] = i[118];
  assign o[60572] = i[118];
  assign o[60573] = i[118];
  assign o[60574] = i[118];
  assign o[60575] = i[118];
  assign o[60576] = i[118];
  assign o[60577] = i[118];
  assign o[60578] = i[118];
  assign o[60579] = i[118];
  assign o[60580] = i[118];
  assign o[60581] = i[118];
  assign o[60582] = i[118];
  assign o[60583] = i[118];
  assign o[60584] = i[118];
  assign o[60585] = i[118];
  assign o[60586] = i[118];
  assign o[60587] = i[118];
  assign o[60588] = i[118];
  assign o[60589] = i[118];
  assign o[60590] = i[118];
  assign o[60591] = i[118];
  assign o[60592] = i[118];
  assign o[60593] = i[118];
  assign o[60594] = i[118];
  assign o[60595] = i[118];
  assign o[60596] = i[118];
  assign o[60597] = i[118];
  assign o[60598] = i[118];
  assign o[60599] = i[118];
  assign o[60600] = i[118];
  assign o[60601] = i[118];
  assign o[60602] = i[118];
  assign o[60603] = i[118];
  assign o[60604] = i[118];
  assign o[60605] = i[118];
  assign o[60606] = i[118];
  assign o[60607] = i[118];
  assign o[60608] = i[118];
  assign o[60609] = i[118];
  assign o[60610] = i[118];
  assign o[60611] = i[118];
  assign o[60612] = i[118];
  assign o[60613] = i[118];
  assign o[60614] = i[118];
  assign o[60615] = i[118];
  assign o[60616] = i[118];
  assign o[60617] = i[118];
  assign o[60618] = i[118];
  assign o[60619] = i[118];
  assign o[60620] = i[118];
  assign o[60621] = i[118];
  assign o[60622] = i[118];
  assign o[60623] = i[118];
  assign o[60624] = i[118];
  assign o[60625] = i[118];
  assign o[60626] = i[118];
  assign o[60627] = i[118];
  assign o[60628] = i[118];
  assign o[60629] = i[118];
  assign o[60630] = i[118];
  assign o[60631] = i[118];
  assign o[60632] = i[118];
  assign o[60633] = i[118];
  assign o[60634] = i[118];
  assign o[60635] = i[118];
  assign o[60636] = i[118];
  assign o[60637] = i[118];
  assign o[60638] = i[118];
  assign o[60639] = i[118];
  assign o[60640] = i[118];
  assign o[60641] = i[118];
  assign o[60642] = i[118];
  assign o[60643] = i[118];
  assign o[60644] = i[118];
  assign o[60645] = i[118];
  assign o[60646] = i[118];
  assign o[60647] = i[118];
  assign o[60648] = i[118];
  assign o[60649] = i[118];
  assign o[60650] = i[118];
  assign o[60651] = i[118];
  assign o[60652] = i[118];
  assign o[60653] = i[118];
  assign o[60654] = i[118];
  assign o[60655] = i[118];
  assign o[60656] = i[118];
  assign o[60657] = i[118];
  assign o[60658] = i[118];
  assign o[60659] = i[118];
  assign o[60660] = i[118];
  assign o[60661] = i[118];
  assign o[60662] = i[118];
  assign o[60663] = i[118];
  assign o[60664] = i[118];
  assign o[60665] = i[118];
  assign o[60666] = i[118];
  assign o[60667] = i[118];
  assign o[60668] = i[118];
  assign o[60669] = i[118];
  assign o[60670] = i[118];
  assign o[60671] = i[118];
  assign o[60672] = i[118];
  assign o[60673] = i[118];
  assign o[60674] = i[118];
  assign o[60675] = i[118];
  assign o[60676] = i[118];
  assign o[60677] = i[118];
  assign o[60678] = i[118];
  assign o[60679] = i[118];
  assign o[60680] = i[118];
  assign o[60681] = i[118];
  assign o[60682] = i[118];
  assign o[60683] = i[118];
  assign o[60684] = i[118];
  assign o[60685] = i[118];
  assign o[60686] = i[118];
  assign o[60687] = i[118];
  assign o[60688] = i[118];
  assign o[60689] = i[118];
  assign o[60690] = i[118];
  assign o[60691] = i[118];
  assign o[60692] = i[118];
  assign o[60693] = i[118];
  assign o[60694] = i[118];
  assign o[60695] = i[118];
  assign o[60696] = i[118];
  assign o[60697] = i[118];
  assign o[60698] = i[118];
  assign o[60699] = i[118];
  assign o[60700] = i[118];
  assign o[60701] = i[118];
  assign o[60702] = i[118];
  assign o[60703] = i[118];
  assign o[60704] = i[118];
  assign o[60705] = i[118];
  assign o[60706] = i[118];
  assign o[60707] = i[118];
  assign o[60708] = i[118];
  assign o[60709] = i[118];
  assign o[60710] = i[118];
  assign o[60711] = i[118];
  assign o[60712] = i[118];
  assign o[60713] = i[118];
  assign o[60714] = i[118];
  assign o[60715] = i[118];
  assign o[60716] = i[118];
  assign o[60717] = i[118];
  assign o[60718] = i[118];
  assign o[60719] = i[118];
  assign o[60720] = i[118];
  assign o[60721] = i[118];
  assign o[60722] = i[118];
  assign o[60723] = i[118];
  assign o[60724] = i[118];
  assign o[60725] = i[118];
  assign o[60726] = i[118];
  assign o[60727] = i[118];
  assign o[60728] = i[118];
  assign o[60729] = i[118];
  assign o[60730] = i[118];
  assign o[60731] = i[118];
  assign o[60732] = i[118];
  assign o[60733] = i[118];
  assign o[60734] = i[118];
  assign o[60735] = i[118];
  assign o[60736] = i[118];
  assign o[60737] = i[118];
  assign o[60738] = i[118];
  assign o[60739] = i[118];
  assign o[60740] = i[118];
  assign o[60741] = i[118];
  assign o[60742] = i[118];
  assign o[60743] = i[118];
  assign o[60744] = i[118];
  assign o[60745] = i[118];
  assign o[60746] = i[118];
  assign o[60747] = i[118];
  assign o[60748] = i[118];
  assign o[60749] = i[118];
  assign o[60750] = i[118];
  assign o[60751] = i[118];
  assign o[60752] = i[118];
  assign o[60753] = i[118];
  assign o[60754] = i[118];
  assign o[60755] = i[118];
  assign o[60756] = i[118];
  assign o[60757] = i[118];
  assign o[60758] = i[118];
  assign o[60759] = i[118];
  assign o[60760] = i[118];
  assign o[60761] = i[118];
  assign o[60762] = i[118];
  assign o[60763] = i[118];
  assign o[60764] = i[118];
  assign o[60765] = i[118];
  assign o[60766] = i[118];
  assign o[60767] = i[118];
  assign o[60768] = i[118];
  assign o[60769] = i[118];
  assign o[60770] = i[118];
  assign o[60771] = i[118];
  assign o[60772] = i[118];
  assign o[60773] = i[118];
  assign o[60774] = i[118];
  assign o[60775] = i[118];
  assign o[60776] = i[118];
  assign o[60777] = i[118];
  assign o[60778] = i[118];
  assign o[60779] = i[118];
  assign o[60780] = i[118];
  assign o[60781] = i[118];
  assign o[60782] = i[118];
  assign o[60783] = i[118];
  assign o[60784] = i[118];
  assign o[60785] = i[118];
  assign o[60786] = i[118];
  assign o[60787] = i[118];
  assign o[60788] = i[118];
  assign o[60789] = i[118];
  assign o[60790] = i[118];
  assign o[60791] = i[118];
  assign o[60792] = i[118];
  assign o[60793] = i[118];
  assign o[60794] = i[118];
  assign o[60795] = i[118];
  assign o[60796] = i[118];
  assign o[60797] = i[118];
  assign o[60798] = i[118];
  assign o[60799] = i[118];
  assign o[60800] = i[118];
  assign o[60801] = i[118];
  assign o[60802] = i[118];
  assign o[60803] = i[118];
  assign o[60804] = i[118];
  assign o[60805] = i[118];
  assign o[60806] = i[118];
  assign o[60807] = i[118];
  assign o[60808] = i[118];
  assign o[60809] = i[118];
  assign o[60810] = i[118];
  assign o[60811] = i[118];
  assign o[60812] = i[118];
  assign o[60813] = i[118];
  assign o[60814] = i[118];
  assign o[60815] = i[118];
  assign o[60816] = i[118];
  assign o[60817] = i[118];
  assign o[60818] = i[118];
  assign o[60819] = i[118];
  assign o[60820] = i[118];
  assign o[60821] = i[118];
  assign o[60822] = i[118];
  assign o[60823] = i[118];
  assign o[60824] = i[118];
  assign o[60825] = i[118];
  assign o[60826] = i[118];
  assign o[60827] = i[118];
  assign o[60828] = i[118];
  assign o[60829] = i[118];
  assign o[60830] = i[118];
  assign o[60831] = i[118];
  assign o[60832] = i[118];
  assign o[60833] = i[118];
  assign o[60834] = i[118];
  assign o[60835] = i[118];
  assign o[60836] = i[118];
  assign o[60837] = i[118];
  assign o[60838] = i[118];
  assign o[60839] = i[118];
  assign o[60840] = i[118];
  assign o[60841] = i[118];
  assign o[60842] = i[118];
  assign o[60843] = i[118];
  assign o[60844] = i[118];
  assign o[60845] = i[118];
  assign o[60846] = i[118];
  assign o[60847] = i[118];
  assign o[60848] = i[118];
  assign o[60849] = i[118];
  assign o[60850] = i[118];
  assign o[60851] = i[118];
  assign o[60852] = i[118];
  assign o[60853] = i[118];
  assign o[60854] = i[118];
  assign o[60855] = i[118];
  assign o[60856] = i[118];
  assign o[60857] = i[118];
  assign o[60858] = i[118];
  assign o[60859] = i[118];
  assign o[60860] = i[118];
  assign o[60861] = i[118];
  assign o[60862] = i[118];
  assign o[60863] = i[118];
  assign o[60864] = i[118];
  assign o[60865] = i[118];
  assign o[60866] = i[118];
  assign o[60867] = i[118];
  assign o[60868] = i[118];
  assign o[60869] = i[118];
  assign o[60870] = i[118];
  assign o[60871] = i[118];
  assign o[60872] = i[118];
  assign o[60873] = i[118];
  assign o[60874] = i[118];
  assign o[60875] = i[118];
  assign o[60876] = i[118];
  assign o[60877] = i[118];
  assign o[60878] = i[118];
  assign o[60879] = i[118];
  assign o[60880] = i[118];
  assign o[60881] = i[118];
  assign o[60882] = i[118];
  assign o[60883] = i[118];
  assign o[60884] = i[118];
  assign o[60885] = i[118];
  assign o[60886] = i[118];
  assign o[60887] = i[118];
  assign o[60888] = i[118];
  assign o[60889] = i[118];
  assign o[60890] = i[118];
  assign o[60891] = i[118];
  assign o[60892] = i[118];
  assign o[60893] = i[118];
  assign o[60894] = i[118];
  assign o[60895] = i[118];
  assign o[60896] = i[118];
  assign o[60897] = i[118];
  assign o[60898] = i[118];
  assign o[60899] = i[118];
  assign o[60900] = i[118];
  assign o[60901] = i[118];
  assign o[60902] = i[118];
  assign o[60903] = i[118];
  assign o[60904] = i[118];
  assign o[60905] = i[118];
  assign o[60906] = i[118];
  assign o[60907] = i[118];
  assign o[60908] = i[118];
  assign o[60909] = i[118];
  assign o[60910] = i[118];
  assign o[60911] = i[118];
  assign o[60912] = i[118];
  assign o[60913] = i[118];
  assign o[60914] = i[118];
  assign o[60915] = i[118];
  assign o[60916] = i[118];
  assign o[60917] = i[118];
  assign o[60918] = i[118];
  assign o[60919] = i[118];
  assign o[60920] = i[118];
  assign o[60921] = i[118];
  assign o[60922] = i[118];
  assign o[60923] = i[118];
  assign o[60924] = i[118];
  assign o[60925] = i[118];
  assign o[60926] = i[118];
  assign o[60927] = i[118];
  assign o[59904] = i[117];
  assign o[59905] = i[117];
  assign o[59906] = i[117];
  assign o[59907] = i[117];
  assign o[59908] = i[117];
  assign o[59909] = i[117];
  assign o[59910] = i[117];
  assign o[59911] = i[117];
  assign o[59912] = i[117];
  assign o[59913] = i[117];
  assign o[59914] = i[117];
  assign o[59915] = i[117];
  assign o[59916] = i[117];
  assign o[59917] = i[117];
  assign o[59918] = i[117];
  assign o[59919] = i[117];
  assign o[59920] = i[117];
  assign o[59921] = i[117];
  assign o[59922] = i[117];
  assign o[59923] = i[117];
  assign o[59924] = i[117];
  assign o[59925] = i[117];
  assign o[59926] = i[117];
  assign o[59927] = i[117];
  assign o[59928] = i[117];
  assign o[59929] = i[117];
  assign o[59930] = i[117];
  assign o[59931] = i[117];
  assign o[59932] = i[117];
  assign o[59933] = i[117];
  assign o[59934] = i[117];
  assign o[59935] = i[117];
  assign o[59936] = i[117];
  assign o[59937] = i[117];
  assign o[59938] = i[117];
  assign o[59939] = i[117];
  assign o[59940] = i[117];
  assign o[59941] = i[117];
  assign o[59942] = i[117];
  assign o[59943] = i[117];
  assign o[59944] = i[117];
  assign o[59945] = i[117];
  assign o[59946] = i[117];
  assign o[59947] = i[117];
  assign o[59948] = i[117];
  assign o[59949] = i[117];
  assign o[59950] = i[117];
  assign o[59951] = i[117];
  assign o[59952] = i[117];
  assign o[59953] = i[117];
  assign o[59954] = i[117];
  assign o[59955] = i[117];
  assign o[59956] = i[117];
  assign o[59957] = i[117];
  assign o[59958] = i[117];
  assign o[59959] = i[117];
  assign o[59960] = i[117];
  assign o[59961] = i[117];
  assign o[59962] = i[117];
  assign o[59963] = i[117];
  assign o[59964] = i[117];
  assign o[59965] = i[117];
  assign o[59966] = i[117];
  assign o[59967] = i[117];
  assign o[59968] = i[117];
  assign o[59969] = i[117];
  assign o[59970] = i[117];
  assign o[59971] = i[117];
  assign o[59972] = i[117];
  assign o[59973] = i[117];
  assign o[59974] = i[117];
  assign o[59975] = i[117];
  assign o[59976] = i[117];
  assign o[59977] = i[117];
  assign o[59978] = i[117];
  assign o[59979] = i[117];
  assign o[59980] = i[117];
  assign o[59981] = i[117];
  assign o[59982] = i[117];
  assign o[59983] = i[117];
  assign o[59984] = i[117];
  assign o[59985] = i[117];
  assign o[59986] = i[117];
  assign o[59987] = i[117];
  assign o[59988] = i[117];
  assign o[59989] = i[117];
  assign o[59990] = i[117];
  assign o[59991] = i[117];
  assign o[59992] = i[117];
  assign o[59993] = i[117];
  assign o[59994] = i[117];
  assign o[59995] = i[117];
  assign o[59996] = i[117];
  assign o[59997] = i[117];
  assign o[59998] = i[117];
  assign o[59999] = i[117];
  assign o[60000] = i[117];
  assign o[60001] = i[117];
  assign o[60002] = i[117];
  assign o[60003] = i[117];
  assign o[60004] = i[117];
  assign o[60005] = i[117];
  assign o[60006] = i[117];
  assign o[60007] = i[117];
  assign o[60008] = i[117];
  assign o[60009] = i[117];
  assign o[60010] = i[117];
  assign o[60011] = i[117];
  assign o[60012] = i[117];
  assign o[60013] = i[117];
  assign o[60014] = i[117];
  assign o[60015] = i[117];
  assign o[60016] = i[117];
  assign o[60017] = i[117];
  assign o[60018] = i[117];
  assign o[60019] = i[117];
  assign o[60020] = i[117];
  assign o[60021] = i[117];
  assign o[60022] = i[117];
  assign o[60023] = i[117];
  assign o[60024] = i[117];
  assign o[60025] = i[117];
  assign o[60026] = i[117];
  assign o[60027] = i[117];
  assign o[60028] = i[117];
  assign o[60029] = i[117];
  assign o[60030] = i[117];
  assign o[60031] = i[117];
  assign o[60032] = i[117];
  assign o[60033] = i[117];
  assign o[60034] = i[117];
  assign o[60035] = i[117];
  assign o[60036] = i[117];
  assign o[60037] = i[117];
  assign o[60038] = i[117];
  assign o[60039] = i[117];
  assign o[60040] = i[117];
  assign o[60041] = i[117];
  assign o[60042] = i[117];
  assign o[60043] = i[117];
  assign o[60044] = i[117];
  assign o[60045] = i[117];
  assign o[60046] = i[117];
  assign o[60047] = i[117];
  assign o[60048] = i[117];
  assign o[60049] = i[117];
  assign o[60050] = i[117];
  assign o[60051] = i[117];
  assign o[60052] = i[117];
  assign o[60053] = i[117];
  assign o[60054] = i[117];
  assign o[60055] = i[117];
  assign o[60056] = i[117];
  assign o[60057] = i[117];
  assign o[60058] = i[117];
  assign o[60059] = i[117];
  assign o[60060] = i[117];
  assign o[60061] = i[117];
  assign o[60062] = i[117];
  assign o[60063] = i[117];
  assign o[60064] = i[117];
  assign o[60065] = i[117];
  assign o[60066] = i[117];
  assign o[60067] = i[117];
  assign o[60068] = i[117];
  assign o[60069] = i[117];
  assign o[60070] = i[117];
  assign o[60071] = i[117];
  assign o[60072] = i[117];
  assign o[60073] = i[117];
  assign o[60074] = i[117];
  assign o[60075] = i[117];
  assign o[60076] = i[117];
  assign o[60077] = i[117];
  assign o[60078] = i[117];
  assign o[60079] = i[117];
  assign o[60080] = i[117];
  assign o[60081] = i[117];
  assign o[60082] = i[117];
  assign o[60083] = i[117];
  assign o[60084] = i[117];
  assign o[60085] = i[117];
  assign o[60086] = i[117];
  assign o[60087] = i[117];
  assign o[60088] = i[117];
  assign o[60089] = i[117];
  assign o[60090] = i[117];
  assign o[60091] = i[117];
  assign o[60092] = i[117];
  assign o[60093] = i[117];
  assign o[60094] = i[117];
  assign o[60095] = i[117];
  assign o[60096] = i[117];
  assign o[60097] = i[117];
  assign o[60098] = i[117];
  assign o[60099] = i[117];
  assign o[60100] = i[117];
  assign o[60101] = i[117];
  assign o[60102] = i[117];
  assign o[60103] = i[117];
  assign o[60104] = i[117];
  assign o[60105] = i[117];
  assign o[60106] = i[117];
  assign o[60107] = i[117];
  assign o[60108] = i[117];
  assign o[60109] = i[117];
  assign o[60110] = i[117];
  assign o[60111] = i[117];
  assign o[60112] = i[117];
  assign o[60113] = i[117];
  assign o[60114] = i[117];
  assign o[60115] = i[117];
  assign o[60116] = i[117];
  assign o[60117] = i[117];
  assign o[60118] = i[117];
  assign o[60119] = i[117];
  assign o[60120] = i[117];
  assign o[60121] = i[117];
  assign o[60122] = i[117];
  assign o[60123] = i[117];
  assign o[60124] = i[117];
  assign o[60125] = i[117];
  assign o[60126] = i[117];
  assign o[60127] = i[117];
  assign o[60128] = i[117];
  assign o[60129] = i[117];
  assign o[60130] = i[117];
  assign o[60131] = i[117];
  assign o[60132] = i[117];
  assign o[60133] = i[117];
  assign o[60134] = i[117];
  assign o[60135] = i[117];
  assign o[60136] = i[117];
  assign o[60137] = i[117];
  assign o[60138] = i[117];
  assign o[60139] = i[117];
  assign o[60140] = i[117];
  assign o[60141] = i[117];
  assign o[60142] = i[117];
  assign o[60143] = i[117];
  assign o[60144] = i[117];
  assign o[60145] = i[117];
  assign o[60146] = i[117];
  assign o[60147] = i[117];
  assign o[60148] = i[117];
  assign o[60149] = i[117];
  assign o[60150] = i[117];
  assign o[60151] = i[117];
  assign o[60152] = i[117];
  assign o[60153] = i[117];
  assign o[60154] = i[117];
  assign o[60155] = i[117];
  assign o[60156] = i[117];
  assign o[60157] = i[117];
  assign o[60158] = i[117];
  assign o[60159] = i[117];
  assign o[60160] = i[117];
  assign o[60161] = i[117];
  assign o[60162] = i[117];
  assign o[60163] = i[117];
  assign o[60164] = i[117];
  assign o[60165] = i[117];
  assign o[60166] = i[117];
  assign o[60167] = i[117];
  assign o[60168] = i[117];
  assign o[60169] = i[117];
  assign o[60170] = i[117];
  assign o[60171] = i[117];
  assign o[60172] = i[117];
  assign o[60173] = i[117];
  assign o[60174] = i[117];
  assign o[60175] = i[117];
  assign o[60176] = i[117];
  assign o[60177] = i[117];
  assign o[60178] = i[117];
  assign o[60179] = i[117];
  assign o[60180] = i[117];
  assign o[60181] = i[117];
  assign o[60182] = i[117];
  assign o[60183] = i[117];
  assign o[60184] = i[117];
  assign o[60185] = i[117];
  assign o[60186] = i[117];
  assign o[60187] = i[117];
  assign o[60188] = i[117];
  assign o[60189] = i[117];
  assign o[60190] = i[117];
  assign o[60191] = i[117];
  assign o[60192] = i[117];
  assign o[60193] = i[117];
  assign o[60194] = i[117];
  assign o[60195] = i[117];
  assign o[60196] = i[117];
  assign o[60197] = i[117];
  assign o[60198] = i[117];
  assign o[60199] = i[117];
  assign o[60200] = i[117];
  assign o[60201] = i[117];
  assign o[60202] = i[117];
  assign o[60203] = i[117];
  assign o[60204] = i[117];
  assign o[60205] = i[117];
  assign o[60206] = i[117];
  assign o[60207] = i[117];
  assign o[60208] = i[117];
  assign o[60209] = i[117];
  assign o[60210] = i[117];
  assign o[60211] = i[117];
  assign o[60212] = i[117];
  assign o[60213] = i[117];
  assign o[60214] = i[117];
  assign o[60215] = i[117];
  assign o[60216] = i[117];
  assign o[60217] = i[117];
  assign o[60218] = i[117];
  assign o[60219] = i[117];
  assign o[60220] = i[117];
  assign o[60221] = i[117];
  assign o[60222] = i[117];
  assign o[60223] = i[117];
  assign o[60224] = i[117];
  assign o[60225] = i[117];
  assign o[60226] = i[117];
  assign o[60227] = i[117];
  assign o[60228] = i[117];
  assign o[60229] = i[117];
  assign o[60230] = i[117];
  assign o[60231] = i[117];
  assign o[60232] = i[117];
  assign o[60233] = i[117];
  assign o[60234] = i[117];
  assign o[60235] = i[117];
  assign o[60236] = i[117];
  assign o[60237] = i[117];
  assign o[60238] = i[117];
  assign o[60239] = i[117];
  assign o[60240] = i[117];
  assign o[60241] = i[117];
  assign o[60242] = i[117];
  assign o[60243] = i[117];
  assign o[60244] = i[117];
  assign o[60245] = i[117];
  assign o[60246] = i[117];
  assign o[60247] = i[117];
  assign o[60248] = i[117];
  assign o[60249] = i[117];
  assign o[60250] = i[117];
  assign o[60251] = i[117];
  assign o[60252] = i[117];
  assign o[60253] = i[117];
  assign o[60254] = i[117];
  assign o[60255] = i[117];
  assign o[60256] = i[117];
  assign o[60257] = i[117];
  assign o[60258] = i[117];
  assign o[60259] = i[117];
  assign o[60260] = i[117];
  assign o[60261] = i[117];
  assign o[60262] = i[117];
  assign o[60263] = i[117];
  assign o[60264] = i[117];
  assign o[60265] = i[117];
  assign o[60266] = i[117];
  assign o[60267] = i[117];
  assign o[60268] = i[117];
  assign o[60269] = i[117];
  assign o[60270] = i[117];
  assign o[60271] = i[117];
  assign o[60272] = i[117];
  assign o[60273] = i[117];
  assign o[60274] = i[117];
  assign o[60275] = i[117];
  assign o[60276] = i[117];
  assign o[60277] = i[117];
  assign o[60278] = i[117];
  assign o[60279] = i[117];
  assign o[60280] = i[117];
  assign o[60281] = i[117];
  assign o[60282] = i[117];
  assign o[60283] = i[117];
  assign o[60284] = i[117];
  assign o[60285] = i[117];
  assign o[60286] = i[117];
  assign o[60287] = i[117];
  assign o[60288] = i[117];
  assign o[60289] = i[117];
  assign o[60290] = i[117];
  assign o[60291] = i[117];
  assign o[60292] = i[117];
  assign o[60293] = i[117];
  assign o[60294] = i[117];
  assign o[60295] = i[117];
  assign o[60296] = i[117];
  assign o[60297] = i[117];
  assign o[60298] = i[117];
  assign o[60299] = i[117];
  assign o[60300] = i[117];
  assign o[60301] = i[117];
  assign o[60302] = i[117];
  assign o[60303] = i[117];
  assign o[60304] = i[117];
  assign o[60305] = i[117];
  assign o[60306] = i[117];
  assign o[60307] = i[117];
  assign o[60308] = i[117];
  assign o[60309] = i[117];
  assign o[60310] = i[117];
  assign o[60311] = i[117];
  assign o[60312] = i[117];
  assign o[60313] = i[117];
  assign o[60314] = i[117];
  assign o[60315] = i[117];
  assign o[60316] = i[117];
  assign o[60317] = i[117];
  assign o[60318] = i[117];
  assign o[60319] = i[117];
  assign o[60320] = i[117];
  assign o[60321] = i[117];
  assign o[60322] = i[117];
  assign o[60323] = i[117];
  assign o[60324] = i[117];
  assign o[60325] = i[117];
  assign o[60326] = i[117];
  assign o[60327] = i[117];
  assign o[60328] = i[117];
  assign o[60329] = i[117];
  assign o[60330] = i[117];
  assign o[60331] = i[117];
  assign o[60332] = i[117];
  assign o[60333] = i[117];
  assign o[60334] = i[117];
  assign o[60335] = i[117];
  assign o[60336] = i[117];
  assign o[60337] = i[117];
  assign o[60338] = i[117];
  assign o[60339] = i[117];
  assign o[60340] = i[117];
  assign o[60341] = i[117];
  assign o[60342] = i[117];
  assign o[60343] = i[117];
  assign o[60344] = i[117];
  assign o[60345] = i[117];
  assign o[60346] = i[117];
  assign o[60347] = i[117];
  assign o[60348] = i[117];
  assign o[60349] = i[117];
  assign o[60350] = i[117];
  assign o[60351] = i[117];
  assign o[60352] = i[117];
  assign o[60353] = i[117];
  assign o[60354] = i[117];
  assign o[60355] = i[117];
  assign o[60356] = i[117];
  assign o[60357] = i[117];
  assign o[60358] = i[117];
  assign o[60359] = i[117];
  assign o[60360] = i[117];
  assign o[60361] = i[117];
  assign o[60362] = i[117];
  assign o[60363] = i[117];
  assign o[60364] = i[117];
  assign o[60365] = i[117];
  assign o[60366] = i[117];
  assign o[60367] = i[117];
  assign o[60368] = i[117];
  assign o[60369] = i[117];
  assign o[60370] = i[117];
  assign o[60371] = i[117];
  assign o[60372] = i[117];
  assign o[60373] = i[117];
  assign o[60374] = i[117];
  assign o[60375] = i[117];
  assign o[60376] = i[117];
  assign o[60377] = i[117];
  assign o[60378] = i[117];
  assign o[60379] = i[117];
  assign o[60380] = i[117];
  assign o[60381] = i[117];
  assign o[60382] = i[117];
  assign o[60383] = i[117];
  assign o[60384] = i[117];
  assign o[60385] = i[117];
  assign o[60386] = i[117];
  assign o[60387] = i[117];
  assign o[60388] = i[117];
  assign o[60389] = i[117];
  assign o[60390] = i[117];
  assign o[60391] = i[117];
  assign o[60392] = i[117];
  assign o[60393] = i[117];
  assign o[60394] = i[117];
  assign o[60395] = i[117];
  assign o[60396] = i[117];
  assign o[60397] = i[117];
  assign o[60398] = i[117];
  assign o[60399] = i[117];
  assign o[60400] = i[117];
  assign o[60401] = i[117];
  assign o[60402] = i[117];
  assign o[60403] = i[117];
  assign o[60404] = i[117];
  assign o[60405] = i[117];
  assign o[60406] = i[117];
  assign o[60407] = i[117];
  assign o[60408] = i[117];
  assign o[60409] = i[117];
  assign o[60410] = i[117];
  assign o[60411] = i[117];
  assign o[60412] = i[117];
  assign o[60413] = i[117];
  assign o[60414] = i[117];
  assign o[60415] = i[117];
  assign o[59392] = i[116];
  assign o[59393] = i[116];
  assign o[59394] = i[116];
  assign o[59395] = i[116];
  assign o[59396] = i[116];
  assign o[59397] = i[116];
  assign o[59398] = i[116];
  assign o[59399] = i[116];
  assign o[59400] = i[116];
  assign o[59401] = i[116];
  assign o[59402] = i[116];
  assign o[59403] = i[116];
  assign o[59404] = i[116];
  assign o[59405] = i[116];
  assign o[59406] = i[116];
  assign o[59407] = i[116];
  assign o[59408] = i[116];
  assign o[59409] = i[116];
  assign o[59410] = i[116];
  assign o[59411] = i[116];
  assign o[59412] = i[116];
  assign o[59413] = i[116];
  assign o[59414] = i[116];
  assign o[59415] = i[116];
  assign o[59416] = i[116];
  assign o[59417] = i[116];
  assign o[59418] = i[116];
  assign o[59419] = i[116];
  assign o[59420] = i[116];
  assign o[59421] = i[116];
  assign o[59422] = i[116];
  assign o[59423] = i[116];
  assign o[59424] = i[116];
  assign o[59425] = i[116];
  assign o[59426] = i[116];
  assign o[59427] = i[116];
  assign o[59428] = i[116];
  assign o[59429] = i[116];
  assign o[59430] = i[116];
  assign o[59431] = i[116];
  assign o[59432] = i[116];
  assign o[59433] = i[116];
  assign o[59434] = i[116];
  assign o[59435] = i[116];
  assign o[59436] = i[116];
  assign o[59437] = i[116];
  assign o[59438] = i[116];
  assign o[59439] = i[116];
  assign o[59440] = i[116];
  assign o[59441] = i[116];
  assign o[59442] = i[116];
  assign o[59443] = i[116];
  assign o[59444] = i[116];
  assign o[59445] = i[116];
  assign o[59446] = i[116];
  assign o[59447] = i[116];
  assign o[59448] = i[116];
  assign o[59449] = i[116];
  assign o[59450] = i[116];
  assign o[59451] = i[116];
  assign o[59452] = i[116];
  assign o[59453] = i[116];
  assign o[59454] = i[116];
  assign o[59455] = i[116];
  assign o[59456] = i[116];
  assign o[59457] = i[116];
  assign o[59458] = i[116];
  assign o[59459] = i[116];
  assign o[59460] = i[116];
  assign o[59461] = i[116];
  assign o[59462] = i[116];
  assign o[59463] = i[116];
  assign o[59464] = i[116];
  assign o[59465] = i[116];
  assign o[59466] = i[116];
  assign o[59467] = i[116];
  assign o[59468] = i[116];
  assign o[59469] = i[116];
  assign o[59470] = i[116];
  assign o[59471] = i[116];
  assign o[59472] = i[116];
  assign o[59473] = i[116];
  assign o[59474] = i[116];
  assign o[59475] = i[116];
  assign o[59476] = i[116];
  assign o[59477] = i[116];
  assign o[59478] = i[116];
  assign o[59479] = i[116];
  assign o[59480] = i[116];
  assign o[59481] = i[116];
  assign o[59482] = i[116];
  assign o[59483] = i[116];
  assign o[59484] = i[116];
  assign o[59485] = i[116];
  assign o[59486] = i[116];
  assign o[59487] = i[116];
  assign o[59488] = i[116];
  assign o[59489] = i[116];
  assign o[59490] = i[116];
  assign o[59491] = i[116];
  assign o[59492] = i[116];
  assign o[59493] = i[116];
  assign o[59494] = i[116];
  assign o[59495] = i[116];
  assign o[59496] = i[116];
  assign o[59497] = i[116];
  assign o[59498] = i[116];
  assign o[59499] = i[116];
  assign o[59500] = i[116];
  assign o[59501] = i[116];
  assign o[59502] = i[116];
  assign o[59503] = i[116];
  assign o[59504] = i[116];
  assign o[59505] = i[116];
  assign o[59506] = i[116];
  assign o[59507] = i[116];
  assign o[59508] = i[116];
  assign o[59509] = i[116];
  assign o[59510] = i[116];
  assign o[59511] = i[116];
  assign o[59512] = i[116];
  assign o[59513] = i[116];
  assign o[59514] = i[116];
  assign o[59515] = i[116];
  assign o[59516] = i[116];
  assign o[59517] = i[116];
  assign o[59518] = i[116];
  assign o[59519] = i[116];
  assign o[59520] = i[116];
  assign o[59521] = i[116];
  assign o[59522] = i[116];
  assign o[59523] = i[116];
  assign o[59524] = i[116];
  assign o[59525] = i[116];
  assign o[59526] = i[116];
  assign o[59527] = i[116];
  assign o[59528] = i[116];
  assign o[59529] = i[116];
  assign o[59530] = i[116];
  assign o[59531] = i[116];
  assign o[59532] = i[116];
  assign o[59533] = i[116];
  assign o[59534] = i[116];
  assign o[59535] = i[116];
  assign o[59536] = i[116];
  assign o[59537] = i[116];
  assign o[59538] = i[116];
  assign o[59539] = i[116];
  assign o[59540] = i[116];
  assign o[59541] = i[116];
  assign o[59542] = i[116];
  assign o[59543] = i[116];
  assign o[59544] = i[116];
  assign o[59545] = i[116];
  assign o[59546] = i[116];
  assign o[59547] = i[116];
  assign o[59548] = i[116];
  assign o[59549] = i[116];
  assign o[59550] = i[116];
  assign o[59551] = i[116];
  assign o[59552] = i[116];
  assign o[59553] = i[116];
  assign o[59554] = i[116];
  assign o[59555] = i[116];
  assign o[59556] = i[116];
  assign o[59557] = i[116];
  assign o[59558] = i[116];
  assign o[59559] = i[116];
  assign o[59560] = i[116];
  assign o[59561] = i[116];
  assign o[59562] = i[116];
  assign o[59563] = i[116];
  assign o[59564] = i[116];
  assign o[59565] = i[116];
  assign o[59566] = i[116];
  assign o[59567] = i[116];
  assign o[59568] = i[116];
  assign o[59569] = i[116];
  assign o[59570] = i[116];
  assign o[59571] = i[116];
  assign o[59572] = i[116];
  assign o[59573] = i[116];
  assign o[59574] = i[116];
  assign o[59575] = i[116];
  assign o[59576] = i[116];
  assign o[59577] = i[116];
  assign o[59578] = i[116];
  assign o[59579] = i[116];
  assign o[59580] = i[116];
  assign o[59581] = i[116];
  assign o[59582] = i[116];
  assign o[59583] = i[116];
  assign o[59584] = i[116];
  assign o[59585] = i[116];
  assign o[59586] = i[116];
  assign o[59587] = i[116];
  assign o[59588] = i[116];
  assign o[59589] = i[116];
  assign o[59590] = i[116];
  assign o[59591] = i[116];
  assign o[59592] = i[116];
  assign o[59593] = i[116];
  assign o[59594] = i[116];
  assign o[59595] = i[116];
  assign o[59596] = i[116];
  assign o[59597] = i[116];
  assign o[59598] = i[116];
  assign o[59599] = i[116];
  assign o[59600] = i[116];
  assign o[59601] = i[116];
  assign o[59602] = i[116];
  assign o[59603] = i[116];
  assign o[59604] = i[116];
  assign o[59605] = i[116];
  assign o[59606] = i[116];
  assign o[59607] = i[116];
  assign o[59608] = i[116];
  assign o[59609] = i[116];
  assign o[59610] = i[116];
  assign o[59611] = i[116];
  assign o[59612] = i[116];
  assign o[59613] = i[116];
  assign o[59614] = i[116];
  assign o[59615] = i[116];
  assign o[59616] = i[116];
  assign o[59617] = i[116];
  assign o[59618] = i[116];
  assign o[59619] = i[116];
  assign o[59620] = i[116];
  assign o[59621] = i[116];
  assign o[59622] = i[116];
  assign o[59623] = i[116];
  assign o[59624] = i[116];
  assign o[59625] = i[116];
  assign o[59626] = i[116];
  assign o[59627] = i[116];
  assign o[59628] = i[116];
  assign o[59629] = i[116];
  assign o[59630] = i[116];
  assign o[59631] = i[116];
  assign o[59632] = i[116];
  assign o[59633] = i[116];
  assign o[59634] = i[116];
  assign o[59635] = i[116];
  assign o[59636] = i[116];
  assign o[59637] = i[116];
  assign o[59638] = i[116];
  assign o[59639] = i[116];
  assign o[59640] = i[116];
  assign o[59641] = i[116];
  assign o[59642] = i[116];
  assign o[59643] = i[116];
  assign o[59644] = i[116];
  assign o[59645] = i[116];
  assign o[59646] = i[116];
  assign o[59647] = i[116];
  assign o[59648] = i[116];
  assign o[59649] = i[116];
  assign o[59650] = i[116];
  assign o[59651] = i[116];
  assign o[59652] = i[116];
  assign o[59653] = i[116];
  assign o[59654] = i[116];
  assign o[59655] = i[116];
  assign o[59656] = i[116];
  assign o[59657] = i[116];
  assign o[59658] = i[116];
  assign o[59659] = i[116];
  assign o[59660] = i[116];
  assign o[59661] = i[116];
  assign o[59662] = i[116];
  assign o[59663] = i[116];
  assign o[59664] = i[116];
  assign o[59665] = i[116];
  assign o[59666] = i[116];
  assign o[59667] = i[116];
  assign o[59668] = i[116];
  assign o[59669] = i[116];
  assign o[59670] = i[116];
  assign o[59671] = i[116];
  assign o[59672] = i[116];
  assign o[59673] = i[116];
  assign o[59674] = i[116];
  assign o[59675] = i[116];
  assign o[59676] = i[116];
  assign o[59677] = i[116];
  assign o[59678] = i[116];
  assign o[59679] = i[116];
  assign o[59680] = i[116];
  assign o[59681] = i[116];
  assign o[59682] = i[116];
  assign o[59683] = i[116];
  assign o[59684] = i[116];
  assign o[59685] = i[116];
  assign o[59686] = i[116];
  assign o[59687] = i[116];
  assign o[59688] = i[116];
  assign o[59689] = i[116];
  assign o[59690] = i[116];
  assign o[59691] = i[116];
  assign o[59692] = i[116];
  assign o[59693] = i[116];
  assign o[59694] = i[116];
  assign o[59695] = i[116];
  assign o[59696] = i[116];
  assign o[59697] = i[116];
  assign o[59698] = i[116];
  assign o[59699] = i[116];
  assign o[59700] = i[116];
  assign o[59701] = i[116];
  assign o[59702] = i[116];
  assign o[59703] = i[116];
  assign o[59704] = i[116];
  assign o[59705] = i[116];
  assign o[59706] = i[116];
  assign o[59707] = i[116];
  assign o[59708] = i[116];
  assign o[59709] = i[116];
  assign o[59710] = i[116];
  assign o[59711] = i[116];
  assign o[59712] = i[116];
  assign o[59713] = i[116];
  assign o[59714] = i[116];
  assign o[59715] = i[116];
  assign o[59716] = i[116];
  assign o[59717] = i[116];
  assign o[59718] = i[116];
  assign o[59719] = i[116];
  assign o[59720] = i[116];
  assign o[59721] = i[116];
  assign o[59722] = i[116];
  assign o[59723] = i[116];
  assign o[59724] = i[116];
  assign o[59725] = i[116];
  assign o[59726] = i[116];
  assign o[59727] = i[116];
  assign o[59728] = i[116];
  assign o[59729] = i[116];
  assign o[59730] = i[116];
  assign o[59731] = i[116];
  assign o[59732] = i[116];
  assign o[59733] = i[116];
  assign o[59734] = i[116];
  assign o[59735] = i[116];
  assign o[59736] = i[116];
  assign o[59737] = i[116];
  assign o[59738] = i[116];
  assign o[59739] = i[116];
  assign o[59740] = i[116];
  assign o[59741] = i[116];
  assign o[59742] = i[116];
  assign o[59743] = i[116];
  assign o[59744] = i[116];
  assign o[59745] = i[116];
  assign o[59746] = i[116];
  assign o[59747] = i[116];
  assign o[59748] = i[116];
  assign o[59749] = i[116];
  assign o[59750] = i[116];
  assign o[59751] = i[116];
  assign o[59752] = i[116];
  assign o[59753] = i[116];
  assign o[59754] = i[116];
  assign o[59755] = i[116];
  assign o[59756] = i[116];
  assign o[59757] = i[116];
  assign o[59758] = i[116];
  assign o[59759] = i[116];
  assign o[59760] = i[116];
  assign o[59761] = i[116];
  assign o[59762] = i[116];
  assign o[59763] = i[116];
  assign o[59764] = i[116];
  assign o[59765] = i[116];
  assign o[59766] = i[116];
  assign o[59767] = i[116];
  assign o[59768] = i[116];
  assign o[59769] = i[116];
  assign o[59770] = i[116];
  assign o[59771] = i[116];
  assign o[59772] = i[116];
  assign o[59773] = i[116];
  assign o[59774] = i[116];
  assign o[59775] = i[116];
  assign o[59776] = i[116];
  assign o[59777] = i[116];
  assign o[59778] = i[116];
  assign o[59779] = i[116];
  assign o[59780] = i[116];
  assign o[59781] = i[116];
  assign o[59782] = i[116];
  assign o[59783] = i[116];
  assign o[59784] = i[116];
  assign o[59785] = i[116];
  assign o[59786] = i[116];
  assign o[59787] = i[116];
  assign o[59788] = i[116];
  assign o[59789] = i[116];
  assign o[59790] = i[116];
  assign o[59791] = i[116];
  assign o[59792] = i[116];
  assign o[59793] = i[116];
  assign o[59794] = i[116];
  assign o[59795] = i[116];
  assign o[59796] = i[116];
  assign o[59797] = i[116];
  assign o[59798] = i[116];
  assign o[59799] = i[116];
  assign o[59800] = i[116];
  assign o[59801] = i[116];
  assign o[59802] = i[116];
  assign o[59803] = i[116];
  assign o[59804] = i[116];
  assign o[59805] = i[116];
  assign o[59806] = i[116];
  assign o[59807] = i[116];
  assign o[59808] = i[116];
  assign o[59809] = i[116];
  assign o[59810] = i[116];
  assign o[59811] = i[116];
  assign o[59812] = i[116];
  assign o[59813] = i[116];
  assign o[59814] = i[116];
  assign o[59815] = i[116];
  assign o[59816] = i[116];
  assign o[59817] = i[116];
  assign o[59818] = i[116];
  assign o[59819] = i[116];
  assign o[59820] = i[116];
  assign o[59821] = i[116];
  assign o[59822] = i[116];
  assign o[59823] = i[116];
  assign o[59824] = i[116];
  assign o[59825] = i[116];
  assign o[59826] = i[116];
  assign o[59827] = i[116];
  assign o[59828] = i[116];
  assign o[59829] = i[116];
  assign o[59830] = i[116];
  assign o[59831] = i[116];
  assign o[59832] = i[116];
  assign o[59833] = i[116];
  assign o[59834] = i[116];
  assign o[59835] = i[116];
  assign o[59836] = i[116];
  assign o[59837] = i[116];
  assign o[59838] = i[116];
  assign o[59839] = i[116];
  assign o[59840] = i[116];
  assign o[59841] = i[116];
  assign o[59842] = i[116];
  assign o[59843] = i[116];
  assign o[59844] = i[116];
  assign o[59845] = i[116];
  assign o[59846] = i[116];
  assign o[59847] = i[116];
  assign o[59848] = i[116];
  assign o[59849] = i[116];
  assign o[59850] = i[116];
  assign o[59851] = i[116];
  assign o[59852] = i[116];
  assign o[59853] = i[116];
  assign o[59854] = i[116];
  assign o[59855] = i[116];
  assign o[59856] = i[116];
  assign o[59857] = i[116];
  assign o[59858] = i[116];
  assign o[59859] = i[116];
  assign o[59860] = i[116];
  assign o[59861] = i[116];
  assign o[59862] = i[116];
  assign o[59863] = i[116];
  assign o[59864] = i[116];
  assign o[59865] = i[116];
  assign o[59866] = i[116];
  assign o[59867] = i[116];
  assign o[59868] = i[116];
  assign o[59869] = i[116];
  assign o[59870] = i[116];
  assign o[59871] = i[116];
  assign o[59872] = i[116];
  assign o[59873] = i[116];
  assign o[59874] = i[116];
  assign o[59875] = i[116];
  assign o[59876] = i[116];
  assign o[59877] = i[116];
  assign o[59878] = i[116];
  assign o[59879] = i[116];
  assign o[59880] = i[116];
  assign o[59881] = i[116];
  assign o[59882] = i[116];
  assign o[59883] = i[116];
  assign o[59884] = i[116];
  assign o[59885] = i[116];
  assign o[59886] = i[116];
  assign o[59887] = i[116];
  assign o[59888] = i[116];
  assign o[59889] = i[116];
  assign o[59890] = i[116];
  assign o[59891] = i[116];
  assign o[59892] = i[116];
  assign o[59893] = i[116];
  assign o[59894] = i[116];
  assign o[59895] = i[116];
  assign o[59896] = i[116];
  assign o[59897] = i[116];
  assign o[59898] = i[116];
  assign o[59899] = i[116];
  assign o[59900] = i[116];
  assign o[59901] = i[116];
  assign o[59902] = i[116];
  assign o[59903] = i[116];
  assign o[58880] = i[115];
  assign o[58881] = i[115];
  assign o[58882] = i[115];
  assign o[58883] = i[115];
  assign o[58884] = i[115];
  assign o[58885] = i[115];
  assign o[58886] = i[115];
  assign o[58887] = i[115];
  assign o[58888] = i[115];
  assign o[58889] = i[115];
  assign o[58890] = i[115];
  assign o[58891] = i[115];
  assign o[58892] = i[115];
  assign o[58893] = i[115];
  assign o[58894] = i[115];
  assign o[58895] = i[115];
  assign o[58896] = i[115];
  assign o[58897] = i[115];
  assign o[58898] = i[115];
  assign o[58899] = i[115];
  assign o[58900] = i[115];
  assign o[58901] = i[115];
  assign o[58902] = i[115];
  assign o[58903] = i[115];
  assign o[58904] = i[115];
  assign o[58905] = i[115];
  assign o[58906] = i[115];
  assign o[58907] = i[115];
  assign o[58908] = i[115];
  assign o[58909] = i[115];
  assign o[58910] = i[115];
  assign o[58911] = i[115];
  assign o[58912] = i[115];
  assign o[58913] = i[115];
  assign o[58914] = i[115];
  assign o[58915] = i[115];
  assign o[58916] = i[115];
  assign o[58917] = i[115];
  assign o[58918] = i[115];
  assign o[58919] = i[115];
  assign o[58920] = i[115];
  assign o[58921] = i[115];
  assign o[58922] = i[115];
  assign o[58923] = i[115];
  assign o[58924] = i[115];
  assign o[58925] = i[115];
  assign o[58926] = i[115];
  assign o[58927] = i[115];
  assign o[58928] = i[115];
  assign o[58929] = i[115];
  assign o[58930] = i[115];
  assign o[58931] = i[115];
  assign o[58932] = i[115];
  assign o[58933] = i[115];
  assign o[58934] = i[115];
  assign o[58935] = i[115];
  assign o[58936] = i[115];
  assign o[58937] = i[115];
  assign o[58938] = i[115];
  assign o[58939] = i[115];
  assign o[58940] = i[115];
  assign o[58941] = i[115];
  assign o[58942] = i[115];
  assign o[58943] = i[115];
  assign o[58944] = i[115];
  assign o[58945] = i[115];
  assign o[58946] = i[115];
  assign o[58947] = i[115];
  assign o[58948] = i[115];
  assign o[58949] = i[115];
  assign o[58950] = i[115];
  assign o[58951] = i[115];
  assign o[58952] = i[115];
  assign o[58953] = i[115];
  assign o[58954] = i[115];
  assign o[58955] = i[115];
  assign o[58956] = i[115];
  assign o[58957] = i[115];
  assign o[58958] = i[115];
  assign o[58959] = i[115];
  assign o[58960] = i[115];
  assign o[58961] = i[115];
  assign o[58962] = i[115];
  assign o[58963] = i[115];
  assign o[58964] = i[115];
  assign o[58965] = i[115];
  assign o[58966] = i[115];
  assign o[58967] = i[115];
  assign o[58968] = i[115];
  assign o[58969] = i[115];
  assign o[58970] = i[115];
  assign o[58971] = i[115];
  assign o[58972] = i[115];
  assign o[58973] = i[115];
  assign o[58974] = i[115];
  assign o[58975] = i[115];
  assign o[58976] = i[115];
  assign o[58977] = i[115];
  assign o[58978] = i[115];
  assign o[58979] = i[115];
  assign o[58980] = i[115];
  assign o[58981] = i[115];
  assign o[58982] = i[115];
  assign o[58983] = i[115];
  assign o[58984] = i[115];
  assign o[58985] = i[115];
  assign o[58986] = i[115];
  assign o[58987] = i[115];
  assign o[58988] = i[115];
  assign o[58989] = i[115];
  assign o[58990] = i[115];
  assign o[58991] = i[115];
  assign o[58992] = i[115];
  assign o[58993] = i[115];
  assign o[58994] = i[115];
  assign o[58995] = i[115];
  assign o[58996] = i[115];
  assign o[58997] = i[115];
  assign o[58998] = i[115];
  assign o[58999] = i[115];
  assign o[59000] = i[115];
  assign o[59001] = i[115];
  assign o[59002] = i[115];
  assign o[59003] = i[115];
  assign o[59004] = i[115];
  assign o[59005] = i[115];
  assign o[59006] = i[115];
  assign o[59007] = i[115];
  assign o[59008] = i[115];
  assign o[59009] = i[115];
  assign o[59010] = i[115];
  assign o[59011] = i[115];
  assign o[59012] = i[115];
  assign o[59013] = i[115];
  assign o[59014] = i[115];
  assign o[59015] = i[115];
  assign o[59016] = i[115];
  assign o[59017] = i[115];
  assign o[59018] = i[115];
  assign o[59019] = i[115];
  assign o[59020] = i[115];
  assign o[59021] = i[115];
  assign o[59022] = i[115];
  assign o[59023] = i[115];
  assign o[59024] = i[115];
  assign o[59025] = i[115];
  assign o[59026] = i[115];
  assign o[59027] = i[115];
  assign o[59028] = i[115];
  assign o[59029] = i[115];
  assign o[59030] = i[115];
  assign o[59031] = i[115];
  assign o[59032] = i[115];
  assign o[59033] = i[115];
  assign o[59034] = i[115];
  assign o[59035] = i[115];
  assign o[59036] = i[115];
  assign o[59037] = i[115];
  assign o[59038] = i[115];
  assign o[59039] = i[115];
  assign o[59040] = i[115];
  assign o[59041] = i[115];
  assign o[59042] = i[115];
  assign o[59043] = i[115];
  assign o[59044] = i[115];
  assign o[59045] = i[115];
  assign o[59046] = i[115];
  assign o[59047] = i[115];
  assign o[59048] = i[115];
  assign o[59049] = i[115];
  assign o[59050] = i[115];
  assign o[59051] = i[115];
  assign o[59052] = i[115];
  assign o[59053] = i[115];
  assign o[59054] = i[115];
  assign o[59055] = i[115];
  assign o[59056] = i[115];
  assign o[59057] = i[115];
  assign o[59058] = i[115];
  assign o[59059] = i[115];
  assign o[59060] = i[115];
  assign o[59061] = i[115];
  assign o[59062] = i[115];
  assign o[59063] = i[115];
  assign o[59064] = i[115];
  assign o[59065] = i[115];
  assign o[59066] = i[115];
  assign o[59067] = i[115];
  assign o[59068] = i[115];
  assign o[59069] = i[115];
  assign o[59070] = i[115];
  assign o[59071] = i[115];
  assign o[59072] = i[115];
  assign o[59073] = i[115];
  assign o[59074] = i[115];
  assign o[59075] = i[115];
  assign o[59076] = i[115];
  assign o[59077] = i[115];
  assign o[59078] = i[115];
  assign o[59079] = i[115];
  assign o[59080] = i[115];
  assign o[59081] = i[115];
  assign o[59082] = i[115];
  assign o[59083] = i[115];
  assign o[59084] = i[115];
  assign o[59085] = i[115];
  assign o[59086] = i[115];
  assign o[59087] = i[115];
  assign o[59088] = i[115];
  assign o[59089] = i[115];
  assign o[59090] = i[115];
  assign o[59091] = i[115];
  assign o[59092] = i[115];
  assign o[59093] = i[115];
  assign o[59094] = i[115];
  assign o[59095] = i[115];
  assign o[59096] = i[115];
  assign o[59097] = i[115];
  assign o[59098] = i[115];
  assign o[59099] = i[115];
  assign o[59100] = i[115];
  assign o[59101] = i[115];
  assign o[59102] = i[115];
  assign o[59103] = i[115];
  assign o[59104] = i[115];
  assign o[59105] = i[115];
  assign o[59106] = i[115];
  assign o[59107] = i[115];
  assign o[59108] = i[115];
  assign o[59109] = i[115];
  assign o[59110] = i[115];
  assign o[59111] = i[115];
  assign o[59112] = i[115];
  assign o[59113] = i[115];
  assign o[59114] = i[115];
  assign o[59115] = i[115];
  assign o[59116] = i[115];
  assign o[59117] = i[115];
  assign o[59118] = i[115];
  assign o[59119] = i[115];
  assign o[59120] = i[115];
  assign o[59121] = i[115];
  assign o[59122] = i[115];
  assign o[59123] = i[115];
  assign o[59124] = i[115];
  assign o[59125] = i[115];
  assign o[59126] = i[115];
  assign o[59127] = i[115];
  assign o[59128] = i[115];
  assign o[59129] = i[115];
  assign o[59130] = i[115];
  assign o[59131] = i[115];
  assign o[59132] = i[115];
  assign o[59133] = i[115];
  assign o[59134] = i[115];
  assign o[59135] = i[115];
  assign o[59136] = i[115];
  assign o[59137] = i[115];
  assign o[59138] = i[115];
  assign o[59139] = i[115];
  assign o[59140] = i[115];
  assign o[59141] = i[115];
  assign o[59142] = i[115];
  assign o[59143] = i[115];
  assign o[59144] = i[115];
  assign o[59145] = i[115];
  assign o[59146] = i[115];
  assign o[59147] = i[115];
  assign o[59148] = i[115];
  assign o[59149] = i[115];
  assign o[59150] = i[115];
  assign o[59151] = i[115];
  assign o[59152] = i[115];
  assign o[59153] = i[115];
  assign o[59154] = i[115];
  assign o[59155] = i[115];
  assign o[59156] = i[115];
  assign o[59157] = i[115];
  assign o[59158] = i[115];
  assign o[59159] = i[115];
  assign o[59160] = i[115];
  assign o[59161] = i[115];
  assign o[59162] = i[115];
  assign o[59163] = i[115];
  assign o[59164] = i[115];
  assign o[59165] = i[115];
  assign o[59166] = i[115];
  assign o[59167] = i[115];
  assign o[59168] = i[115];
  assign o[59169] = i[115];
  assign o[59170] = i[115];
  assign o[59171] = i[115];
  assign o[59172] = i[115];
  assign o[59173] = i[115];
  assign o[59174] = i[115];
  assign o[59175] = i[115];
  assign o[59176] = i[115];
  assign o[59177] = i[115];
  assign o[59178] = i[115];
  assign o[59179] = i[115];
  assign o[59180] = i[115];
  assign o[59181] = i[115];
  assign o[59182] = i[115];
  assign o[59183] = i[115];
  assign o[59184] = i[115];
  assign o[59185] = i[115];
  assign o[59186] = i[115];
  assign o[59187] = i[115];
  assign o[59188] = i[115];
  assign o[59189] = i[115];
  assign o[59190] = i[115];
  assign o[59191] = i[115];
  assign o[59192] = i[115];
  assign o[59193] = i[115];
  assign o[59194] = i[115];
  assign o[59195] = i[115];
  assign o[59196] = i[115];
  assign o[59197] = i[115];
  assign o[59198] = i[115];
  assign o[59199] = i[115];
  assign o[59200] = i[115];
  assign o[59201] = i[115];
  assign o[59202] = i[115];
  assign o[59203] = i[115];
  assign o[59204] = i[115];
  assign o[59205] = i[115];
  assign o[59206] = i[115];
  assign o[59207] = i[115];
  assign o[59208] = i[115];
  assign o[59209] = i[115];
  assign o[59210] = i[115];
  assign o[59211] = i[115];
  assign o[59212] = i[115];
  assign o[59213] = i[115];
  assign o[59214] = i[115];
  assign o[59215] = i[115];
  assign o[59216] = i[115];
  assign o[59217] = i[115];
  assign o[59218] = i[115];
  assign o[59219] = i[115];
  assign o[59220] = i[115];
  assign o[59221] = i[115];
  assign o[59222] = i[115];
  assign o[59223] = i[115];
  assign o[59224] = i[115];
  assign o[59225] = i[115];
  assign o[59226] = i[115];
  assign o[59227] = i[115];
  assign o[59228] = i[115];
  assign o[59229] = i[115];
  assign o[59230] = i[115];
  assign o[59231] = i[115];
  assign o[59232] = i[115];
  assign o[59233] = i[115];
  assign o[59234] = i[115];
  assign o[59235] = i[115];
  assign o[59236] = i[115];
  assign o[59237] = i[115];
  assign o[59238] = i[115];
  assign o[59239] = i[115];
  assign o[59240] = i[115];
  assign o[59241] = i[115];
  assign o[59242] = i[115];
  assign o[59243] = i[115];
  assign o[59244] = i[115];
  assign o[59245] = i[115];
  assign o[59246] = i[115];
  assign o[59247] = i[115];
  assign o[59248] = i[115];
  assign o[59249] = i[115];
  assign o[59250] = i[115];
  assign o[59251] = i[115];
  assign o[59252] = i[115];
  assign o[59253] = i[115];
  assign o[59254] = i[115];
  assign o[59255] = i[115];
  assign o[59256] = i[115];
  assign o[59257] = i[115];
  assign o[59258] = i[115];
  assign o[59259] = i[115];
  assign o[59260] = i[115];
  assign o[59261] = i[115];
  assign o[59262] = i[115];
  assign o[59263] = i[115];
  assign o[59264] = i[115];
  assign o[59265] = i[115];
  assign o[59266] = i[115];
  assign o[59267] = i[115];
  assign o[59268] = i[115];
  assign o[59269] = i[115];
  assign o[59270] = i[115];
  assign o[59271] = i[115];
  assign o[59272] = i[115];
  assign o[59273] = i[115];
  assign o[59274] = i[115];
  assign o[59275] = i[115];
  assign o[59276] = i[115];
  assign o[59277] = i[115];
  assign o[59278] = i[115];
  assign o[59279] = i[115];
  assign o[59280] = i[115];
  assign o[59281] = i[115];
  assign o[59282] = i[115];
  assign o[59283] = i[115];
  assign o[59284] = i[115];
  assign o[59285] = i[115];
  assign o[59286] = i[115];
  assign o[59287] = i[115];
  assign o[59288] = i[115];
  assign o[59289] = i[115];
  assign o[59290] = i[115];
  assign o[59291] = i[115];
  assign o[59292] = i[115];
  assign o[59293] = i[115];
  assign o[59294] = i[115];
  assign o[59295] = i[115];
  assign o[59296] = i[115];
  assign o[59297] = i[115];
  assign o[59298] = i[115];
  assign o[59299] = i[115];
  assign o[59300] = i[115];
  assign o[59301] = i[115];
  assign o[59302] = i[115];
  assign o[59303] = i[115];
  assign o[59304] = i[115];
  assign o[59305] = i[115];
  assign o[59306] = i[115];
  assign o[59307] = i[115];
  assign o[59308] = i[115];
  assign o[59309] = i[115];
  assign o[59310] = i[115];
  assign o[59311] = i[115];
  assign o[59312] = i[115];
  assign o[59313] = i[115];
  assign o[59314] = i[115];
  assign o[59315] = i[115];
  assign o[59316] = i[115];
  assign o[59317] = i[115];
  assign o[59318] = i[115];
  assign o[59319] = i[115];
  assign o[59320] = i[115];
  assign o[59321] = i[115];
  assign o[59322] = i[115];
  assign o[59323] = i[115];
  assign o[59324] = i[115];
  assign o[59325] = i[115];
  assign o[59326] = i[115];
  assign o[59327] = i[115];
  assign o[59328] = i[115];
  assign o[59329] = i[115];
  assign o[59330] = i[115];
  assign o[59331] = i[115];
  assign o[59332] = i[115];
  assign o[59333] = i[115];
  assign o[59334] = i[115];
  assign o[59335] = i[115];
  assign o[59336] = i[115];
  assign o[59337] = i[115];
  assign o[59338] = i[115];
  assign o[59339] = i[115];
  assign o[59340] = i[115];
  assign o[59341] = i[115];
  assign o[59342] = i[115];
  assign o[59343] = i[115];
  assign o[59344] = i[115];
  assign o[59345] = i[115];
  assign o[59346] = i[115];
  assign o[59347] = i[115];
  assign o[59348] = i[115];
  assign o[59349] = i[115];
  assign o[59350] = i[115];
  assign o[59351] = i[115];
  assign o[59352] = i[115];
  assign o[59353] = i[115];
  assign o[59354] = i[115];
  assign o[59355] = i[115];
  assign o[59356] = i[115];
  assign o[59357] = i[115];
  assign o[59358] = i[115];
  assign o[59359] = i[115];
  assign o[59360] = i[115];
  assign o[59361] = i[115];
  assign o[59362] = i[115];
  assign o[59363] = i[115];
  assign o[59364] = i[115];
  assign o[59365] = i[115];
  assign o[59366] = i[115];
  assign o[59367] = i[115];
  assign o[59368] = i[115];
  assign o[59369] = i[115];
  assign o[59370] = i[115];
  assign o[59371] = i[115];
  assign o[59372] = i[115];
  assign o[59373] = i[115];
  assign o[59374] = i[115];
  assign o[59375] = i[115];
  assign o[59376] = i[115];
  assign o[59377] = i[115];
  assign o[59378] = i[115];
  assign o[59379] = i[115];
  assign o[59380] = i[115];
  assign o[59381] = i[115];
  assign o[59382] = i[115];
  assign o[59383] = i[115];
  assign o[59384] = i[115];
  assign o[59385] = i[115];
  assign o[59386] = i[115];
  assign o[59387] = i[115];
  assign o[59388] = i[115];
  assign o[59389] = i[115];
  assign o[59390] = i[115];
  assign o[59391] = i[115];
  assign o[58368] = i[114];
  assign o[58369] = i[114];
  assign o[58370] = i[114];
  assign o[58371] = i[114];
  assign o[58372] = i[114];
  assign o[58373] = i[114];
  assign o[58374] = i[114];
  assign o[58375] = i[114];
  assign o[58376] = i[114];
  assign o[58377] = i[114];
  assign o[58378] = i[114];
  assign o[58379] = i[114];
  assign o[58380] = i[114];
  assign o[58381] = i[114];
  assign o[58382] = i[114];
  assign o[58383] = i[114];
  assign o[58384] = i[114];
  assign o[58385] = i[114];
  assign o[58386] = i[114];
  assign o[58387] = i[114];
  assign o[58388] = i[114];
  assign o[58389] = i[114];
  assign o[58390] = i[114];
  assign o[58391] = i[114];
  assign o[58392] = i[114];
  assign o[58393] = i[114];
  assign o[58394] = i[114];
  assign o[58395] = i[114];
  assign o[58396] = i[114];
  assign o[58397] = i[114];
  assign o[58398] = i[114];
  assign o[58399] = i[114];
  assign o[58400] = i[114];
  assign o[58401] = i[114];
  assign o[58402] = i[114];
  assign o[58403] = i[114];
  assign o[58404] = i[114];
  assign o[58405] = i[114];
  assign o[58406] = i[114];
  assign o[58407] = i[114];
  assign o[58408] = i[114];
  assign o[58409] = i[114];
  assign o[58410] = i[114];
  assign o[58411] = i[114];
  assign o[58412] = i[114];
  assign o[58413] = i[114];
  assign o[58414] = i[114];
  assign o[58415] = i[114];
  assign o[58416] = i[114];
  assign o[58417] = i[114];
  assign o[58418] = i[114];
  assign o[58419] = i[114];
  assign o[58420] = i[114];
  assign o[58421] = i[114];
  assign o[58422] = i[114];
  assign o[58423] = i[114];
  assign o[58424] = i[114];
  assign o[58425] = i[114];
  assign o[58426] = i[114];
  assign o[58427] = i[114];
  assign o[58428] = i[114];
  assign o[58429] = i[114];
  assign o[58430] = i[114];
  assign o[58431] = i[114];
  assign o[58432] = i[114];
  assign o[58433] = i[114];
  assign o[58434] = i[114];
  assign o[58435] = i[114];
  assign o[58436] = i[114];
  assign o[58437] = i[114];
  assign o[58438] = i[114];
  assign o[58439] = i[114];
  assign o[58440] = i[114];
  assign o[58441] = i[114];
  assign o[58442] = i[114];
  assign o[58443] = i[114];
  assign o[58444] = i[114];
  assign o[58445] = i[114];
  assign o[58446] = i[114];
  assign o[58447] = i[114];
  assign o[58448] = i[114];
  assign o[58449] = i[114];
  assign o[58450] = i[114];
  assign o[58451] = i[114];
  assign o[58452] = i[114];
  assign o[58453] = i[114];
  assign o[58454] = i[114];
  assign o[58455] = i[114];
  assign o[58456] = i[114];
  assign o[58457] = i[114];
  assign o[58458] = i[114];
  assign o[58459] = i[114];
  assign o[58460] = i[114];
  assign o[58461] = i[114];
  assign o[58462] = i[114];
  assign o[58463] = i[114];
  assign o[58464] = i[114];
  assign o[58465] = i[114];
  assign o[58466] = i[114];
  assign o[58467] = i[114];
  assign o[58468] = i[114];
  assign o[58469] = i[114];
  assign o[58470] = i[114];
  assign o[58471] = i[114];
  assign o[58472] = i[114];
  assign o[58473] = i[114];
  assign o[58474] = i[114];
  assign o[58475] = i[114];
  assign o[58476] = i[114];
  assign o[58477] = i[114];
  assign o[58478] = i[114];
  assign o[58479] = i[114];
  assign o[58480] = i[114];
  assign o[58481] = i[114];
  assign o[58482] = i[114];
  assign o[58483] = i[114];
  assign o[58484] = i[114];
  assign o[58485] = i[114];
  assign o[58486] = i[114];
  assign o[58487] = i[114];
  assign o[58488] = i[114];
  assign o[58489] = i[114];
  assign o[58490] = i[114];
  assign o[58491] = i[114];
  assign o[58492] = i[114];
  assign o[58493] = i[114];
  assign o[58494] = i[114];
  assign o[58495] = i[114];
  assign o[58496] = i[114];
  assign o[58497] = i[114];
  assign o[58498] = i[114];
  assign o[58499] = i[114];
  assign o[58500] = i[114];
  assign o[58501] = i[114];
  assign o[58502] = i[114];
  assign o[58503] = i[114];
  assign o[58504] = i[114];
  assign o[58505] = i[114];
  assign o[58506] = i[114];
  assign o[58507] = i[114];
  assign o[58508] = i[114];
  assign o[58509] = i[114];
  assign o[58510] = i[114];
  assign o[58511] = i[114];
  assign o[58512] = i[114];
  assign o[58513] = i[114];
  assign o[58514] = i[114];
  assign o[58515] = i[114];
  assign o[58516] = i[114];
  assign o[58517] = i[114];
  assign o[58518] = i[114];
  assign o[58519] = i[114];
  assign o[58520] = i[114];
  assign o[58521] = i[114];
  assign o[58522] = i[114];
  assign o[58523] = i[114];
  assign o[58524] = i[114];
  assign o[58525] = i[114];
  assign o[58526] = i[114];
  assign o[58527] = i[114];
  assign o[58528] = i[114];
  assign o[58529] = i[114];
  assign o[58530] = i[114];
  assign o[58531] = i[114];
  assign o[58532] = i[114];
  assign o[58533] = i[114];
  assign o[58534] = i[114];
  assign o[58535] = i[114];
  assign o[58536] = i[114];
  assign o[58537] = i[114];
  assign o[58538] = i[114];
  assign o[58539] = i[114];
  assign o[58540] = i[114];
  assign o[58541] = i[114];
  assign o[58542] = i[114];
  assign o[58543] = i[114];
  assign o[58544] = i[114];
  assign o[58545] = i[114];
  assign o[58546] = i[114];
  assign o[58547] = i[114];
  assign o[58548] = i[114];
  assign o[58549] = i[114];
  assign o[58550] = i[114];
  assign o[58551] = i[114];
  assign o[58552] = i[114];
  assign o[58553] = i[114];
  assign o[58554] = i[114];
  assign o[58555] = i[114];
  assign o[58556] = i[114];
  assign o[58557] = i[114];
  assign o[58558] = i[114];
  assign o[58559] = i[114];
  assign o[58560] = i[114];
  assign o[58561] = i[114];
  assign o[58562] = i[114];
  assign o[58563] = i[114];
  assign o[58564] = i[114];
  assign o[58565] = i[114];
  assign o[58566] = i[114];
  assign o[58567] = i[114];
  assign o[58568] = i[114];
  assign o[58569] = i[114];
  assign o[58570] = i[114];
  assign o[58571] = i[114];
  assign o[58572] = i[114];
  assign o[58573] = i[114];
  assign o[58574] = i[114];
  assign o[58575] = i[114];
  assign o[58576] = i[114];
  assign o[58577] = i[114];
  assign o[58578] = i[114];
  assign o[58579] = i[114];
  assign o[58580] = i[114];
  assign o[58581] = i[114];
  assign o[58582] = i[114];
  assign o[58583] = i[114];
  assign o[58584] = i[114];
  assign o[58585] = i[114];
  assign o[58586] = i[114];
  assign o[58587] = i[114];
  assign o[58588] = i[114];
  assign o[58589] = i[114];
  assign o[58590] = i[114];
  assign o[58591] = i[114];
  assign o[58592] = i[114];
  assign o[58593] = i[114];
  assign o[58594] = i[114];
  assign o[58595] = i[114];
  assign o[58596] = i[114];
  assign o[58597] = i[114];
  assign o[58598] = i[114];
  assign o[58599] = i[114];
  assign o[58600] = i[114];
  assign o[58601] = i[114];
  assign o[58602] = i[114];
  assign o[58603] = i[114];
  assign o[58604] = i[114];
  assign o[58605] = i[114];
  assign o[58606] = i[114];
  assign o[58607] = i[114];
  assign o[58608] = i[114];
  assign o[58609] = i[114];
  assign o[58610] = i[114];
  assign o[58611] = i[114];
  assign o[58612] = i[114];
  assign o[58613] = i[114];
  assign o[58614] = i[114];
  assign o[58615] = i[114];
  assign o[58616] = i[114];
  assign o[58617] = i[114];
  assign o[58618] = i[114];
  assign o[58619] = i[114];
  assign o[58620] = i[114];
  assign o[58621] = i[114];
  assign o[58622] = i[114];
  assign o[58623] = i[114];
  assign o[58624] = i[114];
  assign o[58625] = i[114];
  assign o[58626] = i[114];
  assign o[58627] = i[114];
  assign o[58628] = i[114];
  assign o[58629] = i[114];
  assign o[58630] = i[114];
  assign o[58631] = i[114];
  assign o[58632] = i[114];
  assign o[58633] = i[114];
  assign o[58634] = i[114];
  assign o[58635] = i[114];
  assign o[58636] = i[114];
  assign o[58637] = i[114];
  assign o[58638] = i[114];
  assign o[58639] = i[114];
  assign o[58640] = i[114];
  assign o[58641] = i[114];
  assign o[58642] = i[114];
  assign o[58643] = i[114];
  assign o[58644] = i[114];
  assign o[58645] = i[114];
  assign o[58646] = i[114];
  assign o[58647] = i[114];
  assign o[58648] = i[114];
  assign o[58649] = i[114];
  assign o[58650] = i[114];
  assign o[58651] = i[114];
  assign o[58652] = i[114];
  assign o[58653] = i[114];
  assign o[58654] = i[114];
  assign o[58655] = i[114];
  assign o[58656] = i[114];
  assign o[58657] = i[114];
  assign o[58658] = i[114];
  assign o[58659] = i[114];
  assign o[58660] = i[114];
  assign o[58661] = i[114];
  assign o[58662] = i[114];
  assign o[58663] = i[114];
  assign o[58664] = i[114];
  assign o[58665] = i[114];
  assign o[58666] = i[114];
  assign o[58667] = i[114];
  assign o[58668] = i[114];
  assign o[58669] = i[114];
  assign o[58670] = i[114];
  assign o[58671] = i[114];
  assign o[58672] = i[114];
  assign o[58673] = i[114];
  assign o[58674] = i[114];
  assign o[58675] = i[114];
  assign o[58676] = i[114];
  assign o[58677] = i[114];
  assign o[58678] = i[114];
  assign o[58679] = i[114];
  assign o[58680] = i[114];
  assign o[58681] = i[114];
  assign o[58682] = i[114];
  assign o[58683] = i[114];
  assign o[58684] = i[114];
  assign o[58685] = i[114];
  assign o[58686] = i[114];
  assign o[58687] = i[114];
  assign o[58688] = i[114];
  assign o[58689] = i[114];
  assign o[58690] = i[114];
  assign o[58691] = i[114];
  assign o[58692] = i[114];
  assign o[58693] = i[114];
  assign o[58694] = i[114];
  assign o[58695] = i[114];
  assign o[58696] = i[114];
  assign o[58697] = i[114];
  assign o[58698] = i[114];
  assign o[58699] = i[114];
  assign o[58700] = i[114];
  assign o[58701] = i[114];
  assign o[58702] = i[114];
  assign o[58703] = i[114];
  assign o[58704] = i[114];
  assign o[58705] = i[114];
  assign o[58706] = i[114];
  assign o[58707] = i[114];
  assign o[58708] = i[114];
  assign o[58709] = i[114];
  assign o[58710] = i[114];
  assign o[58711] = i[114];
  assign o[58712] = i[114];
  assign o[58713] = i[114];
  assign o[58714] = i[114];
  assign o[58715] = i[114];
  assign o[58716] = i[114];
  assign o[58717] = i[114];
  assign o[58718] = i[114];
  assign o[58719] = i[114];
  assign o[58720] = i[114];
  assign o[58721] = i[114];
  assign o[58722] = i[114];
  assign o[58723] = i[114];
  assign o[58724] = i[114];
  assign o[58725] = i[114];
  assign o[58726] = i[114];
  assign o[58727] = i[114];
  assign o[58728] = i[114];
  assign o[58729] = i[114];
  assign o[58730] = i[114];
  assign o[58731] = i[114];
  assign o[58732] = i[114];
  assign o[58733] = i[114];
  assign o[58734] = i[114];
  assign o[58735] = i[114];
  assign o[58736] = i[114];
  assign o[58737] = i[114];
  assign o[58738] = i[114];
  assign o[58739] = i[114];
  assign o[58740] = i[114];
  assign o[58741] = i[114];
  assign o[58742] = i[114];
  assign o[58743] = i[114];
  assign o[58744] = i[114];
  assign o[58745] = i[114];
  assign o[58746] = i[114];
  assign o[58747] = i[114];
  assign o[58748] = i[114];
  assign o[58749] = i[114];
  assign o[58750] = i[114];
  assign o[58751] = i[114];
  assign o[58752] = i[114];
  assign o[58753] = i[114];
  assign o[58754] = i[114];
  assign o[58755] = i[114];
  assign o[58756] = i[114];
  assign o[58757] = i[114];
  assign o[58758] = i[114];
  assign o[58759] = i[114];
  assign o[58760] = i[114];
  assign o[58761] = i[114];
  assign o[58762] = i[114];
  assign o[58763] = i[114];
  assign o[58764] = i[114];
  assign o[58765] = i[114];
  assign o[58766] = i[114];
  assign o[58767] = i[114];
  assign o[58768] = i[114];
  assign o[58769] = i[114];
  assign o[58770] = i[114];
  assign o[58771] = i[114];
  assign o[58772] = i[114];
  assign o[58773] = i[114];
  assign o[58774] = i[114];
  assign o[58775] = i[114];
  assign o[58776] = i[114];
  assign o[58777] = i[114];
  assign o[58778] = i[114];
  assign o[58779] = i[114];
  assign o[58780] = i[114];
  assign o[58781] = i[114];
  assign o[58782] = i[114];
  assign o[58783] = i[114];
  assign o[58784] = i[114];
  assign o[58785] = i[114];
  assign o[58786] = i[114];
  assign o[58787] = i[114];
  assign o[58788] = i[114];
  assign o[58789] = i[114];
  assign o[58790] = i[114];
  assign o[58791] = i[114];
  assign o[58792] = i[114];
  assign o[58793] = i[114];
  assign o[58794] = i[114];
  assign o[58795] = i[114];
  assign o[58796] = i[114];
  assign o[58797] = i[114];
  assign o[58798] = i[114];
  assign o[58799] = i[114];
  assign o[58800] = i[114];
  assign o[58801] = i[114];
  assign o[58802] = i[114];
  assign o[58803] = i[114];
  assign o[58804] = i[114];
  assign o[58805] = i[114];
  assign o[58806] = i[114];
  assign o[58807] = i[114];
  assign o[58808] = i[114];
  assign o[58809] = i[114];
  assign o[58810] = i[114];
  assign o[58811] = i[114];
  assign o[58812] = i[114];
  assign o[58813] = i[114];
  assign o[58814] = i[114];
  assign o[58815] = i[114];
  assign o[58816] = i[114];
  assign o[58817] = i[114];
  assign o[58818] = i[114];
  assign o[58819] = i[114];
  assign o[58820] = i[114];
  assign o[58821] = i[114];
  assign o[58822] = i[114];
  assign o[58823] = i[114];
  assign o[58824] = i[114];
  assign o[58825] = i[114];
  assign o[58826] = i[114];
  assign o[58827] = i[114];
  assign o[58828] = i[114];
  assign o[58829] = i[114];
  assign o[58830] = i[114];
  assign o[58831] = i[114];
  assign o[58832] = i[114];
  assign o[58833] = i[114];
  assign o[58834] = i[114];
  assign o[58835] = i[114];
  assign o[58836] = i[114];
  assign o[58837] = i[114];
  assign o[58838] = i[114];
  assign o[58839] = i[114];
  assign o[58840] = i[114];
  assign o[58841] = i[114];
  assign o[58842] = i[114];
  assign o[58843] = i[114];
  assign o[58844] = i[114];
  assign o[58845] = i[114];
  assign o[58846] = i[114];
  assign o[58847] = i[114];
  assign o[58848] = i[114];
  assign o[58849] = i[114];
  assign o[58850] = i[114];
  assign o[58851] = i[114];
  assign o[58852] = i[114];
  assign o[58853] = i[114];
  assign o[58854] = i[114];
  assign o[58855] = i[114];
  assign o[58856] = i[114];
  assign o[58857] = i[114];
  assign o[58858] = i[114];
  assign o[58859] = i[114];
  assign o[58860] = i[114];
  assign o[58861] = i[114];
  assign o[58862] = i[114];
  assign o[58863] = i[114];
  assign o[58864] = i[114];
  assign o[58865] = i[114];
  assign o[58866] = i[114];
  assign o[58867] = i[114];
  assign o[58868] = i[114];
  assign o[58869] = i[114];
  assign o[58870] = i[114];
  assign o[58871] = i[114];
  assign o[58872] = i[114];
  assign o[58873] = i[114];
  assign o[58874] = i[114];
  assign o[58875] = i[114];
  assign o[58876] = i[114];
  assign o[58877] = i[114];
  assign o[58878] = i[114];
  assign o[58879] = i[114];
  assign o[57856] = i[113];
  assign o[57857] = i[113];
  assign o[57858] = i[113];
  assign o[57859] = i[113];
  assign o[57860] = i[113];
  assign o[57861] = i[113];
  assign o[57862] = i[113];
  assign o[57863] = i[113];
  assign o[57864] = i[113];
  assign o[57865] = i[113];
  assign o[57866] = i[113];
  assign o[57867] = i[113];
  assign o[57868] = i[113];
  assign o[57869] = i[113];
  assign o[57870] = i[113];
  assign o[57871] = i[113];
  assign o[57872] = i[113];
  assign o[57873] = i[113];
  assign o[57874] = i[113];
  assign o[57875] = i[113];
  assign o[57876] = i[113];
  assign o[57877] = i[113];
  assign o[57878] = i[113];
  assign o[57879] = i[113];
  assign o[57880] = i[113];
  assign o[57881] = i[113];
  assign o[57882] = i[113];
  assign o[57883] = i[113];
  assign o[57884] = i[113];
  assign o[57885] = i[113];
  assign o[57886] = i[113];
  assign o[57887] = i[113];
  assign o[57888] = i[113];
  assign o[57889] = i[113];
  assign o[57890] = i[113];
  assign o[57891] = i[113];
  assign o[57892] = i[113];
  assign o[57893] = i[113];
  assign o[57894] = i[113];
  assign o[57895] = i[113];
  assign o[57896] = i[113];
  assign o[57897] = i[113];
  assign o[57898] = i[113];
  assign o[57899] = i[113];
  assign o[57900] = i[113];
  assign o[57901] = i[113];
  assign o[57902] = i[113];
  assign o[57903] = i[113];
  assign o[57904] = i[113];
  assign o[57905] = i[113];
  assign o[57906] = i[113];
  assign o[57907] = i[113];
  assign o[57908] = i[113];
  assign o[57909] = i[113];
  assign o[57910] = i[113];
  assign o[57911] = i[113];
  assign o[57912] = i[113];
  assign o[57913] = i[113];
  assign o[57914] = i[113];
  assign o[57915] = i[113];
  assign o[57916] = i[113];
  assign o[57917] = i[113];
  assign o[57918] = i[113];
  assign o[57919] = i[113];
  assign o[57920] = i[113];
  assign o[57921] = i[113];
  assign o[57922] = i[113];
  assign o[57923] = i[113];
  assign o[57924] = i[113];
  assign o[57925] = i[113];
  assign o[57926] = i[113];
  assign o[57927] = i[113];
  assign o[57928] = i[113];
  assign o[57929] = i[113];
  assign o[57930] = i[113];
  assign o[57931] = i[113];
  assign o[57932] = i[113];
  assign o[57933] = i[113];
  assign o[57934] = i[113];
  assign o[57935] = i[113];
  assign o[57936] = i[113];
  assign o[57937] = i[113];
  assign o[57938] = i[113];
  assign o[57939] = i[113];
  assign o[57940] = i[113];
  assign o[57941] = i[113];
  assign o[57942] = i[113];
  assign o[57943] = i[113];
  assign o[57944] = i[113];
  assign o[57945] = i[113];
  assign o[57946] = i[113];
  assign o[57947] = i[113];
  assign o[57948] = i[113];
  assign o[57949] = i[113];
  assign o[57950] = i[113];
  assign o[57951] = i[113];
  assign o[57952] = i[113];
  assign o[57953] = i[113];
  assign o[57954] = i[113];
  assign o[57955] = i[113];
  assign o[57956] = i[113];
  assign o[57957] = i[113];
  assign o[57958] = i[113];
  assign o[57959] = i[113];
  assign o[57960] = i[113];
  assign o[57961] = i[113];
  assign o[57962] = i[113];
  assign o[57963] = i[113];
  assign o[57964] = i[113];
  assign o[57965] = i[113];
  assign o[57966] = i[113];
  assign o[57967] = i[113];
  assign o[57968] = i[113];
  assign o[57969] = i[113];
  assign o[57970] = i[113];
  assign o[57971] = i[113];
  assign o[57972] = i[113];
  assign o[57973] = i[113];
  assign o[57974] = i[113];
  assign o[57975] = i[113];
  assign o[57976] = i[113];
  assign o[57977] = i[113];
  assign o[57978] = i[113];
  assign o[57979] = i[113];
  assign o[57980] = i[113];
  assign o[57981] = i[113];
  assign o[57982] = i[113];
  assign o[57983] = i[113];
  assign o[57984] = i[113];
  assign o[57985] = i[113];
  assign o[57986] = i[113];
  assign o[57987] = i[113];
  assign o[57988] = i[113];
  assign o[57989] = i[113];
  assign o[57990] = i[113];
  assign o[57991] = i[113];
  assign o[57992] = i[113];
  assign o[57993] = i[113];
  assign o[57994] = i[113];
  assign o[57995] = i[113];
  assign o[57996] = i[113];
  assign o[57997] = i[113];
  assign o[57998] = i[113];
  assign o[57999] = i[113];
  assign o[58000] = i[113];
  assign o[58001] = i[113];
  assign o[58002] = i[113];
  assign o[58003] = i[113];
  assign o[58004] = i[113];
  assign o[58005] = i[113];
  assign o[58006] = i[113];
  assign o[58007] = i[113];
  assign o[58008] = i[113];
  assign o[58009] = i[113];
  assign o[58010] = i[113];
  assign o[58011] = i[113];
  assign o[58012] = i[113];
  assign o[58013] = i[113];
  assign o[58014] = i[113];
  assign o[58015] = i[113];
  assign o[58016] = i[113];
  assign o[58017] = i[113];
  assign o[58018] = i[113];
  assign o[58019] = i[113];
  assign o[58020] = i[113];
  assign o[58021] = i[113];
  assign o[58022] = i[113];
  assign o[58023] = i[113];
  assign o[58024] = i[113];
  assign o[58025] = i[113];
  assign o[58026] = i[113];
  assign o[58027] = i[113];
  assign o[58028] = i[113];
  assign o[58029] = i[113];
  assign o[58030] = i[113];
  assign o[58031] = i[113];
  assign o[58032] = i[113];
  assign o[58033] = i[113];
  assign o[58034] = i[113];
  assign o[58035] = i[113];
  assign o[58036] = i[113];
  assign o[58037] = i[113];
  assign o[58038] = i[113];
  assign o[58039] = i[113];
  assign o[58040] = i[113];
  assign o[58041] = i[113];
  assign o[58042] = i[113];
  assign o[58043] = i[113];
  assign o[58044] = i[113];
  assign o[58045] = i[113];
  assign o[58046] = i[113];
  assign o[58047] = i[113];
  assign o[58048] = i[113];
  assign o[58049] = i[113];
  assign o[58050] = i[113];
  assign o[58051] = i[113];
  assign o[58052] = i[113];
  assign o[58053] = i[113];
  assign o[58054] = i[113];
  assign o[58055] = i[113];
  assign o[58056] = i[113];
  assign o[58057] = i[113];
  assign o[58058] = i[113];
  assign o[58059] = i[113];
  assign o[58060] = i[113];
  assign o[58061] = i[113];
  assign o[58062] = i[113];
  assign o[58063] = i[113];
  assign o[58064] = i[113];
  assign o[58065] = i[113];
  assign o[58066] = i[113];
  assign o[58067] = i[113];
  assign o[58068] = i[113];
  assign o[58069] = i[113];
  assign o[58070] = i[113];
  assign o[58071] = i[113];
  assign o[58072] = i[113];
  assign o[58073] = i[113];
  assign o[58074] = i[113];
  assign o[58075] = i[113];
  assign o[58076] = i[113];
  assign o[58077] = i[113];
  assign o[58078] = i[113];
  assign o[58079] = i[113];
  assign o[58080] = i[113];
  assign o[58081] = i[113];
  assign o[58082] = i[113];
  assign o[58083] = i[113];
  assign o[58084] = i[113];
  assign o[58085] = i[113];
  assign o[58086] = i[113];
  assign o[58087] = i[113];
  assign o[58088] = i[113];
  assign o[58089] = i[113];
  assign o[58090] = i[113];
  assign o[58091] = i[113];
  assign o[58092] = i[113];
  assign o[58093] = i[113];
  assign o[58094] = i[113];
  assign o[58095] = i[113];
  assign o[58096] = i[113];
  assign o[58097] = i[113];
  assign o[58098] = i[113];
  assign o[58099] = i[113];
  assign o[58100] = i[113];
  assign o[58101] = i[113];
  assign o[58102] = i[113];
  assign o[58103] = i[113];
  assign o[58104] = i[113];
  assign o[58105] = i[113];
  assign o[58106] = i[113];
  assign o[58107] = i[113];
  assign o[58108] = i[113];
  assign o[58109] = i[113];
  assign o[58110] = i[113];
  assign o[58111] = i[113];
  assign o[58112] = i[113];
  assign o[58113] = i[113];
  assign o[58114] = i[113];
  assign o[58115] = i[113];
  assign o[58116] = i[113];
  assign o[58117] = i[113];
  assign o[58118] = i[113];
  assign o[58119] = i[113];
  assign o[58120] = i[113];
  assign o[58121] = i[113];
  assign o[58122] = i[113];
  assign o[58123] = i[113];
  assign o[58124] = i[113];
  assign o[58125] = i[113];
  assign o[58126] = i[113];
  assign o[58127] = i[113];
  assign o[58128] = i[113];
  assign o[58129] = i[113];
  assign o[58130] = i[113];
  assign o[58131] = i[113];
  assign o[58132] = i[113];
  assign o[58133] = i[113];
  assign o[58134] = i[113];
  assign o[58135] = i[113];
  assign o[58136] = i[113];
  assign o[58137] = i[113];
  assign o[58138] = i[113];
  assign o[58139] = i[113];
  assign o[58140] = i[113];
  assign o[58141] = i[113];
  assign o[58142] = i[113];
  assign o[58143] = i[113];
  assign o[58144] = i[113];
  assign o[58145] = i[113];
  assign o[58146] = i[113];
  assign o[58147] = i[113];
  assign o[58148] = i[113];
  assign o[58149] = i[113];
  assign o[58150] = i[113];
  assign o[58151] = i[113];
  assign o[58152] = i[113];
  assign o[58153] = i[113];
  assign o[58154] = i[113];
  assign o[58155] = i[113];
  assign o[58156] = i[113];
  assign o[58157] = i[113];
  assign o[58158] = i[113];
  assign o[58159] = i[113];
  assign o[58160] = i[113];
  assign o[58161] = i[113];
  assign o[58162] = i[113];
  assign o[58163] = i[113];
  assign o[58164] = i[113];
  assign o[58165] = i[113];
  assign o[58166] = i[113];
  assign o[58167] = i[113];
  assign o[58168] = i[113];
  assign o[58169] = i[113];
  assign o[58170] = i[113];
  assign o[58171] = i[113];
  assign o[58172] = i[113];
  assign o[58173] = i[113];
  assign o[58174] = i[113];
  assign o[58175] = i[113];
  assign o[58176] = i[113];
  assign o[58177] = i[113];
  assign o[58178] = i[113];
  assign o[58179] = i[113];
  assign o[58180] = i[113];
  assign o[58181] = i[113];
  assign o[58182] = i[113];
  assign o[58183] = i[113];
  assign o[58184] = i[113];
  assign o[58185] = i[113];
  assign o[58186] = i[113];
  assign o[58187] = i[113];
  assign o[58188] = i[113];
  assign o[58189] = i[113];
  assign o[58190] = i[113];
  assign o[58191] = i[113];
  assign o[58192] = i[113];
  assign o[58193] = i[113];
  assign o[58194] = i[113];
  assign o[58195] = i[113];
  assign o[58196] = i[113];
  assign o[58197] = i[113];
  assign o[58198] = i[113];
  assign o[58199] = i[113];
  assign o[58200] = i[113];
  assign o[58201] = i[113];
  assign o[58202] = i[113];
  assign o[58203] = i[113];
  assign o[58204] = i[113];
  assign o[58205] = i[113];
  assign o[58206] = i[113];
  assign o[58207] = i[113];
  assign o[58208] = i[113];
  assign o[58209] = i[113];
  assign o[58210] = i[113];
  assign o[58211] = i[113];
  assign o[58212] = i[113];
  assign o[58213] = i[113];
  assign o[58214] = i[113];
  assign o[58215] = i[113];
  assign o[58216] = i[113];
  assign o[58217] = i[113];
  assign o[58218] = i[113];
  assign o[58219] = i[113];
  assign o[58220] = i[113];
  assign o[58221] = i[113];
  assign o[58222] = i[113];
  assign o[58223] = i[113];
  assign o[58224] = i[113];
  assign o[58225] = i[113];
  assign o[58226] = i[113];
  assign o[58227] = i[113];
  assign o[58228] = i[113];
  assign o[58229] = i[113];
  assign o[58230] = i[113];
  assign o[58231] = i[113];
  assign o[58232] = i[113];
  assign o[58233] = i[113];
  assign o[58234] = i[113];
  assign o[58235] = i[113];
  assign o[58236] = i[113];
  assign o[58237] = i[113];
  assign o[58238] = i[113];
  assign o[58239] = i[113];
  assign o[58240] = i[113];
  assign o[58241] = i[113];
  assign o[58242] = i[113];
  assign o[58243] = i[113];
  assign o[58244] = i[113];
  assign o[58245] = i[113];
  assign o[58246] = i[113];
  assign o[58247] = i[113];
  assign o[58248] = i[113];
  assign o[58249] = i[113];
  assign o[58250] = i[113];
  assign o[58251] = i[113];
  assign o[58252] = i[113];
  assign o[58253] = i[113];
  assign o[58254] = i[113];
  assign o[58255] = i[113];
  assign o[58256] = i[113];
  assign o[58257] = i[113];
  assign o[58258] = i[113];
  assign o[58259] = i[113];
  assign o[58260] = i[113];
  assign o[58261] = i[113];
  assign o[58262] = i[113];
  assign o[58263] = i[113];
  assign o[58264] = i[113];
  assign o[58265] = i[113];
  assign o[58266] = i[113];
  assign o[58267] = i[113];
  assign o[58268] = i[113];
  assign o[58269] = i[113];
  assign o[58270] = i[113];
  assign o[58271] = i[113];
  assign o[58272] = i[113];
  assign o[58273] = i[113];
  assign o[58274] = i[113];
  assign o[58275] = i[113];
  assign o[58276] = i[113];
  assign o[58277] = i[113];
  assign o[58278] = i[113];
  assign o[58279] = i[113];
  assign o[58280] = i[113];
  assign o[58281] = i[113];
  assign o[58282] = i[113];
  assign o[58283] = i[113];
  assign o[58284] = i[113];
  assign o[58285] = i[113];
  assign o[58286] = i[113];
  assign o[58287] = i[113];
  assign o[58288] = i[113];
  assign o[58289] = i[113];
  assign o[58290] = i[113];
  assign o[58291] = i[113];
  assign o[58292] = i[113];
  assign o[58293] = i[113];
  assign o[58294] = i[113];
  assign o[58295] = i[113];
  assign o[58296] = i[113];
  assign o[58297] = i[113];
  assign o[58298] = i[113];
  assign o[58299] = i[113];
  assign o[58300] = i[113];
  assign o[58301] = i[113];
  assign o[58302] = i[113];
  assign o[58303] = i[113];
  assign o[58304] = i[113];
  assign o[58305] = i[113];
  assign o[58306] = i[113];
  assign o[58307] = i[113];
  assign o[58308] = i[113];
  assign o[58309] = i[113];
  assign o[58310] = i[113];
  assign o[58311] = i[113];
  assign o[58312] = i[113];
  assign o[58313] = i[113];
  assign o[58314] = i[113];
  assign o[58315] = i[113];
  assign o[58316] = i[113];
  assign o[58317] = i[113];
  assign o[58318] = i[113];
  assign o[58319] = i[113];
  assign o[58320] = i[113];
  assign o[58321] = i[113];
  assign o[58322] = i[113];
  assign o[58323] = i[113];
  assign o[58324] = i[113];
  assign o[58325] = i[113];
  assign o[58326] = i[113];
  assign o[58327] = i[113];
  assign o[58328] = i[113];
  assign o[58329] = i[113];
  assign o[58330] = i[113];
  assign o[58331] = i[113];
  assign o[58332] = i[113];
  assign o[58333] = i[113];
  assign o[58334] = i[113];
  assign o[58335] = i[113];
  assign o[58336] = i[113];
  assign o[58337] = i[113];
  assign o[58338] = i[113];
  assign o[58339] = i[113];
  assign o[58340] = i[113];
  assign o[58341] = i[113];
  assign o[58342] = i[113];
  assign o[58343] = i[113];
  assign o[58344] = i[113];
  assign o[58345] = i[113];
  assign o[58346] = i[113];
  assign o[58347] = i[113];
  assign o[58348] = i[113];
  assign o[58349] = i[113];
  assign o[58350] = i[113];
  assign o[58351] = i[113];
  assign o[58352] = i[113];
  assign o[58353] = i[113];
  assign o[58354] = i[113];
  assign o[58355] = i[113];
  assign o[58356] = i[113];
  assign o[58357] = i[113];
  assign o[58358] = i[113];
  assign o[58359] = i[113];
  assign o[58360] = i[113];
  assign o[58361] = i[113];
  assign o[58362] = i[113];
  assign o[58363] = i[113];
  assign o[58364] = i[113];
  assign o[58365] = i[113];
  assign o[58366] = i[113];
  assign o[58367] = i[113];
  assign o[57344] = i[112];
  assign o[57345] = i[112];
  assign o[57346] = i[112];
  assign o[57347] = i[112];
  assign o[57348] = i[112];
  assign o[57349] = i[112];
  assign o[57350] = i[112];
  assign o[57351] = i[112];
  assign o[57352] = i[112];
  assign o[57353] = i[112];
  assign o[57354] = i[112];
  assign o[57355] = i[112];
  assign o[57356] = i[112];
  assign o[57357] = i[112];
  assign o[57358] = i[112];
  assign o[57359] = i[112];
  assign o[57360] = i[112];
  assign o[57361] = i[112];
  assign o[57362] = i[112];
  assign o[57363] = i[112];
  assign o[57364] = i[112];
  assign o[57365] = i[112];
  assign o[57366] = i[112];
  assign o[57367] = i[112];
  assign o[57368] = i[112];
  assign o[57369] = i[112];
  assign o[57370] = i[112];
  assign o[57371] = i[112];
  assign o[57372] = i[112];
  assign o[57373] = i[112];
  assign o[57374] = i[112];
  assign o[57375] = i[112];
  assign o[57376] = i[112];
  assign o[57377] = i[112];
  assign o[57378] = i[112];
  assign o[57379] = i[112];
  assign o[57380] = i[112];
  assign o[57381] = i[112];
  assign o[57382] = i[112];
  assign o[57383] = i[112];
  assign o[57384] = i[112];
  assign o[57385] = i[112];
  assign o[57386] = i[112];
  assign o[57387] = i[112];
  assign o[57388] = i[112];
  assign o[57389] = i[112];
  assign o[57390] = i[112];
  assign o[57391] = i[112];
  assign o[57392] = i[112];
  assign o[57393] = i[112];
  assign o[57394] = i[112];
  assign o[57395] = i[112];
  assign o[57396] = i[112];
  assign o[57397] = i[112];
  assign o[57398] = i[112];
  assign o[57399] = i[112];
  assign o[57400] = i[112];
  assign o[57401] = i[112];
  assign o[57402] = i[112];
  assign o[57403] = i[112];
  assign o[57404] = i[112];
  assign o[57405] = i[112];
  assign o[57406] = i[112];
  assign o[57407] = i[112];
  assign o[57408] = i[112];
  assign o[57409] = i[112];
  assign o[57410] = i[112];
  assign o[57411] = i[112];
  assign o[57412] = i[112];
  assign o[57413] = i[112];
  assign o[57414] = i[112];
  assign o[57415] = i[112];
  assign o[57416] = i[112];
  assign o[57417] = i[112];
  assign o[57418] = i[112];
  assign o[57419] = i[112];
  assign o[57420] = i[112];
  assign o[57421] = i[112];
  assign o[57422] = i[112];
  assign o[57423] = i[112];
  assign o[57424] = i[112];
  assign o[57425] = i[112];
  assign o[57426] = i[112];
  assign o[57427] = i[112];
  assign o[57428] = i[112];
  assign o[57429] = i[112];
  assign o[57430] = i[112];
  assign o[57431] = i[112];
  assign o[57432] = i[112];
  assign o[57433] = i[112];
  assign o[57434] = i[112];
  assign o[57435] = i[112];
  assign o[57436] = i[112];
  assign o[57437] = i[112];
  assign o[57438] = i[112];
  assign o[57439] = i[112];
  assign o[57440] = i[112];
  assign o[57441] = i[112];
  assign o[57442] = i[112];
  assign o[57443] = i[112];
  assign o[57444] = i[112];
  assign o[57445] = i[112];
  assign o[57446] = i[112];
  assign o[57447] = i[112];
  assign o[57448] = i[112];
  assign o[57449] = i[112];
  assign o[57450] = i[112];
  assign o[57451] = i[112];
  assign o[57452] = i[112];
  assign o[57453] = i[112];
  assign o[57454] = i[112];
  assign o[57455] = i[112];
  assign o[57456] = i[112];
  assign o[57457] = i[112];
  assign o[57458] = i[112];
  assign o[57459] = i[112];
  assign o[57460] = i[112];
  assign o[57461] = i[112];
  assign o[57462] = i[112];
  assign o[57463] = i[112];
  assign o[57464] = i[112];
  assign o[57465] = i[112];
  assign o[57466] = i[112];
  assign o[57467] = i[112];
  assign o[57468] = i[112];
  assign o[57469] = i[112];
  assign o[57470] = i[112];
  assign o[57471] = i[112];
  assign o[57472] = i[112];
  assign o[57473] = i[112];
  assign o[57474] = i[112];
  assign o[57475] = i[112];
  assign o[57476] = i[112];
  assign o[57477] = i[112];
  assign o[57478] = i[112];
  assign o[57479] = i[112];
  assign o[57480] = i[112];
  assign o[57481] = i[112];
  assign o[57482] = i[112];
  assign o[57483] = i[112];
  assign o[57484] = i[112];
  assign o[57485] = i[112];
  assign o[57486] = i[112];
  assign o[57487] = i[112];
  assign o[57488] = i[112];
  assign o[57489] = i[112];
  assign o[57490] = i[112];
  assign o[57491] = i[112];
  assign o[57492] = i[112];
  assign o[57493] = i[112];
  assign o[57494] = i[112];
  assign o[57495] = i[112];
  assign o[57496] = i[112];
  assign o[57497] = i[112];
  assign o[57498] = i[112];
  assign o[57499] = i[112];
  assign o[57500] = i[112];
  assign o[57501] = i[112];
  assign o[57502] = i[112];
  assign o[57503] = i[112];
  assign o[57504] = i[112];
  assign o[57505] = i[112];
  assign o[57506] = i[112];
  assign o[57507] = i[112];
  assign o[57508] = i[112];
  assign o[57509] = i[112];
  assign o[57510] = i[112];
  assign o[57511] = i[112];
  assign o[57512] = i[112];
  assign o[57513] = i[112];
  assign o[57514] = i[112];
  assign o[57515] = i[112];
  assign o[57516] = i[112];
  assign o[57517] = i[112];
  assign o[57518] = i[112];
  assign o[57519] = i[112];
  assign o[57520] = i[112];
  assign o[57521] = i[112];
  assign o[57522] = i[112];
  assign o[57523] = i[112];
  assign o[57524] = i[112];
  assign o[57525] = i[112];
  assign o[57526] = i[112];
  assign o[57527] = i[112];
  assign o[57528] = i[112];
  assign o[57529] = i[112];
  assign o[57530] = i[112];
  assign o[57531] = i[112];
  assign o[57532] = i[112];
  assign o[57533] = i[112];
  assign o[57534] = i[112];
  assign o[57535] = i[112];
  assign o[57536] = i[112];
  assign o[57537] = i[112];
  assign o[57538] = i[112];
  assign o[57539] = i[112];
  assign o[57540] = i[112];
  assign o[57541] = i[112];
  assign o[57542] = i[112];
  assign o[57543] = i[112];
  assign o[57544] = i[112];
  assign o[57545] = i[112];
  assign o[57546] = i[112];
  assign o[57547] = i[112];
  assign o[57548] = i[112];
  assign o[57549] = i[112];
  assign o[57550] = i[112];
  assign o[57551] = i[112];
  assign o[57552] = i[112];
  assign o[57553] = i[112];
  assign o[57554] = i[112];
  assign o[57555] = i[112];
  assign o[57556] = i[112];
  assign o[57557] = i[112];
  assign o[57558] = i[112];
  assign o[57559] = i[112];
  assign o[57560] = i[112];
  assign o[57561] = i[112];
  assign o[57562] = i[112];
  assign o[57563] = i[112];
  assign o[57564] = i[112];
  assign o[57565] = i[112];
  assign o[57566] = i[112];
  assign o[57567] = i[112];
  assign o[57568] = i[112];
  assign o[57569] = i[112];
  assign o[57570] = i[112];
  assign o[57571] = i[112];
  assign o[57572] = i[112];
  assign o[57573] = i[112];
  assign o[57574] = i[112];
  assign o[57575] = i[112];
  assign o[57576] = i[112];
  assign o[57577] = i[112];
  assign o[57578] = i[112];
  assign o[57579] = i[112];
  assign o[57580] = i[112];
  assign o[57581] = i[112];
  assign o[57582] = i[112];
  assign o[57583] = i[112];
  assign o[57584] = i[112];
  assign o[57585] = i[112];
  assign o[57586] = i[112];
  assign o[57587] = i[112];
  assign o[57588] = i[112];
  assign o[57589] = i[112];
  assign o[57590] = i[112];
  assign o[57591] = i[112];
  assign o[57592] = i[112];
  assign o[57593] = i[112];
  assign o[57594] = i[112];
  assign o[57595] = i[112];
  assign o[57596] = i[112];
  assign o[57597] = i[112];
  assign o[57598] = i[112];
  assign o[57599] = i[112];
  assign o[57600] = i[112];
  assign o[57601] = i[112];
  assign o[57602] = i[112];
  assign o[57603] = i[112];
  assign o[57604] = i[112];
  assign o[57605] = i[112];
  assign o[57606] = i[112];
  assign o[57607] = i[112];
  assign o[57608] = i[112];
  assign o[57609] = i[112];
  assign o[57610] = i[112];
  assign o[57611] = i[112];
  assign o[57612] = i[112];
  assign o[57613] = i[112];
  assign o[57614] = i[112];
  assign o[57615] = i[112];
  assign o[57616] = i[112];
  assign o[57617] = i[112];
  assign o[57618] = i[112];
  assign o[57619] = i[112];
  assign o[57620] = i[112];
  assign o[57621] = i[112];
  assign o[57622] = i[112];
  assign o[57623] = i[112];
  assign o[57624] = i[112];
  assign o[57625] = i[112];
  assign o[57626] = i[112];
  assign o[57627] = i[112];
  assign o[57628] = i[112];
  assign o[57629] = i[112];
  assign o[57630] = i[112];
  assign o[57631] = i[112];
  assign o[57632] = i[112];
  assign o[57633] = i[112];
  assign o[57634] = i[112];
  assign o[57635] = i[112];
  assign o[57636] = i[112];
  assign o[57637] = i[112];
  assign o[57638] = i[112];
  assign o[57639] = i[112];
  assign o[57640] = i[112];
  assign o[57641] = i[112];
  assign o[57642] = i[112];
  assign o[57643] = i[112];
  assign o[57644] = i[112];
  assign o[57645] = i[112];
  assign o[57646] = i[112];
  assign o[57647] = i[112];
  assign o[57648] = i[112];
  assign o[57649] = i[112];
  assign o[57650] = i[112];
  assign o[57651] = i[112];
  assign o[57652] = i[112];
  assign o[57653] = i[112];
  assign o[57654] = i[112];
  assign o[57655] = i[112];
  assign o[57656] = i[112];
  assign o[57657] = i[112];
  assign o[57658] = i[112];
  assign o[57659] = i[112];
  assign o[57660] = i[112];
  assign o[57661] = i[112];
  assign o[57662] = i[112];
  assign o[57663] = i[112];
  assign o[57664] = i[112];
  assign o[57665] = i[112];
  assign o[57666] = i[112];
  assign o[57667] = i[112];
  assign o[57668] = i[112];
  assign o[57669] = i[112];
  assign o[57670] = i[112];
  assign o[57671] = i[112];
  assign o[57672] = i[112];
  assign o[57673] = i[112];
  assign o[57674] = i[112];
  assign o[57675] = i[112];
  assign o[57676] = i[112];
  assign o[57677] = i[112];
  assign o[57678] = i[112];
  assign o[57679] = i[112];
  assign o[57680] = i[112];
  assign o[57681] = i[112];
  assign o[57682] = i[112];
  assign o[57683] = i[112];
  assign o[57684] = i[112];
  assign o[57685] = i[112];
  assign o[57686] = i[112];
  assign o[57687] = i[112];
  assign o[57688] = i[112];
  assign o[57689] = i[112];
  assign o[57690] = i[112];
  assign o[57691] = i[112];
  assign o[57692] = i[112];
  assign o[57693] = i[112];
  assign o[57694] = i[112];
  assign o[57695] = i[112];
  assign o[57696] = i[112];
  assign o[57697] = i[112];
  assign o[57698] = i[112];
  assign o[57699] = i[112];
  assign o[57700] = i[112];
  assign o[57701] = i[112];
  assign o[57702] = i[112];
  assign o[57703] = i[112];
  assign o[57704] = i[112];
  assign o[57705] = i[112];
  assign o[57706] = i[112];
  assign o[57707] = i[112];
  assign o[57708] = i[112];
  assign o[57709] = i[112];
  assign o[57710] = i[112];
  assign o[57711] = i[112];
  assign o[57712] = i[112];
  assign o[57713] = i[112];
  assign o[57714] = i[112];
  assign o[57715] = i[112];
  assign o[57716] = i[112];
  assign o[57717] = i[112];
  assign o[57718] = i[112];
  assign o[57719] = i[112];
  assign o[57720] = i[112];
  assign o[57721] = i[112];
  assign o[57722] = i[112];
  assign o[57723] = i[112];
  assign o[57724] = i[112];
  assign o[57725] = i[112];
  assign o[57726] = i[112];
  assign o[57727] = i[112];
  assign o[57728] = i[112];
  assign o[57729] = i[112];
  assign o[57730] = i[112];
  assign o[57731] = i[112];
  assign o[57732] = i[112];
  assign o[57733] = i[112];
  assign o[57734] = i[112];
  assign o[57735] = i[112];
  assign o[57736] = i[112];
  assign o[57737] = i[112];
  assign o[57738] = i[112];
  assign o[57739] = i[112];
  assign o[57740] = i[112];
  assign o[57741] = i[112];
  assign o[57742] = i[112];
  assign o[57743] = i[112];
  assign o[57744] = i[112];
  assign o[57745] = i[112];
  assign o[57746] = i[112];
  assign o[57747] = i[112];
  assign o[57748] = i[112];
  assign o[57749] = i[112];
  assign o[57750] = i[112];
  assign o[57751] = i[112];
  assign o[57752] = i[112];
  assign o[57753] = i[112];
  assign o[57754] = i[112];
  assign o[57755] = i[112];
  assign o[57756] = i[112];
  assign o[57757] = i[112];
  assign o[57758] = i[112];
  assign o[57759] = i[112];
  assign o[57760] = i[112];
  assign o[57761] = i[112];
  assign o[57762] = i[112];
  assign o[57763] = i[112];
  assign o[57764] = i[112];
  assign o[57765] = i[112];
  assign o[57766] = i[112];
  assign o[57767] = i[112];
  assign o[57768] = i[112];
  assign o[57769] = i[112];
  assign o[57770] = i[112];
  assign o[57771] = i[112];
  assign o[57772] = i[112];
  assign o[57773] = i[112];
  assign o[57774] = i[112];
  assign o[57775] = i[112];
  assign o[57776] = i[112];
  assign o[57777] = i[112];
  assign o[57778] = i[112];
  assign o[57779] = i[112];
  assign o[57780] = i[112];
  assign o[57781] = i[112];
  assign o[57782] = i[112];
  assign o[57783] = i[112];
  assign o[57784] = i[112];
  assign o[57785] = i[112];
  assign o[57786] = i[112];
  assign o[57787] = i[112];
  assign o[57788] = i[112];
  assign o[57789] = i[112];
  assign o[57790] = i[112];
  assign o[57791] = i[112];
  assign o[57792] = i[112];
  assign o[57793] = i[112];
  assign o[57794] = i[112];
  assign o[57795] = i[112];
  assign o[57796] = i[112];
  assign o[57797] = i[112];
  assign o[57798] = i[112];
  assign o[57799] = i[112];
  assign o[57800] = i[112];
  assign o[57801] = i[112];
  assign o[57802] = i[112];
  assign o[57803] = i[112];
  assign o[57804] = i[112];
  assign o[57805] = i[112];
  assign o[57806] = i[112];
  assign o[57807] = i[112];
  assign o[57808] = i[112];
  assign o[57809] = i[112];
  assign o[57810] = i[112];
  assign o[57811] = i[112];
  assign o[57812] = i[112];
  assign o[57813] = i[112];
  assign o[57814] = i[112];
  assign o[57815] = i[112];
  assign o[57816] = i[112];
  assign o[57817] = i[112];
  assign o[57818] = i[112];
  assign o[57819] = i[112];
  assign o[57820] = i[112];
  assign o[57821] = i[112];
  assign o[57822] = i[112];
  assign o[57823] = i[112];
  assign o[57824] = i[112];
  assign o[57825] = i[112];
  assign o[57826] = i[112];
  assign o[57827] = i[112];
  assign o[57828] = i[112];
  assign o[57829] = i[112];
  assign o[57830] = i[112];
  assign o[57831] = i[112];
  assign o[57832] = i[112];
  assign o[57833] = i[112];
  assign o[57834] = i[112];
  assign o[57835] = i[112];
  assign o[57836] = i[112];
  assign o[57837] = i[112];
  assign o[57838] = i[112];
  assign o[57839] = i[112];
  assign o[57840] = i[112];
  assign o[57841] = i[112];
  assign o[57842] = i[112];
  assign o[57843] = i[112];
  assign o[57844] = i[112];
  assign o[57845] = i[112];
  assign o[57846] = i[112];
  assign o[57847] = i[112];
  assign o[57848] = i[112];
  assign o[57849] = i[112];
  assign o[57850] = i[112];
  assign o[57851] = i[112];
  assign o[57852] = i[112];
  assign o[57853] = i[112];
  assign o[57854] = i[112];
  assign o[57855] = i[112];
  assign o[56832] = i[111];
  assign o[56833] = i[111];
  assign o[56834] = i[111];
  assign o[56835] = i[111];
  assign o[56836] = i[111];
  assign o[56837] = i[111];
  assign o[56838] = i[111];
  assign o[56839] = i[111];
  assign o[56840] = i[111];
  assign o[56841] = i[111];
  assign o[56842] = i[111];
  assign o[56843] = i[111];
  assign o[56844] = i[111];
  assign o[56845] = i[111];
  assign o[56846] = i[111];
  assign o[56847] = i[111];
  assign o[56848] = i[111];
  assign o[56849] = i[111];
  assign o[56850] = i[111];
  assign o[56851] = i[111];
  assign o[56852] = i[111];
  assign o[56853] = i[111];
  assign o[56854] = i[111];
  assign o[56855] = i[111];
  assign o[56856] = i[111];
  assign o[56857] = i[111];
  assign o[56858] = i[111];
  assign o[56859] = i[111];
  assign o[56860] = i[111];
  assign o[56861] = i[111];
  assign o[56862] = i[111];
  assign o[56863] = i[111];
  assign o[56864] = i[111];
  assign o[56865] = i[111];
  assign o[56866] = i[111];
  assign o[56867] = i[111];
  assign o[56868] = i[111];
  assign o[56869] = i[111];
  assign o[56870] = i[111];
  assign o[56871] = i[111];
  assign o[56872] = i[111];
  assign o[56873] = i[111];
  assign o[56874] = i[111];
  assign o[56875] = i[111];
  assign o[56876] = i[111];
  assign o[56877] = i[111];
  assign o[56878] = i[111];
  assign o[56879] = i[111];
  assign o[56880] = i[111];
  assign o[56881] = i[111];
  assign o[56882] = i[111];
  assign o[56883] = i[111];
  assign o[56884] = i[111];
  assign o[56885] = i[111];
  assign o[56886] = i[111];
  assign o[56887] = i[111];
  assign o[56888] = i[111];
  assign o[56889] = i[111];
  assign o[56890] = i[111];
  assign o[56891] = i[111];
  assign o[56892] = i[111];
  assign o[56893] = i[111];
  assign o[56894] = i[111];
  assign o[56895] = i[111];
  assign o[56896] = i[111];
  assign o[56897] = i[111];
  assign o[56898] = i[111];
  assign o[56899] = i[111];
  assign o[56900] = i[111];
  assign o[56901] = i[111];
  assign o[56902] = i[111];
  assign o[56903] = i[111];
  assign o[56904] = i[111];
  assign o[56905] = i[111];
  assign o[56906] = i[111];
  assign o[56907] = i[111];
  assign o[56908] = i[111];
  assign o[56909] = i[111];
  assign o[56910] = i[111];
  assign o[56911] = i[111];
  assign o[56912] = i[111];
  assign o[56913] = i[111];
  assign o[56914] = i[111];
  assign o[56915] = i[111];
  assign o[56916] = i[111];
  assign o[56917] = i[111];
  assign o[56918] = i[111];
  assign o[56919] = i[111];
  assign o[56920] = i[111];
  assign o[56921] = i[111];
  assign o[56922] = i[111];
  assign o[56923] = i[111];
  assign o[56924] = i[111];
  assign o[56925] = i[111];
  assign o[56926] = i[111];
  assign o[56927] = i[111];
  assign o[56928] = i[111];
  assign o[56929] = i[111];
  assign o[56930] = i[111];
  assign o[56931] = i[111];
  assign o[56932] = i[111];
  assign o[56933] = i[111];
  assign o[56934] = i[111];
  assign o[56935] = i[111];
  assign o[56936] = i[111];
  assign o[56937] = i[111];
  assign o[56938] = i[111];
  assign o[56939] = i[111];
  assign o[56940] = i[111];
  assign o[56941] = i[111];
  assign o[56942] = i[111];
  assign o[56943] = i[111];
  assign o[56944] = i[111];
  assign o[56945] = i[111];
  assign o[56946] = i[111];
  assign o[56947] = i[111];
  assign o[56948] = i[111];
  assign o[56949] = i[111];
  assign o[56950] = i[111];
  assign o[56951] = i[111];
  assign o[56952] = i[111];
  assign o[56953] = i[111];
  assign o[56954] = i[111];
  assign o[56955] = i[111];
  assign o[56956] = i[111];
  assign o[56957] = i[111];
  assign o[56958] = i[111];
  assign o[56959] = i[111];
  assign o[56960] = i[111];
  assign o[56961] = i[111];
  assign o[56962] = i[111];
  assign o[56963] = i[111];
  assign o[56964] = i[111];
  assign o[56965] = i[111];
  assign o[56966] = i[111];
  assign o[56967] = i[111];
  assign o[56968] = i[111];
  assign o[56969] = i[111];
  assign o[56970] = i[111];
  assign o[56971] = i[111];
  assign o[56972] = i[111];
  assign o[56973] = i[111];
  assign o[56974] = i[111];
  assign o[56975] = i[111];
  assign o[56976] = i[111];
  assign o[56977] = i[111];
  assign o[56978] = i[111];
  assign o[56979] = i[111];
  assign o[56980] = i[111];
  assign o[56981] = i[111];
  assign o[56982] = i[111];
  assign o[56983] = i[111];
  assign o[56984] = i[111];
  assign o[56985] = i[111];
  assign o[56986] = i[111];
  assign o[56987] = i[111];
  assign o[56988] = i[111];
  assign o[56989] = i[111];
  assign o[56990] = i[111];
  assign o[56991] = i[111];
  assign o[56992] = i[111];
  assign o[56993] = i[111];
  assign o[56994] = i[111];
  assign o[56995] = i[111];
  assign o[56996] = i[111];
  assign o[56997] = i[111];
  assign o[56998] = i[111];
  assign o[56999] = i[111];
  assign o[57000] = i[111];
  assign o[57001] = i[111];
  assign o[57002] = i[111];
  assign o[57003] = i[111];
  assign o[57004] = i[111];
  assign o[57005] = i[111];
  assign o[57006] = i[111];
  assign o[57007] = i[111];
  assign o[57008] = i[111];
  assign o[57009] = i[111];
  assign o[57010] = i[111];
  assign o[57011] = i[111];
  assign o[57012] = i[111];
  assign o[57013] = i[111];
  assign o[57014] = i[111];
  assign o[57015] = i[111];
  assign o[57016] = i[111];
  assign o[57017] = i[111];
  assign o[57018] = i[111];
  assign o[57019] = i[111];
  assign o[57020] = i[111];
  assign o[57021] = i[111];
  assign o[57022] = i[111];
  assign o[57023] = i[111];
  assign o[57024] = i[111];
  assign o[57025] = i[111];
  assign o[57026] = i[111];
  assign o[57027] = i[111];
  assign o[57028] = i[111];
  assign o[57029] = i[111];
  assign o[57030] = i[111];
  assign o[57031] = i[111];
  assign o[57032] = i[111];
  assign o[57033] = i[111];
  assign o[57034] = i[111];
  assign o[57035] = i[111];
  assign o[57036] = i[111];
  assign o[57037] = i[111];
  assign o[57038] = i[111];
  assign o[57039] = i[111];
  assign o[57040] = i[111];
  assign o[57041] = i[111];
  assign o[57042] = i[111];
  assign o[57043] = i[111];
  assign o[57044] = i[111];
  assign o[57045] = i[111];
  assign o[57046] = i[111];
  assign o[57047] = i[111];
  assign o[57048] = i[111];
  assign o[57049] = i[111];
  assign o[57050] = i[111];
  assign o[57051] = i[111];
  assign o[57052] = i[111];
  assign o[57053] = i[111];
  assign o[57054] = i[111];
  assign o[57055] = i[111];
  assign o[57056] = i[111];
  assign o[57057] = i[111];
  assign o[57058] = i[111];
  assign o[57059] = i[111];
  assign o[57060] = i[111];
  assign o[57061] = i[111];
  assign o[57062] = i[111];
  assign o[57063] = i[111];
  assign o[57064] = i[111];
  assign o[57065] = i[111];
  assign o[57066] = i[111];
  assign o[57067] = i[111];
  assign o[57068] = i[111];
  assign o[57069] = i[111];
  assign o[57070] = i[111];
  assign o[57071] = i[111];
  assign o[57072] = i[111];
  assign o[57073] = i[111];
  assign o[57074] = i[111];
  assign o[57075] = i[111];
  assign o[57076] = i[111];
  assign o[57077] = i[111];
  assign o[57078] = i[111];
  assign o[57079] = i[111];
  assign o[57080] = i[111];
  assign o[57081] = i[111];
  assign o[57082] = i[111];
  assign o[57083] = i[111];
  assign o[57084] = i[111];
  assign o[57085] = i[111];
  assign o[57086] = i[111];
  assign o[57087] = i[111];
  assign o[57088] = i[111];
  assign o[57089] = i[111];
  assign o[57090] = i[111];
  assign o[57091] = i[111];
  assign o[57092] = i[111];
  assign o[57093] = i[111];
  assign o[57094] = i[111];
  assign o[57095] = i[111];
  assign o[57096] = i[111];
  assign o[57097] = i[111];
  assign o[57098] = i[111];
  assign o[57099] = i[111];
  assign o[57100] = i[111];
  assign o[57101] = i[111];
  assign o[57102] = i[111];
  assign o[57103] = i[111];
  assign o[57104] = i[111];
  assign o[57105] = i[111];
  assign o[57106] = i[111];
  assign o[57107] = i[111];
  assign o[57108] = i[111];
  assign o[57109] = i[111];
  assign o[57110] = i[111];
  assign o[57111] = i[111];
  assign o[57112] = i[111];
  assign o[57113] = i[111];
  assign o[57114] = i[111];
  assign o[57115] = i[111];
  assign o[57116] = i[111];
  assign o[57117] = i[111];
  assign o[57118] = i[111];
  assign o[57119] = i[111];
  assign o[57120] = i[111];
  assign o[57121] = i[111];
  assign o[57122] = i[111];
  assign o[57123] = i[111];
  assign o[57124] = i[111];
  assign o[57125] = i[111];
  assign o[57126] = i[111];
  assign o[57127] = i[111];
  assign o[57128] = i[111];
  assign o[57129] = i[111];
  assign o[57130] = i[111];
  assign o[57131] = i[111];
  assign o[57132] = i[111];
  assign o[57133] = i[111];
  assign o[57134] = i[111];
  assign o[57135] = i[111];
  assign o[57136] = i[111];
  assign o[57137] = i[111];
  assign o[57138] = i[111];
  assign o[57139] = i[111];
  assign o[57140] = i[111];
  assign o[57141] = i[111];
  assign o[57142] = i[111];
  assign o[57143] = i[111];
  assign o[57144] = i[111];
  assign o[57145] = i[111];
  assign o[57146] = i[111];
  assign o[57147] = i[111];
  assign o[57148] = i[111];
  assign o[57149] = i[111];
  assign o[57150] = i[111];
  assign o[57151] = i[111];
  assign o[57152] = i[111];
  assign o[57153] = i[111];
  assign o[57154] = i[111];
  assign o[57155] = i[111];
  assign o[57156] = i[111];
  assign o[57157] = i[111];
  assign o[57158] = i[111];
  assign o[57159] = i[111];
  assign o[57160] = i[111];
  assign o[57161] = i[111];
  assign o[57162] = i[111];
  assign o[57163] = i[111];
  assign o[57164] = i[111];
  assign o[57165] = i[111];
  assign o[57166] = i[111];
  assign o[57167] = i[111];
  assign o[57168] = i[111];
  assign o[57169] = i[111];
  assign o[57170] = i[111];
  assign o[57171] = i[111];
  assign o[57172] = i[111];
  assign o[57173] = i[111];
  assign o[57174] = i[111];
  assign o[57175] = i[111];
  assign o[57176] = i[111];
  assign o[57177] = i[111];
  assign o[57178] = i[111];
  assign o[57179] = i[111];
  assign o[57180] = i[111];
  assign o[57181] = i[111];
  assign o[57182] = i[111];
  assign o[57183] = i[111];
  assign o[57184] = i[111];
  assign o[57185] = i[111];
  assign o[57186] = i[111];
  assign o[57187] = i[111];
  assign o[57188] = i[111];
  assign o[57189] = i[111];
  assign o[57190] = i[111];
  assign o[57191] = i[111];
  assign o[57192] = i[111];
  assign o[57193] = i[111];
  assign o[57194] = i[111];
  assign o[57195] = i[111];
  assign o[57196] = i[111];
  assign o[57197] = i[111];
  assign o[57198] = i[111];
  assign o[57199] = i[111];
  assign o[57200] = i[111];
  assign o[57201] = i[111];
  assign o[57202] = i[111];
  assign o[57203] = i[111];
  assign o[57204] = i[111];
  assign o[57205] = i[111];
  assign o[57206] = i[111];
  assign o[57207] = i[111];
  assign o[57208] = i[111];
  assign o[57209] = i[111];
  assign o[57210] = i[111];
  assign o[57211] = i[111];
  assign o[57212] = i[111];
  assign o[57213] = i[111];
  assign o[57214] = i[111];
  assign o[57215] = i[111];
  assign o[57216] = i[111];
  assign o[57217] = i[111];
  assign o[57218] = i[111];
  assign o[57219] = i[111];
  assign o[57220] = i[111];
  assign o[57221] = i[111];
  assign o[57222] = i[111];
  assign o[57223] = i[111];
  assign o[57224] = i[111];
  assign o[57225] = i[111];
  assign o[57226] = i[111];
  assign o[57227] = i[111];
  assign o[57228] = i[111];
  assign o[57229] = i[111];
  assign o[57230] = i[111];
  assign o[57231] = i[111];
  assign o[57232] = i[111];
  assign o[57233] = i[111];
  assign o[57234] = i[111];
  assign o[57235] = i[111];
  assign o[57236] = i[111];
  assign o[57237] = i[111];
  assign o[57238] = i[111];
  assign o[57239] = i[111];
  assign o[57240] = i[111];
  assign o[57241] = i[111];
  assign o[57242] = i[111];
  assign o[57243] = i[111];
  assign o[57244] = i[111];
  assign o[57245] = i[111];
  assign o[57246] = i[111];
  assign o[57247] = i[111];
  assign o[57248] = i[111];
  assign o[57249] = i[111];
  assign o[57250] = i[111];
  assign o[57251] = i[111];
  assign o[57252] = i[111];
  assign o[57253] = i[111];
  assign o[57254] = i[111];
  assign o[57255] = i[111];
  assign o[57256] = i[111];
  assign o[57257] = i[111];
  assign o[57258] = i[111];
  assign o[57259] = i[111];
  assign o[57260] = i[111];
  assign o[57261] = i[111];
  assign o[57262] = i[111];
  assign o[57263] = i[111];
  assign o[57264] = i[111];
  assign o[57265] = i[111];
  assign o[57266] = i[111];
  assign o[57267] = i[111];
  assign o[57268] = i[111];
  assign o[57269] = i[111];
  assign o[57270] = i[111];
  assign o[57271] = i[111];
  assign o[57272] = i[111];
  assign o[57273] = i[111];
  assign o[57274] = i[111];
  assign o[57275] = i[111];
  assign o[57276] = i[111];
  assign o[57277] = i[111];
  assign o[57278] = i[111];
  assign o[57279] = i[111];
  assign o[57280] = i[111];
  assign o[57281] = i[111];
  assign o[57282] = i[111];
  assign o[57283] = i[111];
  assign o[57284] = i[111];
  assign o[57285] = i[111];
  assign o[57286] = i[111];
  assign o[57287] = i[111];
  assign o[57288] = i[111];
  assign o[57289] = i[111];
  assign o[57290] = i[111];
  assign o[57291] = i[111];
  assign o[57292] = i[111];
  assign o[57293] = i[111];
  assign o[57294] = i[111];
  assign o[57295] = i[111];
  assign o[57296] = i[111];
  assign o[57297] = i[111];
  assign o[57298] = i[111];
  assign o[57299] = i[111];
  assign o[57300] = i[111];
  assign o[57301] = i[111];
  assign o[57302] = i[111];
  assign o[57303] = i[111];
  assign o[57304] = i[111];
  assign o[57305] = i[111];
  assign o[57306] = i[111];
  assign o[57307] = i[111];
  assign o[57308] = i[111];
  assign o[57309] = i[111];
  assign o[57310] = i[111];
  assign o[57311] = i[111];
  assign o[57312] = i[111];
  assign o[57313] = i[111];
  assign o[57314] = i[111];
  assign o[57315] = i[111];
  assign o[57316] = i[111];
  assign o[57317] = i[111];
  assign o[57318] = i[111];
  assign o[57319] = i[111];
  assign o[57320] = i[111];
  assign o[57321] = i[111];
  assign o[57322] = i[111];
  assign o[57323] = i[111];
  assign o[57324] = i[111];
  assign o[57325] = i[111];
  assign o[57326] = i[111];
  assign o[57327] = i[111];
  assign o[57328] = i[111];
  assign o[57329] = i[111];
  assign o[57330] = i[111];
  assign o[57331] = i[111];
  assign o[57332] = i[111];
  assign o[57333] = i[111];
  assign o[57334] = i[111];
  assign o[57335] = i[111];
  assign o[57336] = i[111];
  assign o[57337] = i[111];
  assign o[57338] = i[111];
  assign o[57339] = i[111];
  assign o[57340] = i[111];
  assign o[57341] = i[111];
  assign o[57342] = i[111];
  assign o[57343] = i[111];
  assign o[56320] = i[110];
  assign o[56321] = i[110];
  assign o[56322] = i[110];
  assign o[56323] = i[110];
  assign o[56324] = i[110];
  assign o[56325] = i[110];
  assign o[56326] = i[110];
  assign o[56327] = i[110];
  assign o[56328] = i[110];
  assign o[56329] = i[110];
  assign o[56330] = i[110];
  assign o[56331] = i[110];
  assign o[56332] = i[110];
  assign o[56333] = i[110];
  assign o[56334] = i[110];
  assign o[56335] = i[110];
  assign o[56336] = i[110];
  assign o[56337] = i[110];
  assign o[56338] = i[110];
  assign o[56339] = i[110];
  assign o[56340] = i[110];
  assign o[56341] = i[110];
  assign o[56342] = i[110];
  assign o[56343] = i[110];
  assign o[56344] = i[110];
  assign o[56345] = i[110];
  assign o[56346] = i[110];
  assign o[56347] = i[110];
  assign o[56348] = i[110];
  assign o[56349] = i[110];
  assign o[56350] = i[110];
  assign o[56351] = i[110];
  assign o[56352] = i[110];
  assign o[56353] = i[110];
  assign o[56354] = i[110];
  assign o[56355] = i[110];
  assign o[56356] = i[110];
  assign o[56357] = i[110];
  assign o[56358] = i[110];
  assign o[56359] = i[110];
  assign o[56360] = i[110];
  assign o[56361] = i[110];
  assign o[56362] = i[110];
  assign o[56363] = i[110];
  assign o[56364] = i[110];
  assign o[56365] = i[110];
  assign o[56366] = i[110];
  assign o[56367] = i[110];
  assign o[56368] = i[110];
  assign o[56369] = i[110];
  assign o[56370] = i[110];
  assign o[56371] = i[110];
  assign o[56372] = i[110];
  assign o[56373] = i[110];
  assign o[56374] = i[110];
  assign o[56375] = i[110];
  assign o[56376] = i[110];
  assign o[56377] = i[110];
  assign o[56378] = i[110];
  assign o[56379] = i[110];
  assign o[56380] = i[110];
  assign o[56381] = i[110];
  assign o[56382] = i[110];
  assign o[56383] = i[110];
  assign o[56384] = i[110];
  assign o[56385] = i[110];
  assign o[56386] = i[110];
  assign o[56387] = i[110];
  assign o[56388] = i[110];
  assign o[56389] = i[110];
  assign o[56390] = i[110];
  assign o[56391] = i[110];
  assign o[56392] = i[110];
  assign o[56393] = i[110];
  assign o[56394] = i[110];
  assign o[56395] = i[110];
  assign o[56396] = i[110];
  assign o[56397] = i[110];
  assign o[56398] = i[110];
  assign o[56399] = i[110];
  assign o[56400] = i[110];
  assign o[56401] = i[110];
  assign o[56402] = i[110];
  assign o[56403] = i[110];
  assign o[56404] = i[110];
  assign o[56405] = i[110];
  assign o[56406] = i[110];
  assign o[56407] = i[110];
  assign o[56408] = i[110];
  assign o[56409] = i[110];
  assign o[56410] = i[110];
  assign o[56411] = i[110];
  assign o[56412] = i[110];
  assign o[56413] = i[110];
  assign o[56414] = i[110];
  assign o[56415] = i[110];
  assign o[56416] = i[110];
  assign o[56417] = i[110];
  assign o[56418] = i[110];
  assign o[56419] = i[110];
  assign o[56420] = i[110];
  assign o[56421] = i[110];
  assign o[56422] = i[110];
  assign o[56423] = i[110];
  assign o[56424] = i[110];
  assign o[56425] = i[110];
  assign o[56426] = i[110];
  assign o[56427] = i[110];
  assign o[56428] = i[110];
  assign o[56429] = i[110];
  assign o[56430] = i[110];
  assign o[56431] = i[110];
  assign o[56432] = i[110];
  assign o[56433] = i[110];
  assign o[56434] = i[110];
  assign o[56435] = i[110];
  assign o[56436] = i[110];
  assign o[56437] = i[110];
  assign o[56438] = i[110];
  assign o[56439] = i[110];
  assign o[56440] = i[110];
  assign o[56441] = i[110];
  assign o[56442] = i[110];
  assign o[56443] = i[110];
  assign o[56444] = i[110];
  assign o[56445] = i[110];
  assign o[56446] = i[110];
  assign o[56447] = i[110];
  assign o[56448] = i[110];
  assign o[56449] = i[110];
  assign o[56450] = i[110];
  assign o[56451] = i[110];
  assign o[56452] = i[110];
  assign o[56453] = i[110];
  assign o[56454] = i[110];
  assign o[56455] = i[110];
  assign o[56456] = i[110];
  assign o[56457] = i[110];
  assign o[56458] = i[110];
  assign o[56459] = i[110];
  assign o[56460] = i[110];
  assign o[56461] = i[110];
  assign o[56462] = i[110];
  assign o[56463] = i[110];
  assign o[56464] = i[110];
  assign o[56465] = i[110];
  assign o[56466] = i[110];
  assign o[56467] = i[110];
  assign o[56468] = i[110];
  assign o[56469] = i[110];
  assign o[56470] = i[110];
  assign o[56471] = i[110];
  assign o[56472] = i[110];
  assign o[56473] = i[110];
  assign o[56474] = i[110];
  assign o[56475] = i[110];
  assign o[56476] = i[110];
  assign o[56477] = i[110];
  assign o[56478] = i[110];
  assign o[56479] = i[110];
  assign o[56480] = i[110];
  assign o[56481] = i[110];
  assign o[56482] = i[110];
  assign o[56483] = i[110];
  assign o[56484] = i[110];
  assign o[56485] = i[110];
  assign o[56486] = i[110];
  assign o[56487] = i[110];
  assign o[56488] = i[110];
  assign o[56489] = i[110];
  assign o[56490] = i[110];
  assign o[56491] = i[110];
  assign o[56492] = i[110];
  assign o[56493] = i[110];
  assign o[56494] = i[110];
  assign o[56495] = i[110];
  assign o[56496] = i[110];
  assign o[56497] = i[110];
  assign o[56498] = i[110];
  assign o[56499] = i[110];
  assign o[56500] = i[110];
  assign o[56501] = i[110];
  assign o[56502] = i[110];
  assign o[56503] = i[110];
  assign o[56504] = i[110];
  assign o[56505] = i[110];
  assign o[56506] = i[110];
  assign o[56507] = i[110];
  assign o[56508] = i[110];
  assign o[56509] = i[110];
  assign o[56510] = i[110];
  assign o[56511] = i[110];
  assign o[56512] = i[110];
  assign o[56513] = i[110];
  assign o[56514] = i[110];
  assign o[56515] = i[110];
  assign o[56516] = i[110];
  assign o[56517] = i[110];
  assign o[56518] = i[110];
  assign o[56519] = i[110];
  assign o[56520] = i[110];
  assign o[56521] = i[110];
  assign o[56522] = i[110];
  assign o[56523] = i[110];
  assign o[56524] = i[110];
  assign o[56525] = i[110];
  assign o[56526] = i[110];
  assign o[56527] = i[110];
  assign o[56528] = i[110];
  assign o[56529] = i[110];
  assign o[56530] = i[110];
  assign o[56531] = i[110];
  assign o[56532] = i[110];
  assign o[56533] = i[110];
  assign o[56534] = i[110];
  assign o[56535] = i[110];
  assign o[56536] = i[110];
  assign o[56537] = i[110];
  assign o[56538] = i[110];
  assign o[56539] = i[110];
  assign o[56540] = i[110];
  assign o[56541] = i[110];
  assign o[56542] = i[110];
  assign o[56543] = i[110];
  assign o[56544] = i[110];
  assign o[56545] = i[110];
  assign o[56546] = i[110];
  assign o[56547] = i[110];
  assign o[56548] = i[110];
  assign o[56549] = i[110];
  assign o[56550] = i[110];
  assign o[56551] = i[110];
  assign o[56552] = i[110];
  assign o[56553] = i[110];
  assign o[56554] = i[110];
  assign o[56555] = i[110];
  assign o[56556] = i[110];
  assign o[56557] = i[110];
  assign o[56558] = i[110];
  assign o[56559] = i[110];
  assign o[56560] = i[110];
  assign o[56561] = i[110];
  assign o[56562] = i[110];
  assign o[56563] = i[110];
  assign o[56564] = i[110];
  assign o[56565] = i[110];
  assign o[56566] = i[110];
  assign o[56567] = i[110];
  assign o[56568] = i[110];
  assign o[56569] = i[110];
  assign o[56570] = i[110];
  assign o[56571] = i[110];
  assign o[56572] = i[110];
  assign o[56573] = i[110];
  assign o[56574] = i[110];
  assign o[56575] = i[110];
  assign o[56576] = i[110];
  assign o[56577] = i[110];
  assign o[56578] = i[110];
  assign o[56579] = i[110];
  assign o[56580] = i[110];
  assign o[56581] = i[110];
  assign o[56582] = i[110];
  assign o[56583] = i[110];
  assign o[56584] = i[110];
  assign o[56585] = i[110];
  assign o[56586] = i[110];
  assign o[56587] = i[110];
  assign o[56588] = i[110];
  assign o[56589] = i[110];
  assign o[56590] = i[110];
  assign o[56591] = i[110];
  assign o[56592] = i[110];
  assign o[56593] = i[110];
  assign o[56594] = i[110];
  assign o[56595] = i[110];
  assign o[56596] = i[110];
  assign o[56597] = i[110];
  assign o[56598] = i[110];
  assign o[56599] = i[110];
  assign o[56600] = i[110];
  assign o[56601] = i[110];
  assign o[56602] = i[110];
  assign o[56603] = i[110];
  assign o[56604] = i[110];
  assign o[56605] = i[110];
  assign o[56606] = i[110];
  assign o[56607] = i[110];
  assign o[56608] = i[110];
  assign o[56609] = i[110];
  assign o[56610] = i[110];
  assign o[56611] = i[110];
  assign o[56612] = i[110];
  assign o[56613] = i[110];
  assign o[56614] = i[110];
  assign o[56615] = i[110];
  assign o[56616] = i[110];
  assign o[56617] = i[110];
  assign o[56618] = i[110];
  assign o[56619] = i[110];
  assign o[56620] = i[110];
  assign o[56621] = i[110];
  assign o[56622] = i[110];
  assign o[56623] = i[110];
  assign o[56624] = i[110];
  assign o[56625] = i[110];
  assign o[56626] = i[110];
  assign o[56627] = i[110];
  assign o[56628] = i[110];
  assign o[56629] = i[110];
  assign o[56630] = i[110];
  assign o[56631] = i[110];
  assign o[56632] = i[110];
  assign o[56633] = i[110];
  assign o[56634] = i[110];
  assign o[56635] = i[110];
  assign o[56636] = i[110];
  assign o[56637] = i[110];
  assign o[56638] = i[110];
  assign o[56639] = i[110];
  assign o[56640] = i[110];
  assign o[56641] = i[110];
  assign o[56642] = i[110];
  assign o[56643] = i[110];
  assign o[56644] = i[110];
  assign o[56645] = i[110];
  assign o[56646] = i[110];
  assign o[56647] = i[110];
  assign o[56648] = i[110];
  assign o[56649] = i[110];
  assign o[56650] = i[110];
  assign o[56651] = i[110];
  assign o[56652] = i[110];
  assign o[56653] = i[110];
  assign o[56654] = i[110];
  assign o[56655] = i[110];
  assign o[56656] = i[110];
  assign o[56657] = i[110];
  assign o[56658] = i[110];
  assign o[56659] = i[110];
  assign o[56660] = i[110];
  assign o[56661] = i[110];
  assign o[56662] = i[110];
  assign o[56663] = i[110];
  assign o[56664] = i[110];
  assign o[56665] = i[110];
  assign o[56666] = i[110];
  assign o[56667] = i[110];
  assign o[56668] = i[110];
  assign o[56669] = i[110];
  assign o[56670] = i[110];
  assign o[56671] = i[110];
  assign o[56672] = i[110];
  assign o[56673] = i[110];
  assign o[56674] = i[110];
  assign o[56675] = i[110];
  assign o[56676] = i[110];
  assign o[56677] = i[110];
  assign o[56678] = i[110];
  assign o[56679] = i[110];
  assign o[56680] = i[110];
  assign o[56681] = i[110];
  assign o[56682] = i[110];
  assign o[56683] = i[110];
  assign o[56684] = i[110];
  assign o[56685] = i[110];
  assign o[56686] = i[110];
  assign o[56687] = i[110];
  assign o[56688] = i[110];
  assign o[56689] = i[110];
  assign o[56690] = i[110];
  assign o[56691] = i[110];
  assign o[56692] = i[110];
  assign o[56693] = i[110];
  assign o[56694] = i[110];
  assign o[56695] = i[110];
  assign o[56696] = i[110];
  assign o[56697] = i[110];
  assign o[56698] = i[110];
  assign o[56699] = i[110];
  assign o[56700] = i[110];
  assign o[56701] = i[110];
  assign o[56702] = i[110];
  assign o[56703] = i[110];
  assign o[56704] = i[110];
  assign o[56705] = i[110];
  assign o[56706] = i[110];
  assign o[56707] = i[110];
  assign o[56708] = i[110];
  assign o[56709] = i[110];
  assign o[56710] = i[110];
  assign o[56711] = i[110];
  assign o[56712] = i[110];
  assign o[56713] = i[110];
  assign o[56714] = i[110];
  assign o[56715] = i[110];
  assign o[56716] = i[110];
  assign o[56717] = i[110];
  assign o[56718] = i[110];
  assign o[56719] = i[110];
  assign o[56720] = i[110];
  assign o[56721] = i[110];
  assign o[56722] = i[110];
  assign o[56723] = i[110];
  assign o[56724] = i[110];
  assign o[56725] = i[110];
  assign o[56726] = i[110];
  assign o[56727] = i[110];
  assign o[56728] = i[110];
  assign o[56729] = i[110];
  assign o[56730] = i[110];
  assign o[56731] = i[110];
  assign o[56732] = i[110];
  assign o[56733] = i[110];
  assign o[56734] = i[110];
  assign o[56735] = i[110];
  assign o[56736] = i[110];
  assign o[56737] = i[110];
  assign o[56738] = i[110];
  assign o[56739] = i[110];
  assign o[56740] = i[110];
  assign o[56741] = i[110];
  assign o[56742] = i[110];
  assign o[56743] = i[110];
  assign o[56744] = i[110];
  assign o[56745] = i[110];
  assign o[56746] = i[110];
  assign o[56747] = i[110];
  assign o[56748] = i[110];
  assign o[56749] = i[110];
  assign o[56750] = i[110];
  assign o[56751] = i[110];
  assign o[56752] = i[110];
  assign o[56753] = i[110];
  assign o[56754] = i[110];
  assign o[56755] = i[110];
  assign o[56756] = i[110];
  assign o[56757] = i[110];
  assign o[56758] = i[110];
  assign o[56759] = i[110];
  assign o[56760] = i[110];
  assign o[56761] = i[110];
  assign o[56762] = i[110];
  assign o[56763] = i[110];
  assign o[56764] = i[110];
  assign o[56765] = i[110];
  assign o[56766] = i[110];
  assign o[56767] = i[110];
  assign o[56768] = i[110];
  assign o[56769] = i[110];
  assign o[56770] = i[110];
  assign o[56771] = i[110];
  assign o[56772] = i[110];
  assign o[56773] = i[110];
  assign o[56774] = i[110];
  assign o[56775] = i[110];
  assign o[56776] = i[110];
  assign o[56777] = i[110];
  assign o[56778] = i[110];
  assign o[56779] = i[110];
  assign o[56780] = i[110];
  assign o[56781] = i[110];
  assign o[56782] = i[110];
  assign o[56783] = i[110];
  assign o[56784] = i[110];
  assign o[56785] = i[110];
  assign o[56786] = i[110];
  assign o[56787] = i[110];
  assign o[56788] = i[110];
  assign o[56789] = i[110];
  assign o[56790] = i[110];
  assign o[56791] = i[110];
  assign o[56792] = i[110];
  assign o[56793] = i[110];
  assign o[56794] = i[110];
  assign o[56795] = i[110];
  assign o[56796] = i[110];
  assign o[56797] = i[110];
  assign o[56798] = i[110];
  assign o[56799] = i[110];
  assign o[56800] = i[110];
  assign o[56801] = i[110];
  assign o[56802] = i[110];
  assign o[56803] = i[110];
  assign o[56804] = i[110];
  assign o[56805] = i[110];
  assign o[56806] = i[110];
  assign o[56807] = i[110];
  assign o[56808] = i[110];
  assign o[56809] = i[110];
  assign o[56810] = i[110];
  assign o[56811] = i[110];
  assign o[56812] = i[110];
  assign o[56813] = i[110];
  assign o[56814] = i[110];
  assign o[56815] = i[110];
  assign o[56816] = i[110];
  assign o[56817] = i[110];
  assign o[56818] = i[110];
  assign o[56819] = i[110];
  assign o[56820] = i[110];
  assign o[56821] = i[110];
  assign o[56822] = i[110];
  assign o[56823] = i[110];
  assign o[56824] = i[110];
  assign o[56825] = i[110];
  assign o[56826] = i[110];
  assign o[56827] = i[110];
  assign o[56828] = i[110];
  assign o[56829] = i[110];
  assign o[56830] = i[110];
  assign o[56831] = i[110];
  assign o[55808] = i[109];
  assign o[55809] = i[109];
  assign o[55810] = i[109];
  assign o[55811] = i[109];
  assign o[55812] = i[109];
  assign o[55813] = i[109];
  assign o[55814] = i[109];
  assign o[55815] = i[109];
  assign o[55816] = i[109];
  assign o[55817] = i[109];
  assign o[55818] = i[109];
  assign o[55819] = i[109];
  assign o[55820] = i[109];
  assign o[55821] = i[109];
  assign o[55822] = i[109];
  assign o[55823] = i[109];
  assign o[55824] = i[109];
  assign o[55825] = i[109];
  assign o[55826] = i[109];
  assign o[55827] = i[109];
  assign o[55828] = i[109];
  assign o[55829] = i[109];
  assign o[55830] = i[109];
  assign o[55831] = i[109];
  assign o[55832] = i[109];
  assign o[55833] = i[109];
  assign o[55834] = i[109];
  assign o[55835] = i[109];
  assign o[55836] = i[109];
  assign o[55837] = i[109];
  assign o[55838] = i[109];
  assign o[55839] = i[109];
  assign o[55840] = i[109];
  assign o[55841] = i[109];
  assign o[55842] = i[109];
  assign o[55843] = i[109];
  assign o[55844] = i[109];
  assign o[55845] = i[109];
  assign o[55846] = i[109];
  assign o[55847] = i[109];
  assign o[55848] = i[109];
  assign o[55849] = i[109];
  assign o[55850] = i[109];
  assign o[55851] = i[109];
  assign o[55852] = i[109];
  assign o[55853] = i[109];
  assign o[55854] = i[109];
  assign o[55855] = i[109];
  assign o[55856] = i[109];
  assign o[55857] = i[109];
  assign o[55858] = i[109];
  assign o[55859] = i[109];
  assign o[55860] = i[109];
  assign o[55861] = i[109];
  assign o[55862] = i[109];
  assign o[55863] = i[109];
  assign o[55864] = i[109];
  assign o[55865] = i[109];
  assign o[55866] = i[109];
  assign o[55867] = i[109];
  assign o[55868] = i[109];
  assign o[55869] = i[109];
  assign o[55870] = i[109];
  assign o[55871] = i[109];
  assign o[55872] = i[109];
  assign o[55873] = i[109];
  assign o[55874] = i[109];
  assign o[55875] = i[109];
  assign o[55876] = i[109];
  assign o[55877] = i[109];
  assign o[55878] = i[109];
  assign o[55879] = i[109];
  assign o[55880] = i[109];
  assign o[55881] = i[109];
  assign o[55882] = i[109];
  assign o[55883] = i[109];
  assign o[55884] = i[109];
  assign o[55885] = i[109];
  assign o[55886] = i[109];
  assign o[55887] = i[109];
  assign o[55888] = i[109];
  assign o[55889] = i[109];
  assign o[55890] = i[109];
  assign o[55891] = i[109];
  assign o[55892] = i[109];
  assign o[55893] = i[109];
  assign o[55894] = i[109];
  assign o[55895] = i[109];
  assign o[55896] = i[109];
  assign o[55897] = i[109];
  assign o[55898] = i[109];
  assign o[55899] = i[109];
  assign o[55900] = i[109];
  assign o[55901] = i[109];
  assign o[55902] = i[109];
  assign o[55903] = i[109];
  assign o[55904] = i[109];
  assign o[55905] = i[109];
  assign o[55906] = i[109];
  assign o[55907] = i[109];
  assign o[55908] = i[109];
  assign o[55909] = i[109];
  assign o[55910] = i[109];
  assign o[55911] = i[109];
  assign o[55912] = i[109];
  assign o[55913] = i[109];
  assign o[55914] = i[109];
  assign o[55915] = i[109];
  assign o[55916] = i[109];
  assign o[55917] = i[109];
  assign o[55918] = i[109];
  assign o[55919] = i[109];
  assign o[55920] = i[109];
  assign o[55921] = i[109];
  assign o[55922] = i[109];
  assign o[55923] = i[109];
  assign o[55924] = i[109];
  assign o[55925] = i[109];
  assign o[55926] = i[109];
  assign o[55927] = i[109];
  assign o[55928] = i[109];
  assign o[55929] = i[109];
  assign o[55930] = i[109];
  assign o[55931] = i[109];
  assign o[55932] = i[109];
  assign o[55933] = i[109];
  assign o[55934] = i[109];
  assign o[55935] = i[109];
  assign o[55936] = i[109];
  assign o[55937] = i[109];
  assign o[55938] = i[109];
  assign o[55939] = i[109];
  assign o[55940] = i[109];
  assign o[55941] = i[109];
  assign o[55942] = i[109];
  assign o[55943] = i[109];
  assign o[55944] = i[109];
  assign o[55945] = i[109];
  assign o[55946] = i[109];
  assign o[55947] = i[109];
  assign o[55948] = i[109];
  assign o[55949] = i[109];
  assign o[55950] = i[109];
  assign o[55951] = i[109];
  assign o[55952] = i[109];
  assign o[55953] = i[109];
  assign o[55954] = i[109];
  assign o[55955] = i[109];
  assign o[55956] = i[109];
  assign o[55957] = i[109];
  assign o[55958] = i[109];
  assign o[55959] = i[109];
  assign o[55960] = i[109];
  assign o[55961] = i[109];
  assign o[55962] = i[109];
  assign o[55963] = i[109];
  assign o[55964] = i[109];
  assign o[55965] = i[109];
  assign o[55966] = i[109];
  assign o[55967] = i[109];
  assign o[55968] = i[109];
  assign o[55969] = i[109];
  assign o[55970] = i[109];
  assign o[55971] = i[109];
  assign o[55972] = i[109];
  assign o[55973] = i[109];
  assign o[55974] = i[109];
  assign o[55975] = i[109];
  assign o[55976] = i[109];
  assign o[55977] = i[109];
  assign o[55978] = i[109];
  assign o[55979] = i[109];
  assign o[55980] = i[109];
  assign o[55981] = i[109];
  assign o[55982] = i[109];
  assign o[55983] = i[109];
  assign o[55984] = i[109];
  assign o[55985] = i[109];
  assign o[55986] = i[109];
  assign o[55987] = i[109];
  assign o[55988] = i[109];
  assign o[55989] = i[109];
  assign o[55990] = i[109];
  assign o[55991] = i[109];
  assign o[55992] = i[109];
  assign o[55993] = i[109];
  assign o[55994] = i[109];
  assign o[55995] = i[109];
  assign o[55996] = i[109];
  assign o[55997] = i[109];
  assign o[55998] = i[109];
  assign o[55999] = i[109];
  assign o[56000] = i[109];
  assign o[56001] = i[109];
  assign o[56002] = i[109];
  assign o[56003] = i[109];
  assign o[56004] = i[109];
  assign o[56005] = i[109];
  assign o[56006] = i[109];
  assign o[56007] = i[109];
  assign o[56008] = i[109];
  assign o[56009] = i[109];
  assign o[56010] = i[109];
  assign o[56011] = i[109];
  assign o[56012] = i[109];
  assign o[56013] = i[109];
  assign o[56014] = i[109];
  assign o[56015] = i[109];
  assign o[56016] = i[109];
  assign o[56017] = i[109];
  assign o[56018] = i[109];
  assign o[56019] = i[109];
  assign o[56020] = i[109];
  assign o[56021] = i[109];
  assign o[56022] = i[109];
  assign o[56023] = i[109];
  assign o[56024] = i[109];
  assign o[56025] = i[109];
  assign o[56026] = i[109];
  assign o[56027] = i[109];
  assign o[56028] = i[109];
  assign o[56029] = i[109];
  assign o[56030] = i[109];
  assign o[56031] = i[109];
  assign o[56032] = i[109];
  assign o[56033] = i[109];
  assign o[56034] = i[109];
  assign o[56035] = i[109];
  assign o[56036] = i[109];
  assign o[56037] = i[109];
  assign o[56038] = i[109];
  assign o[56039] = i[109];
  assign o[56040] = i[109];
  assign o[56041] = i[109];
  assign o[56042] = i[109];
  assign o[56043] = i[109];
  assign o[56044] = i[109];
  assign o[56045] = i[109];
  assign o[56046] = i[109];
  assign o[56047] = i[109];
  assign o[56048] = i[109];
  assign o[56049] = i[109];
  assign o[56050] = i[109];
  assign o[56051] = i[109];
  assign o[56052] = i[109];
  assign o[56053] = i[109];
  assign o[56054] = i[109];
  assign o[56055] = i[109];
  assign o[56056] = i[109];
  assign o[56057] = i[109];
  assign o[56058] = i[109];
  assign o[56059] = i[109];
  assign o[56060] = i[109];
  assign o[56061] = i[109];
  assign o[56062] = i[109];
  assign o[56063] = i[109];
  assign o[56064] = i[109];
  assign o[56065] = i[109];
  assign o[56066] = i[109];
  assign o[56067] = i[109];
  assign o[56068] = i[109];
  assign o[56069] = i[109];
  assign o[56070] = i[109];
  assign o[56071] = i[109];
  assign o[56072] = i[109];
  assign o[56073] = i[109];
  assign o[56074] = i[109];
  assign o[56075] = i[109];
  assign o[56076] = i[109];
  assign o[56077] = i[109];
  assign o[56078] = i[109];
  assign o[56079] = i[109];
  assign o[56080] = i[109];
  assign o[56081] = i[109];
  assign o[56082] = i[109];
  assign o[56083] = i[109];
  assign o[56084] = i[109];
  assign o[56085] = i[109];
  assign o[56086] = i[109];
  assign o[56087] = i[109];
  assign o[56088] = i[109];
  assign o[56089] = i[109];
  assign o[56090] = i[109];
  assign o[56091] = i[109];
  assign o[56092] = i[109];
  assign o[56093] = i[109];
  assign o[56094] = i[109];
  assign o[56095] = i[109];
  assign o[56096] = i[109];
  assign o[56097] = i[109];
  assign o[56098] = i[109];
  assign o[56099] = i[109];
  assign o[56100] = i[109];
  assign o[56101] = i[109];
  assign o[56102] = i[109];
  assign o[56103] = i[109];
  assign o[56104] = i[109];
  assign o[56105] = i[109];
  assign o[56106] = i[109];
  assign o[56107] = i[109];
  assign o[56108] = i[109];
  assign o[56109] = i[109];
  assign o[56110] = i[109];
  assign o[56111] = i[109];
  assign o[56112] = i[109];
  assign o[56113] = i[109];
  assign o[56114] = i[109];
  assign o[56115] = i[109];
  assign o[56116] = i[109];
  assign o[56117] = i[109];
  assign o[56118] = i[109];
  assign o[56119] = i[109];
  assign o[56120] = i[109];
  assign o[56121] = i[109];
  assign o[56122] = i[109];
  assign o[56123] = i[109];
  assign o[56124] = i[109];
  assign o[56125] = i[109];
  assign o[56126] = i[109];
  assign o[56127] = i[109];
  assign o[56128] = i[109];
  assign o[56129] = i[109];
  assign o[56130] = i[109];
  assign o[56131] = i[109];
  assign o[56132] = i[109];
  assign o[56133] = i[109];
  assign o[56134] = i[109];
  assign o[56135] = i[109];
  assign o[56136] = i[109];
  assign o[56137] = i[109];
  assign o[56138] = i[109];
  assign o[56139] = i[109];
  assign o[56140] = i[109];
  assign o[56141] = i[109];
  assign o[56142] = i[109];
  assign o[56143] = i[109];
  assign o[56144] = i[109];
  assign o[56145] = i[109];
  assign o[56146] = i[109];
  assign o[56147] = i[109];
  assign o[56148] = i[109];
  assign o[56149] = i[109];
  assign o[56150] = i[109];
  assign o[56151] = i[109];
  assign o[56152] = i[109];
  assign o[56153] = i[109];
  assign o[56154] = i[109];
  assign o[56155] = i[109];
  assign o[56156] = i[109];
  assign o[56157] = i[109];
  assign o[56158] = i[109];
  assign o[56159] = i[109];
  assign o[56160] = i[109];
  assign o[56161] = i[109];
  assign o[56162] = i[109];
  assign o[56163] = i[109];
  assign o[56164] = i[109];
  assign o[56165] = i[109];
  assign o[56166] = i[109];
  assign o[56167] = i[109];
  assign o[56168] = i[109];
  assign o[56169] = i[109];
  assign o[56170] = i[109];
  assign o[56171] = i[109];
  assign o[56172] = i[109];
  assign o[56173] = i[109];
  assign o[56174] = i[109];
  assign o[56175] = i[109];
  assign o[56176] = i[109];
  assign o[56177] = i[109];
  assign o[56178] = i[109];
  assign o[56179] = i[109];
  assign o[56180] = i[109];
  assign o[56181] = i[109];
  assign o[56182] = i[109];
  assign o[56183] = i[109];
  assign o[56184] = i[109];
  assign o[56185] = i[109];
  assign o[56186] = i[109];
  assign o[56187] = i[109];
  assign o[56188] = i[109];
  assign o[56189] = i[109];
  assign o[56190] = i[109];
  assign o[56191] = i[109];
  assign o[56192] = i[109];
  assign o[56193] = i[109];
  assign o[56194] = i[109];
  assign o[56195] = i[109];
  assign o[56196] = i[109];
  assign o[56197] = i[109];
  assign o[56198] = i[109];
  assign o[56199] = i[109];
  assign o[56200] = i[109];
  assign o[56201] = i[109];
  assign o[56202] = i[109];
  assign o[56203] = i[109];
  assign o[56204] = i[109];
  assign o[56205] = i[109];
  assign o[56206] = i[109];
  assign o[56207] = i[109];
  assign o[56208] = i[109];
  assign o[56209] = i[109];
  assign o[56210] = i[109];
  assign o[56211] = i[109];
  assign o[56212] = i[109];
  assign o[56213] = i[109];
  assign o[56214] = i[109];
  assign o[56215] = i[109];
  assign o[56216] = i[109];
  assign o[56217] = i[109];
  assign o[56218] = i[109];
  assign o[56219] = i[109];
  assign o[56220] = i[109];
  assign o[56221] = i[109];
  assign o[56222] = i[109];
  assign o[56223] = i[109];
  assign o[56224] = i[109];
  assign o[56225] = i[109];
  assign o[56226] = i[109];
  assign o[56227] = i[109];
  assign o[56228] = i[109];
  assign o[56229] = i[109];
  assign o[56230] = i[109];
  assign o[56231] = i[109];
  assign o[56232] = i[109];
  assign o[56233] = i[109];
  assign o[56234] = i[109];
  assign o[56235] = i[109];
  assign o[56236] = i[109];
  assign o[56237] = i[109];
  assign o[56238] = i[109];
  assign o[56239] = i[109];
  assign o[56240] = i[109];
  assign o[56241] = i[109];
  assign o[56242] = i[109];
  assign o[56243] = i[109];
  assign o[56244] = i[109];
  assign o[56245] = i[109];
  assign o[56246] = i[109];
  assign o[56247] = i[109];
  assign o[56248] = i[109];
  assign o[56249] = i[109];
  assign o[56250] = i[109];
  assign o[56251] = i[109];
  assign o[56252] = i[109];
  assign o[56253] = i[109];
  assign o[56254] = i[109];
  assign o[56255] = i[109];
  assign o[56256] = i[109];
  assign o[56257] = i[109];
  assign o[56258] = i[109];
  assign o[56259] = i[109];
  assign o[56260] = i[109];
  assign o[56261] = i[109];
  assign o[56262] = i[109];
  assign o[56263] = i[109];
  assign o[56264] = i[109];
  assign o[56265] = i[109];
  assign o[56266] = i[109];
  assign o[56267] = i[109];
  assign o[56268] = i[109];
  assign o[56269] = i[109];
  assign o[56270] = i[109];
  assign o[56271] = i[109];
  assign o[56272] = i[109];
  assign o[56273] = i[109];
  assign o[56274] = i[109];
  assign o[56275] = i[109];
  assign o[56276] = i[109];
  assign o[56277] = i[109];
  assign o[56278] = i[109];
  assign o[56279] = i[109];
  assign o[56280] = i[109];
  assign o[56281] = i[109];
  assign o[56282] = i[109];
  assign o[56283] = i[109];
  assign o[56284] = i[109];
  assign o[56285] = i[109];
  assign o[56286] = i[109];
  assign o[56287] = i[109];
  assign o[56288] = i[109];
  assign o[56289] = i[109];
  assign o[56290] = i[109];
  assign o[56291] = i[109];
  assign o[56292] = i[109];
  assign o[56293] = i[109];
  assign o[56294] = i[109];
  assign o[56295] = i[109];
  assign o[56296] = i[109];
  assign o[56297] = i[109];
  assign o[56298] = i[109];
  assign o[56299] = i[109];
  assign o[56300] = i[109];
  assign o[56301] = i[109];
  assign o[56302] = i[109];
  assign o[56303] = i[109];
  assign o[56304] = i[109];
  assign o[56305] = i[109];
  assign o[56306] = i[109];
  assign o[56307] = i[109];
  assign o[56308] = i[109];
  assign o[56309] = i[109];
  assign o[56310] = i[109];
  assign o[56311] = i[109];
  assign o[56312] = i[109];
  assign o[56313] = i[109];
  assign o[56314] = i[109];
  assign o[56315] = i[109];
  assign o[56316] = i[109];
  assign o[56317] = i[109];
  assign o[56318] = i[109];
  assign o[56319] = i[109];
  assign o[55296] = i[108];
  assign o[55297] = i[108];
  assign o[55298] = i[108];
  assign o[55299] = i[108];
  assign o[55300] = i[108];
  assign o[55301] = i[108];
  assign o[55302] = i[108];
  assign o[55303] = i[108];
  assign o[55304] = i[108];
  assign o[55305] = i[108];
  assign o[55306] = i[108];
  assign o[55307] = i[108];
  assign o[55308] = i[108];
  assign o[55309] = i[108];
  assign o[55310] = i[108];
  assign o[55311] = i[108];
  assign o[55312] = i[108];
  assign o[55313] = i[108];
  assign o[55314] = i[108];
  assign o[55315] = i[108];
  assign o[55316] = i[108];
  assign o[55317] = i[108];
  assign o[55318] = i[108];
  assign o[55319] = i[108];
  assign o[55320] = i[108];
  assign o[55321] = i[108];
  assign o[55322] = i[108];
  assign o[55323] = i[108];
  assign o[55324] = i[108];
  assign o[55325] = i[108];
  assign o[55326] = i[108];
  assign o[55327] = i[108];
  assign o[55328] = i[108];
  assign o[55329] = i[108];
  assign o[55330] = i[108];
  assign o[55331] = i[108];
  assign o[55332] = i[108];
  assign o[55333] = i[108];
  assign o[55334] = i[108];
  assign o[55335] = i[108];
  assign o[55336] = i[108];
  assign o[55337] = i[108];
  assign o[55338] = i[108];
  assign o[55339] = i[108];
  assign o[55340] = i[108];
  assign o[55341] = i[108];
  assign o[55342] = i[108];
  assign o[55343] = i[108];
  assign o[55344] = i[108];
  assign o[55345] = i[108];
  assign o[55346] = i[108];
  assign o[55347] = i[108];
  assign o[55348] = i[108];
  assign o[55349] = i[108];
  assign o[55350] = i[108];
  assign o[55351] = i[108];
  assign o[55352] = i[108];
  assign o[55353] = i[108];
  assign o[55354] = i[108];
  assign o[55355] = i[108];
  assign o[55356] = i[108];
  assign o[55357] = i[108];
  assign o[55358] = i[108];
  assign o[55359] = i[108];
  assign o[55360] = i[108];
  assign o[55361] = i[108];
  assign o[55362] = i[108];
  assign o[55363] = i[108];
  assign o[55364] = i[108];
  assign o[55365] = i[108];
  assign o[55366] = i[108];
  assign o[55367] = i[108];
  assign o[55368] = i[108];
  assign o[55369] = i[108];
  assign o[55370] = i[108];
  assign o[55371] = i[108];
  assign o[55372] = i[108];
  assign o[55373] = i[108];
  assign o[55374] = i[108];
  assign o[55375] = i[108];
  assign o[55376] = i[108];
  assign o[55377] = i[108];
  assign o[55378] = i[108];
  assign o[55379] = i[108];
  assign o[55380] = i[108];
  assign o[55381] = i[108];
  assign o[55382] = i[108];
  assign o[55383] = i[108];
  assign o[55384] = i[108];
  assign o[55385] = i[108];
  assign o[55386] = i[108];
  assign o[55387] = i[108];
  assign o[55388] = i[108];
  assign o[55389] = i[108];
  assign o[55390] = i[108];
  assign o[55391] = i[108];
  assign o[55392] = i[108];
  assign o[55393] = i[108];
  assign o[55394] = i[108];
  assign o[55395] = i[108];
  assign o[55396] = i[108];
  assign o[55397] = i[108];
  assign o[55398] = i[108];
  assign o[55399] = i[108];
  assign o[55400] = i[108];
  assign o[55401] = i[108];
  assign o[55402] = i[108];
  assign o[55403] = i[108];
  assign o[55404] = i[108];
  assign o[55405] = i[108];
  assign o[55406] = i[108];
  assign o[55407] = i[108];
  assign o[55408] = i[108];
  assign o[55409] = i[108];
  assign o[55410] = i[108];
  assign o[55411] = i[108];
  assign o[55412] = i[108];
  assign o[55413] = i[108];
  assign o[55414] = i[108];
  assign o[55415] = i[108];
  assign o[55416] = i[108];
  assign o[55417] = i[108];
  assign o[55418] = i[108];
  assign o[55419] = i[108];
  assign o[55420] = i[108];
  assign o[55421] = i[108];
  assign o[55422] = i[108];
  assign o[55423] = i[108];
  assign o[55424] = i[108];
  assign o[55425] = i[108];
  assign o[55426] = i[108];
  assign o[55427] = i[108];
  assign o[55428] = i[108];
  assign o[55429] = i[108];
  assign o[55430] = i[108];
  assign o[55431] = i[108];
  assign o[55432] = i[108];
  assign o[55433] = i[108];
  assign o[55434] = i[108];
  assign o[55435] = i[108];
  assign o[55436] = i[108];
  assign o[55437] = i[108];
  assign o[55438] = i[108];
  assign o[55439] = i[108];
  assign o[55440] = i[108];
  assign o[55441] = i[108];
  assign o[55442] = i[108];
  assign o[55443] = i[108];
  assign o[55444] = i[108];
  assign o[55445] = i[108];
  assign o[55446] = i[108];
  assign o[55447] = i[108];
  assign o[55448] = i[108];
  assign o[55449] = i[108];
  assign o[55450] = i[108];
  assign o[55451] = i[108];
  assign o[55452] = i[108];
  assign o[55453] = i[108];
  assign o[55454] = i[108];
  assign o[55455] = i[108];
  assign o[55456] = i[108];
  assign o[55457] = i[108];
  assign o[55458] = i[108];
  assign o[55459] = i[108];
  assign o[55460] = i[108];
  assign o[55461] = i[108];
  assign o[55462] = i[108];
  assign o[55463] = i[108];
  assign o[55464] = i[108];
  assign o[55465] = i[108];
  assign o[55466] = i[108];
  assign o[55467] = i[108];
  assign o[55468] = i[108];
  assign o[55469] = i[108];
  assign o[55470] = i[108];
  assign o[55471] = i[108];
  assign o[55472] = i[108];
  assign o[55473] = i[108];
  assign o[55474] = i[108];
  assign o[55475] = i[108];
  assign o[55476] = i[108];
  assign o[55477] = i[108];
  assign o[55478] = i[108];
  assign o[55479] = i[108];
  assign o[55480] = i[108];
  assign o[55481] = i[108];
  assign o[55482] = i[108];
  assign o[55483] = i[108];
  assign o[55484] = i[108];
  assign o[55485] = i[108];
  assign o[55486] = i[108];
  assign o[55487] = i[108];
  assign o[55488] = i[108];
  assign o[55489] = i[108];
  assign o[55490] = i[108];
  assign o[55491] = i[108];
  assign o[55492] = i[108];
  assign o[55493] = i[108];
  assign o[55494] = i[108];
  assign o[55495] = i[108];
  assign o[55496] = i[108];
  assign o[55497] = i[108];
  assign o[55498] = i[108];
  assign o[55499] = i[108];
  assign o[55500] = i[108];
  assign o[55501] = i[108];
  assign o[55502] = i[108];
  assign o[55503] = i[108];
  assign o[55504] = i[108];
  assign o[55505] = i[108];
  assign o[55506] = i[108];
  assign o[55507] = i[108];
  assign o[55508] = i[108];
  assign o[55509] = i[108];
  assign o[55510] = i[108];
  assign o[55511] = i[108];
  assign o[55512] = i[108];
  assign o[55513] = i[108];
  assign o[55514] = i[108];
  assign o[55515] = i[108];
  assign o[55516] = i[108];
  assign o[55517] = i[108];
  assign o[55518] = i[108];
  assign o[55519] = i[108];
  assign o[55520] = i[108];
  assign o[55521] = i[108];
  assign o[55522] = i[108];
  assign o[55523] = i[108];
  assign o[55524] = i[108];
  assign o[55525] = i[108];
  assign o[55526] = i[108];
  assign o[55527] = i[108];
  assign o[55528] = i[108];
  assign o[55529] = i[108];
  assign o[55530] = i[108];
  assign o[55531] = i[108];
  assign o[55532] = i[108];
  assign o[55533] = i[108];
  assign o[55534] = i[108];
  assign o[55535] = i[108];
  assign o[55536] = i[108];
  assign o[55537] = i[108];
  assign o[55538] = i[108];
  assign o[55539] = i[108];
  assign o[55540] = i[108];
  assign o[55541] = i[108];
  assign o[55542] = i[108];
  assign o[55543] = i[108];
  assign o[55544] = i[108];
  assign o[55545] = i[108];
  assign o[55546] = i[108];
  assign o[55547] = i[108];
  assign o[55548] = i[108];
  assign o[55549] = i[108];
  assign o[55550] = i[108];
  assign o[55551] = i[108];
  assign o[55552] = i[108];
  assign o[55553] = i[108];
  assign o[55554] = i[108];
  assign o[55555] = i[108];
  assign o[55556] = i[108];
  assign o[55557] = i[108];
  assign o[55558] = i[108];
  assign o[55559] = i[108];
  assign o[55560] = i[108];
  assign o[55561] = i[108];
  assign o[55562] = i[108];
  assign o[55563] = i[108];
  assign o[55564] = i[108];
  assign o[55565] = i[108];
  assign o[55566] = i[108];
  assign o[55567] = i[108];
  assign o[55568] = i[108];
  assign o[55569] = i[108];
  assign o[55570] = i[108];
  assign o[55571] = i[108];
  assign o[55572] = i[108];
  assign o[55573] = i[108];
  assign o[55574] = i[108];
  assign o[55575] = i[108];
  assign o[55576] = i[108];
  assign o[55577] = i[108];
  assign o[55578] = i[108];
  assign o[55579] = i[108];
  assign o[55580] = i[108];
  assign o[55581] = i[108];
  assign o[55582] = i[108];
  assign o[55583] = i[108];
  assign o[55584] = i[108];
  assign o[55585] = i[108];
  assign o[55586] = i[108];
  assign o[55587] = i[108];
  assign o[55588] = i[108];
  assign o[55589] = i[108];
  assign o[55590] = i[108];
  assign o[55591] = i[108];
  assign o[55592] = i[108];
  assign o[55593] = i[108];
  assign o[55594] = i[108];
  assign o[55595] = i[108];
  assign o[55596] = i[108];
  assign o[55597] = i[108];
  assign o[55598] = i[108];
  assign o[55599] = i[108];
  assign o[55600] = i[108];
  assign o[55601] = i[108];
  assign o[55602] = i[108];
  assign o[55603] = i[108];
  assign o[55604] = i[108];
  assign o[55605] = i[108];
  assign o[55606] = i[108];
  assign o[55607] = i[108];
  assign o[55608] = i[108];
  assign o[55609] = i[108];
  assign o[55610] = i[108];
  assign o[55611] = i[108];
  assign o[55612] = i[108];
  assign o[55613] = i[108];
  assign o[55614] = i[108];
  assign o[55615] = i[108];
  assign o[55616] = i[108];
  assign o[55617] = i[108];
  assign o[55618] = i[108];
  assign o[55619] = i[108];
  assign o[55620] = i[108];
  assign o[55621] = i[108];
  assign o[55622] = i[108];
  assign o[55623] = i[108];
  assign o[55624] = i[108];
  assign o[55625] = i[108];
  assign o[55626] = i[108];
  assign o[55627] = i[108];
  assign o[55628] = i[108];
  assign o[55629] = i[108];
  assign o[55630] = i[108];
  assign o[55631] = i[108];
  assign o[55632] = i[108];
  assign o[55633] = i[108];
  assign o[55634] = i[108];
  assign o[55635] = i[108];
  assign o[55636] = i[108];
  assign o[55637] = i[108];
  assign o[55638] = i[108];
  assign o[55639] = i[108];
  assign o[55640] = i[108];
  assign o[55641] = i[108];
  assign o[55642] = i[108];
  assign o[55643] = i[108];
  assign o[55644] = i[108];
  assign o[55645] = i[108];
  assign o[55646] = i[108];
  assign o[55647] = i[108];
  assign o[55648] = i[108];
  assign o[55649] = i[108];
  assign o[55650] = i[108];
  assign o[55651] = i[108];
  assign o[55652] = i[108];
  assign o[55653] = i[108];
  assign o[55654] = i[108];
  assign o[55655] = i[108];
  assign o[55656] = i[108];
  assign o[55657] = i[108];
  assign o[55658] = i[108];
  assign o[55659] = i[108];
  assign o[55660] = i[108];
  assign o[55661] = i[108];
  assign o[55662] = i[108];
  assign o[55663] = i[108];
  assign o[55664] = i[108];
  assign o[55665] = i[108];
  assign o[55666] = i[108];
  assign o[55667] = i[108];
  assign o[55668] = i[108];
  assign o[55669] = i[108];
  assign o[55670] = i[108];
  assign o[55671] = i[108];
  assign o[55672] = i[108];
  assign o[55673] = i[108];
  assign o[55674] = i[108];
  assign o[55675] = i[108];
  assign o[55676] = i[108];
  assign o[55677] = i[108];
  assign o[55678] = i[108];
  assign o[55679] = i[108];
  assign o[55680] = i[108];
  assign o[55681] = i[108];
  assign o[55682] = i[108];
  assign o[55683] = i[108];
  assign o[55684] = i[108];
  assign o[55685] = i[108];
  assign o[55686] = i[108];
  assign o[55687] = i[108];
  assign o[55688] = i[108];
  assign o[55689] = i[108];
  assign o[55690] = i[108];
  assign o[55691] = i[108];
  assign o[55692] = i[108];
  assign o[55693] = i[108];
  assign o[55694] = i[108];
  assign o[55695] = i[108];
  assign o[55696] = i[108];
  assign o[55697] = i[108];
  assign o[55698] = i[108];
  assign o[55699] = i[108];
  assign o[55700] = i[108];
  assign o[55701] = i[108];
  assign o[55702] = i[108];
  assign o[55703] = i[108];
  assign o[55704] = i[108];
  assign o[55705] = i[108];
  assign o[55706] = i[108];
  assign o[55707] = i[108];
  assign o[55708] = i[108];
  assign o[55709] = i[108];
  assign o[55710] = i[108];
  assign o[55711] = i[108];
  assign o[55712] = i[108];
  assign o[55713] = i[108];
  assign o[55714] = i[108];
  assign o[55715] = i[108];
  assign o[55716] = i[108];
  assign o[55717] = i[108];
  assign o[55718] = i[108];
  assign o[55719] = i[108];
  assign o[55720] = i[108];
  assign o[55721] = i[108];
  assign o[55722] = i[108];
  assign o[55723] = i[108];
  assign o[55724] = i[108];
  assign o[55725] = i[108];
  assign o[55726] = i[108];
  assign o[55727] = i[108];
  assign o[55728] = i[108];
  assign o[55729] = i[108];
  assign o[55730] = i[108];
  assign o[55731] = i[108];
  assign o[55732] = i[108];
  assign o[55733] = i[108];
  assign o[55734] = i[108];
  assign o[55735] = i[108];
  assign o[55736] = i[108];
  assign o[55737] = i[108];
  assign o[55738] = i[108];
  assign o[55739] = i[108];
  assign o[55740] = i[108];
  assign o[55741] = i[108];
  assign o[55742] = i[108];
  assign o[55743] = i[108];
  assign o[55744] = i[108];
  assign o[55745] = i[108];
  assign o[55746] = i[108];
  assign o[55747] = i[108];
  assign o[55748] = i[108];
  assign o[55749] = i[108];
  assign o[55750] = i[108];
  assign o[55751] = i[108];
  assign o[55752] = i[108];
  assign o[55753] = i[108];
  assign o[55754] = i[108];
  assign o[55755] = i[108];
  assign o[55756] = i[108];
  assign o[55757] = i[108];
  assign o[55758] = i[108];
  assign o[55759] = i[108];
  assign o[55760] = i[108];
  assign o[55761] = i[108];
  assign o[55762] = i[108];
  assign o[55763] = i[108];
  assign o[55764] = i[108];
  assign o[55765] = i[108];
  assign o[55766] = i[108];
  assign o[55767] = i[108];
  assign o[55768] = i[108];
  assign o[55769] = i[108];
  assign o[55770] = i[108];
  assign o[55771] = i[108];
  assign o[55772] = i[108];
  assign o[55773] = i[108];
  assign o[55774] = i[108];
  assign o[55775] = i[108];
  assign o[55776] = i[108];
  assign o[55777] = i[108];
  assign o[55778] = i[108];
  assign o[55779] = i[108];
  assign o[55780] = i[108];
  assign o[55781] = i[108];
  assign o[55782] = i[108];
  assign o[55783] = i[108];
  assign o[55784] = i[108];
  assign o[55785] = i[108];
  assign o[55786] = i[108];
  assign o[55787] = i[108];
  assign o[55788] = i[108];
  assign o[55789] = i[108];
  assign o[55790] = i[108];
  assign o[55791] = i[108];
  assign o[55792] = i[108];
  assign o[55793] = i[108];
  assign o[55794] = i[108];
  assign o[55795] = i[108];
  assign o[55796] = i[108];
  assign o[55797] = i[108];
  assign o[55798] = i[108];
  assign o[55799] = i[108];
  assign o[55800] = i[108];
  assign o[55801] = i[108];
  assign o[55802] = i[108];
  assign o[55803] = i[108];
  assign o[55804] = i[108];
  assign o[55805] = i[108];
  assign o[55806] = i[108];
  assign o[55807] = i[108];
  assign o[54784] = i[107];
  assign o[54785] = i[107];
  assign o[54786] = i[107];
  assign o[54787] = i[107];
  assign o[54788] = i[107];
  assign o[54789] = i[107];
  assign o[54790] = i[107];
  assign o[54791] = i[107];
  assign o[54792] = i[107];
  assign o[54793] = i[107];
  assign o[54794] = i[107];
  assign o[54795] = i[107];
  assign o[54796] = i[107];
  assign o[54797] = i[107];
  assign o[54798] = i[107];
  assign o[54799] = i[107];
  assign o[54800] = i[107];
  assign o[54801] = i[107];
  assign o[54802] = i[107];
  assign o[54803] = i[107];
  assign o[54804] = i[107];
  assign o[54805] = i[107];
  assign o[54806] = i[107];
  assign o[54807] = i[107];
  assign o[54808] = i[107];
  assign o[54809] = i[107];
  assign o[54810] = i[107];
  assign o[54811] = i[107];
  assign o[54812] = i[107];
  assign o[54813] = i[107];
  assign o[54814] = i[107];
  assign o[54815] = i[107];
  assign o[54816] = i[107];
  assign o[54817] = i[107];
  assign o[54818] = i[107];
  assign o[54819] = i[107];
  assign o[54820] = i[107];
  assign o[54821] = i[107];
  assign o[54822] = i[107];
  assign o[54823] = i[107];
  assign o[54824] = i[107];
  assign o[54825] = i[107];
  assign o[54826] = i[107];
  assign o[54827] = i[107];
  assign o[54828] = i[107];
  assign o[54829] = i[107];
  assign o[54830] = i[107];
  assign o[54831] = i[107];
  assign o[54832] = i[107];
  assign o[54833] = i[107];
  assign o[54834] = i[107];
  assign o[54835] = i[107];
  assign o[54836] = i[107];
  assign o[54837] = i[107];
  assign o[54838] = i[107];
  assign o[54839] = i[107];
  assign o[54840] = i[107];
  assign o[54841] = i[107];
  assign o[54842] = i[107];
  assign o[54843] = i[107];
  assign o[54844] = i[107];
  assign o[54845] = i[107];
  assign o[54846] = i[107];
  assign o[54847] = i[107];
  assign o[54848] = i[107];
  assign o[54849] = i[107];
  assign o[54850] = i[107];
  assign o[54851] = i[107];
  assign o[54852] = i[107];
  assign o[54853] = i[107];
  assign o[54854] = i[107];
  assign o[54855] = i[107];
  assign o[54856] = i[107];
  assign o[54857] = i[107];
  assign o[54858] = i[107];
  assign o[54859] = i[107];
  assign o[54860] = i[107];
  assign o[54861] = i[107];
  assign o[54862] = i[107];
  assign o[54863] = i[107];
  assign o[54864] = i[107];
  assign o[54865] = i[107];
  assign o[54866] = i[107];
  assign o[54867] = i[107];
  assign o[54868] = i[107];
  assign o[54869] = i[107];
  assign o[54870] = i[107];
  assign o[54871] = i[107];
  assign o[54872] = i[107];
  assign o[54873] = i[107];
  assign o[54874] = i[107];
  assign o[54875] = i[107];
  assign o[54876] = i[107];
  assign o[54877] = i[107];
  assign o[54878] = i[107];
  assign o[54879] = i[107];
  assign o[54880] = i[107];
  assign o[54881] = i[107];
  assign o[54882] = i[107];
  assign o[54883] = i[107];
  assign o[54884] = i[107];
  assign o[54885] = i[107];
  assign o[54886] = i[107];
  assign o[54887] = i[107];
  assign o[54888] = i[107];
  assign o[54889] = i[107];
  assign o[54890] = i[107];
  assign o[54891] = i[107];
  assign o[54892] = i[107];
  assign o[54893] = i[107];
  assign o[54894] = i[107];
  assign o[54895] = i[107];
  assign o[54896] = i[107];
  assign o[54897] = i[107];
  assign o[54898] = i[107];
  assign o[54899] = i[107];
  assign o[54900] = i[107];
  assign o[54901] = i[107];
  assign o[54902] = i[107];
  assign o[54903] = i[107];
  assign o[54904] = i[107];
  assign o[54905] = i[107];
  assign o[54906] = i[107];
  assign o[54907] = i[107];
  assign o[54908] = i[107];
  assign o[54909] = i[107];
  assign o[54910] = i[107];
  assign o[54911] = i[107];
  assign o[54912] = i[107];
  assign o[54913] = i[107];
  assign o[54914] = i[107];
  assign o[54915] = i[107];
  assign o[54916] = i[107];
  assign o[54917] = i[107];
  assign o[54918] = i[107];
  assign o[54919] = i[107];
  assign o[54920] = i[107];
  assign o[54921] = i[107];
  assign o[54922] = i[107];
  assign o[54923] = i[107];
  assign o[54924] = i[107];
  assign o[54925] = i[107];
  assign o[54926] = i[107];
  assign o[54927] = i[107];
  assign o[54928] = i[107];
  assign o[54929] = i[107];
  assign o[54930] = i[107];
  assign o[54931] = i[107];
  assign o[54932] = i[107];
  assign o[54933] = i[107];
  assign o[54934] = i[107];
  assign o[54935] = i[107];
  assign o[54936] = i[107];
  assign o[54937] = i[107];
  assign o[54938] = i[107];
  assign o[54939] = i[107];
  assign o[54940] = i[107];
  assign o[54941] = i[107];
  assign o[54942] = i[107];
  assign o[54943] = i[107];
  assign o[54944] = i[107];
  assign o[54945] = i[107];
  assign o[54946] = i[107];
  assign o[54947] = i[107];
  assign o[54948] = i[107];
  assign o[54949] = i[107];
  assign o[54950] = i[107];
  assign o[54951] = i[107];
  assign o[54952] = i[107];
  assign o[54953] = i[107];
  assign o[54954] = i[107];
  assign o[54955] = i[107];
  assign o[54956] = i[107];
  assign o[54957] = i[107];
  assign o[54958] = i[107];
  assign o[54959] = i[107];
  assign o[54960] = i[107];
  assign o[54961] = i[107];
  assign o[54962] = i[107];
  assign o[54963] = i[107];
  assign o[54964] = i[107];
  assign o[54965] = i[107];
  assign o[54966] = i[107];
  assign o[54967] = i[107];
  assign o[54968] = i[107];
  assign o[54969] = i[107];
  assign o[54970] = i[107];
  assign o[54971] = i[107];
  assign o[54972] = i[107];
  assign o[54973] = i[107];
  assign o[54974] = i[107];
  assign o[54975] = i[107];
  assign o[54976] = i[107];
  assign o[54977] = i[107];
  assign o[54978] = i[107];
  assign o[54979] = i[107];
  assign o[54980] = i[107];
  assign o[54981] = i[107];
  assign o[54982] = i[107];
  assign o[54983] = i[107];
  assign o[54984] = i[107];
  assign o[54985] = i[107];
  assign o[54986] = i[107];
  assign o[54987] = i[107];
  assign o[54988] = i[107];
  assign o[54989] = i[107];
  assign o[54990] = i[107];
  assign o[54991] = i[107];
  assign o[54992] = i[107];
  assign o[54993] = i[107];
  assign o[54994] = i[107];
  assign o[54995] = i[107];
  assign o[54996] = i[107];
  assign o[54997] = i[107];
  assign o[54998] = i[107];
  assign o[54999] = i[107];
  assign o[55000] = i[107];
  assign o[55001] = i[107];
  assign o[55002] = i[107];
  assign o[55003] = i[107];
  assign o[55004] = i[107];
  assign o[55005] = i[107];
  assign o[55006] = i[107];
  assign o[55007] = i[107];
  assign o[55008] = i[107];
  assign o[55009] = i[107];
  assign o[55010] = i[107];
  assign o[55011] = i[107];
  assign o[55012] = i[107];
  assign o[55013] = i[107];
  assign o[55014] = i[107];
  assign o[55015] = i[107];
  assign o[55016] = i[107];
  assign o[55017] = i[107];
  assign o[55018] = i[107];
  assign o[55019] = i[107];
  assign o[55020] = i[107];
  assign o[55021] = i[107];
  assign o[55022] = i[107];
  assign o[55023] = i[107];
  assign o[55024] = i[107];
  assign o[55025] = i[107];
  assign o[55026] = i[107];
  assign o[55027] = i[107];
  assign o[55028] = i[107];
  assign o[55029] = i[107];
  assign o[55030] = i[107];
  assign o[55031] = i[107];
  assign o[55032] = i[107];
  assign o[55033] = i[107];
  assign o[55034] = i[107];
  assign o[55035] = i[107];
  assign o[55036] = i[107];
  assign o[55037] = i[107];
  assign o[55038] = i[107];
  assign o[55039] = i[107];
  assign o[55040] = i[107];
  assign o[55041] = i[107];
  assign o[55042] = i[107];
  assign o[55043] = i[107];
  assign o[55044] = i[107];
  assign o[55045] = i[107];
  assign o[55046] = i[107];
  assign o[55047] = i[107];
  assign o[55048] = i[107];
  assign o[55049] = i[107];
  assign o[55050] = i[107];
  assign o[55051] = i[107];
  assign o[55052] = i[107];
  assign o[55053] = i[107];
  assign o[55054] = i[107];
  assign o[55055] = i[107];
  assign o[55056] = i[107];
  assign o[55057] = i[107];
  assign o[55058] = i[107];
  assign o[55059] = i[107];
  assign o[55060] = i[107];
  assign o[55061] = i[107];
  assign o[55062] = i[107];
  assign o[55063] = i[107];
  assign o[55064] = i[107];
  assign o[55065] = i[107];
  assign o[55066] = i[107];
  assign o[55067] = i[107];
  assign o[55068] = i[107];
  assign o[55069] = i[107];
  assign o[55070] = i[107];
  assign o[55071] = i[107];
  assign o[55072] = i[107];
  assign o[55073] = i[107];
  assign o[55074] = i[107];
  assign o[55075] = i[107];
  assign o[55076] = i[107];
  assign o[55077] = i[107];
  assign o[55078] = i[107];
  assign o[55079] = i[107];
  assign o[55080] = i[107];
  assign o[55081] = i[107];
  assign o[55082] = i[107];
  assign o[55083] = i[107];
  assign o[55084] = i[107];
  assign o[55085] = i[107];
  assign o[55086] = i[107];
  assign o[55087] = i[107];
  assign o[55088] = i[107];
  assign o[55089] = i[107];
  assign o[55090] = i[107];
  assign o[55091] = i[107];
  assign o[55092] = i[107];
  assign o[55093] = i[107];
  assign o[55094] = i[107];
  assign o[55095] = i[107];
  assign o[55096] = i[107];
  assign o[55097] = i[107];
  assign o[55098] = i[107];
  assign o[55099] = i[107];
  assign o[55100] = i[107];
  assign o[55101] = i[107];
  assign o[55102] = i[107];
  assign o[55103] = i[107];
  assign o[55104] = i[107];
  assign o[55105] = i[107];
  assign o[55106] = i[107];
  assign o[55107] = i[107];
  assign o[55108] = i[107];
  assign o[55109] = i[107];
  assign o[55110] = i[107];
  assign o[55111] = i[107];
  assign o[55112] = i[107];
  assign o[55113] = i[107];
  assign o[55114] = i[107];
  assign o[55115] = i[107];
  assign o[55116] = i[107];
  assign o[55117] = i[107];
  assign o[55118] = i[107];
  assign o[55119] = i[107];
  assign o[55120] = i[107];
  assign o[55121] = i[107];
  assign o[55122] = i[107];
  assign o[55123] = i[107];
  assign o[55124] = i[107];
  assign o[55125] = i[107];
  assign o[55126] = i[107];
  assign o[55127] = i[107];
  assign o[55128] = i[107];
  assign o[55129] = i[107];
  assign o[55130] = i[107];
  assign o[55131] = i[107];
  assign o[55132] = i[107];
  assign o[55133] = i[107];
  assign o[55134] = i[107];
  assign o[55135] = i[107];
  assign o[55136] = i[107];
  assign o[55137] = i[107];
  assign o[55138] = i[107];
  assign o[55139] = i[107];
  assign o[55140] = i[107];
  assign o[55141] = i[107];
  assign o[55142] = i[107];
  assign o[55143] = i[107];
  assign o[55144] = i[107];
  assign o[55145] = i[107];
  assign o[55146] = i[107];
  assign o[55147] = i[107];
  assign o[55148] = i[107];
  assign o[55149] = i[107];
  assign o[55150] = i[107];
  assign o[55151] = i[107];
  assign o[55152] = i[107];
  assign o[55153] = i[107];
  assign o[55154] = i[107];
  assign o[55155] = i[107];
  assign o[55156] = i[107];
  assign o[55157] = i[107];
  assign o[55158] = i[107];
  assign o[55159] = i[107];
  assign o[55160] = i[107];
  assign o[55161] = i[107];
  assign o[55162] = i[107];
  assign o[55163] = i[107];
  assign o[55164] = i[107];
  assign o[55165] = i[107];
  assign o[55166] = i[107];
  assign o[55167] = i[107];
  assign o[55168] = i[107];
  assign o[55169] = i[107];
  assign o[55170] = i[107];
  assign o[55171] = i[107];
  assign o[55172] = i[107];
  assign o[55173] = i[107];
  assign o[55174] = i[107];
  assign o[55175] = i[107];
  assign o[55176] = i[107];
  assign o[55177] = i[107];
  assign o[55178] = i[107];
  assign o[55179] = i[107];
  assign o[55180] = i[107];
  assign o[55181] = i[107];
  assign o[55182] = i[107];
  assign o[55183] = i[107];
  assign o[55184] = i[107];
  assign o[55185] = i[107];
  assign o[55186] = i[107];
  assign o[55187] = i[107];
  assign o[55188] = i[107];
  assign o[55189] = i[107];
  assign o[55190] = i[107];
  assign o[55191] = i[107];
  assign o[55192] = i[107];
  assign o[55193] = i[107];
  assign o[55194] = i[107];
  assign o[55195] = i[107];
  assign o[55196] = i[107];
  assign o[55197] = i[107];
  assign o[55198] = i[107];
  assign o[55199] = i[107];
  assign o[55200] = i[107];
  assign o[55201] = i[107];
  assign o[55202] = i[107];
  assign o[55203] = i[107];
  assign o[55204] = i[107];
  assign o[55205] = i[107];
  assign o[55206] = i[107];
  assign o[55207] = i[107];
  assign o[55208] = i[107];
  assign o[55209] = i[107];
  assign o[55210] = i[107];
  assign o[55211] = i[107];
  assign o[55212] = i[107];
  assign o[55213] = i[107];
  assign o[55214] = i[107];
  assign o[55215] = i[107];
  assign o[55216] = i[107];
  assign o[55217] = i[107];
  assign o[55218] = i[107];
  assign o[55219] = i[107];
  assign o[55220] = i[107];
  assign o[55221] = i[107];
  assign o[55222] = i[107];
  assign o[55223] = i[107];
  assign o[55224] = i[107];
  assign o[55225] = i[107];
  assign o[55226] = i[107];
  assign o[55227] = i[107];
  assign o[55228] = i[107];
  assign o[55229] = i[107];
  assign o[55230] = i[107];
  assign o[55231] = i[107];
  assign o[55232] = i[107];
  assign o[55233] = i[107];
  assign o[55234] = i[107];
  assign o[55235] = i[107];
  assign o[55236] = i[107];
  assign o[55237] = i[107];
  assign o[55238] = i[107];
  assign o[55239] = i[107];
  assign o[55240] = i[107];
  assign o[55241] = i[107];
  assign o[55242] = i[107];
  assign o[55243] = i[107];
  assign o[55244] = i[107];
  assign o[55245] = i[107];
  assign o[55246] = i[107];
  assign o[55247] = i[107];
  assign o[55248] = i[107];
  assign o[55249] = i[107];
  assign o[55250] = i[107];
  assign o[55251] = i[107];
  assign o[55252] = i[107];
  assign o[55253] = i[107];
  assign o[55254] = i[107];
  assign o[55255] = i[107];
  assign o[55256] = i[107];
  assign o[55257] = i[107];
  assign o[55258] = i[107];
  assign o[55259] = i[107];
  assign o[55260] = i[107];
  assign o[55261] = i[107];
  assign o[55262] = i[107];
  assign o[55263] = i[107];
  assign o[55264] = i[107];
  assign o[55265] = i[107];
  assign o[55266] = i[107];
  assign o[55267] = i[107];
  assign o[55268] = i[107];
  assign o[55269] = i[107];
  assign o[55270] = i[107];
  assign o[55271] = i[107];
  assign o[55272] = i[107];
  assign o[55273] = i[107];
  assign o[55274] = i[107];
  assign o[55275] = i[107];
  assign o[55276] = i[107];
  assign o[55277] = i[107];
  assign o[55278] = i[107];
  assign o[55279] = i[107];
  assign o[55280] = i[107];
  assign o[55281] = i[107];
  assign o[55282] = i[107];
  assign o[55283] = i[107];
  assign o[55284] = i[107];
  assign o[55285] = i[107];
  assign o[55286] = i[107];
  assign o[55287] = i[107];
  assign o[55288] = i[107];
  assign o[55289] = i[107];
  assign o[55290] = i[107];
  assign o[55291] = i[107];
  assign o[55292] = i[107];
  assign o[55293] = i[107];
  assign o[55294] = i[107];
  assign o[55295] = i[107];
  assign o[54272] = i[106];
  assign o[54273] = i[106];
  assign o[54274] = i[106];
  assign o[54275] = i[106];
  assign o[54276] = i[106];
  assign o[54277] = i[106];
  assign o[54278] = i[106];
  assign o[54279] = i[106];
  assign o[54280] = i[106];
  assign o[54281] = i[106];
  assign o[54282] = i[106];
  assign o[54283] = i[106];
  assign o[54284] = i[106];
  assign o[54285] = i[106];
  assign o[54286] = i[106];
  assign o[54287] = i[106];
  assign o[54288] = i[106];
  assign o[54289] = i[106];
  assign o[54290] = i[106];
  assign o[54291] = i[106];
  assign o[54292] = i[106];
  assign o[54293] = i[106];
  assign o[54294] = i[106];
  assign o[54295] = i[106];
  assign o[54296] = i[106];
  assign o[54297] = i[106];
  assign o[54298] = i[106];
  assign o[54299] = i[106];
  assign o[54300] = i[106];
  assign o[54301] = i[106];
  assign o[54302] = i[106];
  assign o[54303] = i[106];
  assign o[54304] = i[106];
  assign o[54305] = i[106];
  assign o[54306] = i[106];
  assign o[54307] = i[106];
  assign o[54308] = i[106];
  assign o[54309] = i[106];
  assign o[54310] = i[106];
  assign o[54311] = i[106];
  assign o[54312] = i[106];
  assign o[54313] = i[106];
  assign o[54314] = i[106];
  assign o[54315] = i[106];
  assign o[54316] = i[106];
  assign o[54317] = i[106];
  assign o[54318] = i[106];
  assign o[54319] = i[106];
  assign o[54320] = i[106];
  assign o[54321] = i[106];
  assign o[54322] = i[106];
  assign o[54323] = i[106];
  assign o[54324] = i[106];
  assign o[54325] = i[106];
  assign o[54326] = i[106];
  assign o[54327] = i[106];
  assign o[54328] = i[106];
  assign o[54329] = i[106];
  assign o[54330] = i[106];
  assign o[54331] = i[106];
  assign o[54332] = i[106];
  assign o[54333] = i[106];
  assign o[54334] = i[106];
  assign o[54335] = i[106];
  assign o[54336] = i[106];
  assign o[54337] = i[106];
  assign o[54338] = i[106];
  assign o[54339] = i[106];
  assign o[54340] = i[106];
  assign o[54341] = i[106];
  assign o[54342] = i[106];
  assign o[54343] = i[106];
  assign o[54344] = i[106];
  assign o[54345] = i[106];
  assign o[54346] = i[106];
  assign o[54347] = i[106];
  assign o[54348] = i[106];
  assign o[54349] = i[106];
  assign o[54350] = i[106];
  assign o[54351] = i[106];
  assign o[54352] = i[106];
  assign o[54353] = i[106];
  assign o[54354] = i[106];
  assign o[54355] = i[106];
  assign o[54356] = i[106];
  assign o[54357] = i[106];
  assign o[54358] = i[106];
  assign o[54359] = i[106];
  assign o[54360] = i[106];
  assign o[54361] = i[106];
  assign o[54362] = i[106];
  assign o[54363] = i[106];
  assign o[54364] = i[106];
  assign o[54365] = i[106];
  assign o[54366] = i[106];
  assign o[54367] = i[106];
  assign o[54368] = i[106];
  assign o[54369] = i[106];
  assign o[54370] = i[106];
  assign o[54371] = i[106];
  assign o[54372] = i[106];
  assign o[54373] = i[106];
  assign o[54374] = i[106];
  assign o[54375] = i[106];
  assign o[54376] = i[106];
  assign o[54377] = i[106];
  assign o[54378] = i[106];
  assign o[54379] = i[106];
  assign o[54380] = i[106];
  assign o[54381] = i[106];
  assign o[54382] = i[106];
  assign o[54383] = i[106];
  assign o[54384] = i[106];
  assign o[54385] = i[106];
  assign o[54386] = i[106];
  assign o[54387] = i[106];
  assign o[54388] = i[106];
  assign o[54389] = i[106];
  assign o[54390] = i[106];
  assign o[54391] = i[106];
  assign o[54392] = i[106];
  assign o[54393] = i[106];
  assign o[54394] = i[106];
  assign o[54395] = i[106];
  assign o[54396] = i[106];
  assign o[54397] = i[106];
  assign o[54398] = i[106];
  assign o[54399] = i[106];
  assign o[54400] = i[106];
  assign o[54401] = i[106];
  assign o[54402] = i[106];
  assign o[54403] = i[106];
  assign o[54404] = i[106];
  assign o[54405] = i[106];
  assign o[54406] = i[106];
  assign o[54407] = i[106];
  assign o[54408] = i[106];
  assign o[54409] = i[106];
  assign o[54410] = i[106];
  assign o[54411] = i[106];
  assign o[54412] = i[106];
  assign o[54413] = i[106];
  assign o[54414] = i[106];
  assign o[54415] = i[106];
  assign o[54416] = i[106];
  assign o[54417] = i[106];
  assign o[54418] = i[106];
  assign o[54419] = i[106];
  assign o[54420] = i[106];
  assign o[54421] = i[106];
  assign o[54422] = i[106];
  assign o[54423] = i[106];
  assign o[54424] = i[106];
  assign o[54425] = i[106];
  assign o[54426] = i[106];
  assign o[54427] = i[106];
  assign o[54428] = i[106];
  assign o[54429] = i[106];
  assign o[54430] = i[106];
  assign o[54431] = i[106];
  assign o[54432] = i[106];
  assign o[54433] = i[106];
  assign o[54434] = i[106];
  assign o[54435] = i[106];
  assign o[54436] = i[106];
  assign o[54437] = i[106];
  assign o[54438] = i[106];
  assign o[54439] = i[106];
  assign o[54440] = i[106];
  assign o[54441] = i[106];
  assign o[54442] = i[106];
  assign o[54443] = i[106];
  assign o[54444] = i[106];
  assign o[54445] = i[106];
  assign o[54446] = i[106];
  assign o[54447] = i[106];
  assign o[54448] = i[106];
  assign o[54449] = i[106];
  assign o[54450] = i[106];
  assign o[54451] = i[106];
  assign o[54452] = i[106];
  assign o[54453] = i[106];
  assign o[54454] = i[106];
  assign o[54455] = i[106];
  assign o[54456] = i[106];
  assign o[54457] = i[106];
  assign o[54458] = i[106];
  assign o[54459] = i[106];
  assign o[54460] = i[106];
  assign o[54461] = i[106];
  assign o[54462] = i[106];
  assign o[54463] = i[106];
  assign o[54464] = i[106];
  assign o[54465] = i[106];
  assign o[54466] = i[106];
  assign o[54467] = i[106];
  assign o[54468] = i[106];
  assign o[54469] = i[106];
  assign o[54470] = i[106];
  assign o[54471] = i[106];
  assign o[54472] = i[106];
  assign o[54473] = i[106];
  assign o[54474] = i[106];
  assign o[54475] = i[106];
  assign o[54476] = i[106];
  assign o[54477] = i[106];
  assign o[54478] = i[106];
  assign o[54479] = i[106];
  assign o[54480] = i[106];
  assign o[54481] = i[106];
  assign o[54482] = i[106];
  assign o[54483] = i[106];
  assign o[54484] = i[106];
  assign o[54485] = i[106];
  assign o[54486] = i[106];
  assign o[54487] = i[106];
  assign o[54488] = i[106];
  assign o[54489] = i[106];
  assign o[54490] = i[106];
  assign o[54491] = i[106];
  assign o[54492] = i[106];
  assign o[54493] = i[106];
  assign o[54494] = i[106];
  assign o[54495] = i[106];
  assign o[54496] = i[106];
  assign o[54497] = i[106];
  assign o[54498] = i[106];
  assign o[54499] = i[106];
  assign o[54500] = i[106];
  assign o[54501] = i[106];
  assign o[54502] = i[106];
  assign o[54503] = i[106];
  assign o[54504] = i[106];
  assign o[54505] = i[106];
  assign o[54506] = i[106];
  assign o[54507] = i[106];
  assign o[54508] = i[106];
  assign o[54509] = i[106];
  assign o[54510] = i[106];
  assign o[54511] = i[106];
  assign o[54512] = i[106];
  assign o[54513] = i[106];
  assign o[54514] = i[106];
  assign o[54515] = i[106];
  assign o[54516] = i[106];
  assign o[54517] = i[106];
  assign o[54518] = i[106];
  assign o[54519] = i[106];
  assign o[54520] = i[106];
  assign o[54521] = i[106];
  assign o[54522] = i[106];
  assign o[54523] = i[106];
  assign o[54524] = i[106];
  assign o[54525] = i[106];
  assign o[54526] = i[106];
  assign o[54527] = i[106];
  assign o[54528] = i[106];
  assign o[54529] = i[106];
  assign o[54530] = i[106];
  assign o[54531] = i[106];
  assign o[54532] = i[106];
  assign o[54533] = i[106];
  assign o[54534] = i[106];
  assign o[54535] = i[106];
  assign o[54536] = i[106];
  assign o[54537] = i[106];
  assign o[54538] = i[106];
  assign o[54539] = i[106];
  assign o[54540] = i[106];
  assign o[54541] = i[106];
  assign o[54542] = i[106];
  assign o[54543] = i[106];
  assign o[54544] = i[106];
  assign o[54545] = i[106];
  assign o[54546] = i[106];
  assign o[54547] = i[106];
  assign o[54548] = i[106];
  assign o[54549] = i[106];
  assign o[54550] = i[106];
  assign o[54551] = i[106];
  assign o[54552] = i[106];
  assign o[54553] = i[106];
  assign o[54554] = i[106];
  assign o[54555] = i[106];
  assign o[54556] = i[106];
  assign o[54557] = i[106];
  assign o[54558] = i[106];
  assign o[54559] = i[106];
  assign o[54560] = i[106];
  assign o[54561] = i[106];
  assign o[54562] = i[106];
  assign o[54563] = i[106];
  assign o[54564] = i[106];
  assign o[54565] = i[106];
  assign o[54566] = i[106];
  assign o[54567] = i[106];
  assign o[54568] = i[106];
  assign o[54569] = i[106];
  assign o[54570] = i[106];
  assign o[54571] = i[106];
  assign o[54572] = i[106];
  assign o[54573] = i[106];
  assign o[54574] = i[106];
  assign o[54575] = i[106];
  assign o[54576] = i[106];
  assign o[54577] = i[106];
  assign o[54578] = i[106];
  assign o[54579] = i[106];
  assign o[54580] = i[106];
  assign o[54581] = i[106];
  assign o[54582] = i[106];
  assign o[54583] = i[106];
  assign o[54584] = i[106];
  assign o[54585] = i[106];
  assign o[54586] = i[106];
  assign o[54587] = i[106];
  assign o[54588] = i[106];
  assign o[54589] = i[106];
  assign o[54590] = i[106];
  assign o[54591] = i[106];
  assign o[54592] = i[106];
  assign o[54593] = i[106];
  assign o[54594] = i[106];
  assign o[54595] = i[106];
  assign o[54596] = i[106];
  assign o[54597] = i[106];
  assign o[54598] = i[106];
  assign o[54599] = i[106];
  assign o[54600] = i[106];
  assign o[54601] = i[106];
  assign o[54602] = i[106];
  assign o[54603] = i[106];
  assign o[54604] = i[106];
  assign o[54605] = i[106];
  assign o[54606] = i[106];
  assign o[54607] = i[106];
  assign o[54608] = i[106];
  assign o[54609] = i[106];
  assign o[54610] = i[106];
  assign o[54611] = i[106];
  assign o[54612] = i[106];
  assign o[54613] = i[106];
  assign o[54614] = i[106];
  assign o[54615] = i[106];
  assign o[54616] = i[106];
  assign o[54617] = i[106];
  assign o[54618] = i[106];
  assign o[54619] = i[106];
  assign o[54620] = i[106];
  assign o[54621] = i[106];
  assign o[54622] = i[106];
  assign o[54623] = i[106];
  assign o[54624] = i[106];
  assign o[54625] = i[106];
  assign o[54626] = i[106];
  assign o[54627] = i[106];
  assign o[54628] = i[106];
  assign o[54629] = i[106];
  assign o[54630] = i[106];
  assign o[54631] = i[106];
  assign o[54632] = i[106];
  assign o[54633] = i[106];
  assign o[54634] = i[106];
  assign o[54635] = i[106];
  assign o[54636] = i[106];
  assign o[54637] = i[106];
  assign o[54638] = i[106];
  assign o[54639] = i[106];
  assign o[54640] = i[106];
  assign o[54641] = i[106];
  assign o[54642] = i[106];
  assign o[54643] = i[106];
  assign o[54644] = i[106];
  assign o[54645] = i[106];
  assign o[54646] = i[106];
  assign o[54647] = i[106];
  assign o[54648] = i[106];
  assign o[54649] = i[106];
  assign o[54650] = i[106];
  assign o[54651] = i[106];
  assign o[54652] = i[106];
  assign o[54653] = i[106];
  assign o[54654] = i[106];
  assign o[54655] = i[106];
  assign o[54656] = i[106];
  assign o[54657] = i[106];
  assign o[54658] = i[106];
  assign o[54659] = i[106];
  assign o[54660] = i[106];
  assign o[54661] = i[106];
  assign o[54662] = i[106];
  assign o[54663] = i[106];
  assign o[54664] = i[106];
  assign o[54665] = i[106];
  assign o[54666] = i[106];
  assign o[54667] = i[106];
  assign o[54668] = i[106];
  assign o[54669] = i[106];
  assign o[54670] = i[106];
  assign o[54671] = i[106];
  assign o[54672] = i[106];
  assign o[54673] = i[106];
  assign o[54674] = i[106];
  assign o[54675] = i[106];
  assign o[54676] = i[106];
  assign o[54677] = i[106];
  assign o[54678] = i[106];
  assign o[54679] = i[106];
  assign o[54680] = i[106];
  assign o[54681] = i[106];
  assign o[54682] = i[106];
  assign o[54683] = i[106];
  assign o[54684] = i[106];
  assign o[54685] = i[106];
  assign o[54686] = i[106];
  assign o[54687] = i[106];
  assign o[54688] = i[106];
  assign o[54689] = i[106];
  assign o[54690] = i[106];
  assign o[54691] = i[106];
  assign o[54692] = i[106];
  assign o[54693] = i[106];
  assign o[54694] = i[106];
  assign o[54695] = i[106];
  assign o[54696] = i[106];
  assign o[54697] = i[106];
  assign o[54698] = i[106];
  assign o[54699] = i[106];
  assign o[54700] = i[106];
  assign o[54701] = i[106];
  assign o[54702] = i[106];
  assign o[54703] = i[106];
  assign o[54704] = i[106];
  assign o[54705] = i[106];
  assign o[54706] = i[106];
  assign o[54707] = i[106];
  assign o[54708] = i[106];
  assign o[54709] = i[106];
  assign o[54710] = i[106];
  assign o[54711] = i[106];
  assign o[54712] = i[106];
  assign o[54713] = i[106];
  assign o[54714] = i[106];
  assign o[54715] = i[106];
  assign o[54716] = i[106];
  assign o[54717] = i[106];
  assign o[54718] = i[106];
  assign o[54719] = i[106];
  assign o[54720] = i[106];
  assign o[54721] = i[106];
  assign o[54722] = i[106];
  assign o[54723] = i[106];
  assign o[54724] = i[106];
  assign o[54725] = i[106];
  assign o[54726] = i[106];
  assign o[54727] = i[106];
  assign o[54728] = i[106];
  assign o[54729] = i[106];
  assign o[54730] = i[106];
  assign o[54731] = i[106];
  assign o[54732] = i[106];
  assign o[54733] = i[106];
  assign o[54734] = i[106];
  assign o[54735] = i[106];
  assign o[54736] = i[106];
  assign o[54737] = i[106];
  assign o[54738] = i[106];
  assign o[54739] = i[106];
  assign o[54740] = i[106];
  assign o[54741] = i[106];
  assign o[54742] = i[106];
  assign o[54743] = i[106];
  assign o[54744] = i[106];
  assign o[54745] = i[106];
  assign o[54746] = i[106];
  assign o[54747] = i[106];
  assign o[54748] = i[106];
  assign o[54749] = i[106];
  assign o[54750] = i[106];
  assign o[54751] = i[106];
  assign o[54752] = i[106];
  assign o[54753] = i[106];
  assign o[54754] = i[106];
  assign o[54755] = i[106];
  assign o[54756] = i[106];
  assign o[54757] = i[106];
  assign o[54758] = i[106];
  assign o[54759] = i[106];
  assign o[54760] = i[106];
  assign o[54761] = i[106];
  assign o[54762] = i[106];
  assign o[54763] = i[106];
  assign o[54764] = i[106];
  assign o[54765] = i[106];
  assign o[54766] = i[106];
  assign o[54767] = i[106];
  assign o[54768] = i[106];
  assign o[54769] = i[106];
  assign o[54770] = i[106];
  assign o[54771] = i[106];
  assign o[54772] = i[106];
  assign o[54773] = i[106];
  assign o[54774] = i[106];
  assign o[54775] = i[106];
  assign o[54776] = i[106];
  assign o[54777] = i[106];
  assign o[54778] = i[106];
  assign o[54779] = i[106];
  assign o[54780] = i[106];
  assign o[54781] = i[106];
  assign o[54782] = i[106];
  assign o[54783] = i[106];
  assign o[53760] = i[105];
  assign o[53761] = i[105];
  assign o[53762] = i[105];
  assign o[53763] = i[105];
  assign o[53764] = i[105];
  assign o[53765] = i[105];
  assign o[53766] = i[105];
  assign o[53767] = i[105];
  assign o[53768] = i[105];
  assign o[53769] = i[105];
  assign o[53770] = i[105];
  assign o[53771] = i[105];
  assign o[53772] = i[105];
  assign o[53773] = i[105];
  assign o[53774] = i[105];
  assign o[53775] = i[105];
  assign o[53776] = i[105];
  assign o[53777] = i[105];
  assign o[53778] = i[105];
  assign o[53779] = i[105];
  assign o[53780] = i[105];
  assign o[53781] = i[105];
  assign o[53782] = i[105];
  assign o[53783] = i[105];
  assign o[53784] = i[105];
  assign o[53785] = i[105];
  assign o[53786] = i[105];
  assign o[53787] = i[105];
  assign o[53788] = i[105];
  assign o[53789] = i[105];
  assign o[53790] = i[105];
  assign o[53791] = i[105];
  assign o[53792] = i[105];
  assign o[53793] = i[105];
  assign o[53794] = i[105];
  assign o[53795] = i[105];
  assign o[53796] = i[105];
  assign o[53797] = i[105];
  assign o[53798] = i[105];
  assign o[53799] = i[105];
  assign o[53800] = i[105];
  assign o[53801] = i[105];
  assign o[53802] = i[105];
  assign o[53803] = i[105];
  assign o[53804] = i[105];
  assign o[53805] = i[105];
  assign o[53806] = i[105];
  assign o[53807] = i[105];
  assign o[53808] = i[105];
  assign o[53809] = i[105];
  assign o[53810] = i[105];
  assign o[53811] = i[105];
  assign o[53812] = i[105];
  assign o[53813] = i[105];
  assign o[53814] = i[105];
  assign o[53815] = i[105];
  assign o[53816] = i[105];
  assign o[53817] = i[105];
  assign o[53818] = i[105];
  assign o[53819] = i[105];
  assign o[53820] = i[105];
  assign o[53821] = i[105];
  assign o[53822] = i[105];
  assign o[53823] = i[105];
  assign o[53824] = i[105];
  assign o[53825] = i[105];
  assign o[53826] = i[105];
  assign o[53827] = i[105];
  assign o[53828] = i[105];
  assign o[53829] = i[105];
  assign o[53830] = i[105];
  assign o[53831] = i[105];
  assign o[53832] = i[105];
  assign o[53833] = i[105];
  assign o[53834] = i[105];
  assign o[53835] = i[105];
  assign o[53836] = i[105];
  assign o[53837] = i[105];
  assign o[53838] = i[105];
  assign o[53839] = i[105];
  assign o[53840] = i[105];
  assign o[53841] = i[105];
  assign o[53842] = i[105];
  assign o[53843] = i[105];
  assign o[53844] = i[105];
  assign o[53845] = i[105];
  assign o[53846] = i[105];
  assign o[53847] = i[105];
  assign o[53848] = i[105];
  assign o[53849] = i[105];
  assign o[53850] = i[105];
  assign o[53851] = i[105];
  assign o[53852] = i[105];
  assign o[53853] = i[105];
  assign o[53854] = i[105];
  assign o[53855] = i[105];
  assign o[53856] = i[105];
  assign o[53857] = i[105];
  assign o[53858] = i[105];
  assign o[53859] = i[105];
  assign o[53860] = i[105];
  assign o[53861] = i[105];
  assign o[53862] = i[105];
  assign o[53863] = i[105];
  assign o[53864] = i[105];
  assign o[53865] = i[105];
  assign o[53866] = i[105];
  assign o[53867] = i[105];
  assign o[53868] = i[105];
  assign o[53869] = i[105];
  assign o[53870] = i[105];
  assign o[53871] = i[105];
  assign o[53872] = i[105];
  assign o[53873] = i[105];
  assign o[53874] = i[105];
  assign o[53875] = i[105];
  assign o[53876] = i[105];
  assign o[53877] = i[105];
  assign o[53878] = i[105];
  assign o[53879] = i[105];
  assign o[53880] = i[105];
  assign o[53881] = i[105];
  assign o[53882] = i[105];
  assign o[53883] = i[105];
  assign o[53884] = i[105];
  assign o[53885] = i[105];
  assign o[53886] = i[105];
  assign o[53887] = i[105];
  assign o[53888] = i[105];
  assign o[53889] = i[105];
  assign o[53890] = i[105];
  assign o[53891] = i[105];
  assign o[53892] = i[105];
  assign o[53893] = i[105];
  assign o[53894] = i[105];
  assign o[53895] = i[105];
  assign o[53896] = i[105];
  assign o[53897] = i[105];
  assign o[53898] = i[105];
  assign o[53899] = i[105];
  assign o[53900] = i[105];
  assign o[53901] = i[105];
  assign o[53902] = i[105];
  assign o[53903] = i[105];
  assign o[53904] = i[105];
  assign o[53905] = i[105];
  assign o[53906] = i[105];
  assign o[53907] = i[105];
  assign o[53908] = i[105];
  assign o[53909] = i[105];
  assign o[53910] = i[105];
  assign o[53911] = i[105];
  assign o[53912] = i[105];
  assign o[53913] = i[105];
  assign o[53914] = i[105];
  assign o[53915] = i[105];
  assign o[53916] = i[105];
  assign o[53917] = i[105];
  assign o[53918] = i[105];
  assign o[53919] = i[105];
  assign o[53920] = i[105];
  assign o[53921] = i[105];
  assign o[53922] = i[105];
  assign o[53923] = i[105];
  assign o[53924] = i[105];
  assign o[53925] = i[105];
  assign o[53926] = i[105];
  assign o[53927] = i[105];
  assign o[53928] = i[105];
  assign o[53929] = i[105];
  assign o[53930] = i[105];
  assign o[53931] = i[105];
  assign o[53932] = i[105];
  assign o[53933] = i[105];
  assign o[53934] = i[105];
  assign o[53935] = i[105];
  assign o[53936] = i[105];
  assign o[53937] = i[105];
  assign o[53938] = i[105];
  assign o[53939] = i[105];
  assign o[53940] = i[105];
  assign o[53941] = i[105];
  assign o[53942] = i[105];
  assign o[53943] = i[105];
  assign o[53944] = i[105];
  assign o[53945] = i[105];
  assign o[53946] = i[105];
  assign o[53947] = i[105];
  assign o[53948] = i[105];
  assign o[53949] = i[105];
  assign o[53950] = i[105];
  assign o[53951] = i[105];
  assign o[53952] = i[105];
  assign o[53953] = i[105];
  assign o[53954] = i[105];
  assign o[53955] = i[105];
  assign o[53956] = i[105];
  assign o[53957] = i[105];
  assign o[53958] = i[105];
  assign o[53959] = i[105];
  assign o[53960] = i[105];
  assign o[53961] = i[105];
  assign o[53962] = i[105];
  assign o[53963] = i[105];
  assign o[53964] = i[105];
  assign o[53965] = i[105];
  assign o[53966] = i[105];
  assign o[53967] = i[105];
  assign o[53968] = i[105];
  assign o[53969] = i[105];
  assign o[53970] = i[105];
  assign o[53971] = i[105];
  assign o[53972] = i[105];
  assign o[53973] = i[105];
  assign o[53974] = i[105];
  assign o[53975] = i[105];
  assign o[53976] = i[105];
  assign o[53977] = i[105];
  assign o[53978] = i[105];
  assign o[53979] = i[105];
  assign o[53980] = i[105];
  assign o[53981] = i[105];
  assign o[53982] = i[105];
  assign o[53983] = i[105];
  assign o[53984] = i[105];
  assign o[53985] = i[105];
  assign o[53986] = i[105];
  assign o[53987] = i[105];
  assign o[53988] = i[105];
  assign o[53989] = i[105];
  assign o[53990] = i[105];
  assign o[53991] = i[105];
  assign o[53992] = i[105];
  assign o[53993] = i[105];
  assign o[53994] = i[105];
  assign o[53995] = i[105];
  assign o[53996] = i[105];
  assign o[53997] = i[105];
  assign o[53998] = i[105];
  assign o[53999] = i[105];
  assign o[54000] = i[105];
  assign o[54001] = i[105];
  assign o[54002] = i[105];
  assign o[54003] = i[105];
  assign o[54004] = i[105];
  assign o[54005] = i[105];
  assign o[54006] = i[105];
  assign o[54007] = i[105];
  assign o[54008] = i[105];
  assign o[54009] = i[105];
  assign o[54010] = i[105];
  assign o[54011] = i[105];
  assign o[54012] = i[105];
  assign o[54013] = i[105];
  assign o[54014] = i[105];
  assign o[54015] = i[105];
  assign o[54016] = i[105];
  assign o[54017] = i[105];
  assign o[54018] = i[105];
  assign o[54019] = i[105];
  assign o[54020] = i[105];
  assign o[54021] = i[105];
  assign o[54022] = i[105];
  assign o[54023] = i[105];
  assign o[54024] = i[105];
  assign o[54025] = i[105];
  assign o[54026] = i[105];
  assign o[54027] = i[105];
  assign o[54028] = i[105];
  assign o[54029] = i[105];
  assign o[54030] = i[105];
  assign o[54031] = i[105];
  assign o[54032] = i[105];
  assign o[54033] = i[105];
  assign o[54034] = i[105];
  assign o[54035] = i[105];
  assign o[54036] = i[105];
  assign o[54037] = i[105];
  assign o[54038] = i[105];
  assign o[54039] = i[105];
  assign o[54040] = i[105];
  assign o[54041] = i[105];
  assign o[54042] = i[105];
  assign o[54043] = i[105];
  assign o[54044] = i[105];
  assign o[54045] = i[105];
  assign o[54046] = i[105];
  assign o[54047] = i[105];
  assign o[54048] = i[105];
  assign o[54049] = i[105];
  assign o[54050] = i[105];
  assign o[54051] = i[105];
  assign o[54052] = i[105];
  assign o[54053] = i[105];
  assign o[54054] = i[105];
  assign o[54055] = i[105];
  assign o[54056] = i[105];
  assign o[54057] = i[105];
  assign o[54058] = i[105];
  assign o[54059] = i[105];
  assign o[54060] = i[105];
  assign o[54061] = i[105];
  assign o[54062] = i[105];
  assign o[54063] = i[105];
  assign o[54064] = i[105];
  assign o[54065] = i[105];
  assign o[54066] = i[105];
  assign o[54067] = i[105];
  assign o[54068] = i[105];
  assign o[54069] = i[105];
  assign o[54070] = i[105];
  assign o[54071] = i[105];
  assign o[54072] = i[105];
  assign o[54073] = i[105];
  assign o[54074] = i[105];
  assign o[54075] = i[105];
  assign o[54076] = i[105];
  assign o[54077] = i[105];
  assign o[54078] = i[105];
  assign o[54079] = i[105];
  assign o[54080] = i[105];
  assign o[54081] = i[105];
  assign o[54082] = i[105];
  assign o[54083] = i[105];
  assign o[54084] = i[105];
  assign o[54085] = i[105];
  assign o[54086] = i[105];
  assign o[54087] = i[105];
  assign o[54088] = i[105];
  assign o[54089] = i[105];
  assign o[54090] = i[105];
  assign o[54091] = i[105];
  assign o[54092] = i[105];
  assign o[54093] = i[105];
  assign o[54094] = i[105];
  assign o[54095] = i[105];
  assign o[54096] = i[105];
  assign o[54097] = i[105];
  assign o[54098] = i[105];
  assign o[54099] = i[105];
  assign o[54100] = i[105];
  assign o[54101] = i[105];
  assign o[54102] = i[105];
  assign o[54103] = i[105];
  assign o[54104] = i[105];
  assign o[54105] = i[105];
  assign o[54106] = i[105];
  assign o[54107] = i[105];
  assign o[54108] = i[105];
  assign o[54109] = i[105];
  assign o[54110] = i[105];
  assign o[54111] = i[105];
  assign o[54112] = i[105];
  assign o[54113] = i[105];
  assign o[54114] = i[105];
  assign o[54115] = i[105];
  assign o[54116] = i[105];
  assign o[54117] = i[105];
  assign o[54118] = i[105];
  assign o[54119] = i[105];
  assign o[54120] = i[105];
  assign o[54121] = i[105];
  assign o[54122] = i[105];
  assign o[54123] = i[105];
  assign o[54124] = i[105];
  assign o[54125] = i[105];
  assign o[54126] = i[105];
  assign o[54127] = i[105];
  assign o[54128] = i[105];
  assign o[54129] = i[105];
  assign o[54130] = i[105];
  assign o[54131] = i[105];
  assign o[54132] = i[105];
  assign o[54133] = i[105];
  assign o[54134] = i[105];
  assign o[54135] = i[105];
  assign o[54136] = i[105];
  assign o[54137] = i[105];
  assign o[54138] = i[105];
  assign o[54139] = i[105];
  assign o[54140] = i[105];
  assign o[54141] = i[105];
  assign o[54142] = i[105];
  assign o[54143] = i[105];
  assign o[54144] = i[105];
  assign o[54145] = i[105];
  assign o[54146] = i[105];
  assign o[54147] = i[105];
  assign o[54148] = i[105];
  assign o[54149] = i[105];
  assign o[54150] = i[105];
  assign o[54151] = i[105];
  assign o[54152] = i[105];
  assign o[54153] = i[105];
  assign o[54154] = i[105];
  assign o[54155] = i[105];
  assign o[54156] = i[105];
  assign o[54157] = i[105];
  assign o[54158] = i[105];
  assign o[54159] = i[105];
  assign o[54160] = i[105];
  assign o[54161] = i[105];
  assign o[54162] = i[105];
  assign o[54163] = i[105];
  assign o[54164] = i[105];
  assign o[54165] = i[105];
  assign o[54166] = i[105];
  assign o[54167] = i[105];
  assign o[54168] = i[105];
  assign o[54169] = i[105];
  assign o[54170] = i[105];
  assign o[54171] = i[105];
  assign o[54172] = i[105];
  assign o[54173] = i[105];
  assign o[54174] = i[105];
  assign o[54175] = i[105];
  assign o[54176] = i[105];
  assign o[54177] = i[105];
  assign o[54178] = i[105];
  assign o[54179] = i[105];
  assign o[54180] = i[105];
  assign o[54181] = i[105];
  assign o[54182] = i[105];
  assign o[54183] = i[105];
  assign o[54184] = i[105];
  assign o[54185] = i[105];
  assign o[54186] = i[105];
  assign o[54187] = i[105];
  assign o[54188] = i[105];
  assign o[54189] = i[105];
  assign o[54190] = i[105];
  assign o[54191] = i[105];
  assign o[54192] = i[105];
  assign o[54193] = i[105];
  assign o[54194] = i[105];
  assign o[54195] = i[105];
  assign o[54196] = i[105];
  assign o[54197] = i[105];
  assign o[54198] = i[105];
  assign o[54199] = i[105];
  assign o[54200] = i[105];
  assign o[54201] = i[105];
  assign o[54202] = i[105];
  assign o[54203] = i[105];
  assign o[54204] = i[105];
  assign o[54205] = i[105];
  assign o[54206] = i[105];
  assign o[54207] = i[105];
  assign o[54208] = i[105];
  assign o[54209] = i[105];
  assign o[54210] = i[105];
  assign o[54211] = i[105];
  assign o[54212] = i[105];
  assign o[54213] = i[105];
  assign o[54214] = i[105];
  assign o[54215] = i[105];
  assign o[54216] = i[105];
  assign o[54217] = i[105];
  assign o[54218] = i[105];
  assign o[54219] = i[105];
  assign o[54220] = i[105];
  assign o[54221] = i[105];
  assign o[54222] = i[105];
  assign o[54223] = i[105];
  assign o[54224] = i[105];
  assign o[54225] = i[105];
  assign o[54226] = i[105];
  assign o[54227] = i[105];
  assign o[54228] = i[105];
  assign o[54229] = i[105];
  assign o[54230] = i[105];
  assign o[54231] = i[105];
  assign o[54232] = i[105];
  assign o[54233] = i[105];
  assign o[54234] = i[105];
  assign o[54235] = i[105];
  assign o[54236] = i[105];
  assign o[54237] = i[105];
  assign o[54238] = i[105];
  assign o[54239] = i[105];
  assign o[54240] = i[105];
  assign o[54241] = i[105];
  assign o[54242] = i[105];
  assign o[54243] = i[105];
  assign o[54244] = i[105];
  assign o[54245] = i[105];
  assign o[54246] = i[105];
  assign o[54247] = i[105];
  assign o[54248] = i[105];
  assign o[54249] = i[105];
  assign o[54250] = i[105];
  assign o[54251] = i[105];
  assign o[54252] = i[105];
  assign o[54253] = i[105];
  assign o[54254] = i[105];
  assign o[54255] = i[105];
  assign o[54256] = i[105];
  assign o[54257] = i[105];
  assign o[54258] = i[105];
  assign o[54259] = i[105];
  assign o[54260] = i[105];
  assign o[54261] = i[105];
  assign o[54262] = i[105];
  assign o[54263] = i[105];
  assign o[54264] = i[105];
  assign o[54265] = i[105];
  assign o[54266] = i[105];
  assign o[54267] = i[105];
  assign o[54268] = i[105];
  assign o[54269] = i[105];
  assign o[54270] = i[105];
  assign o[54271] = i[105];
  assign o[53248] = i[104];
  assign o[53249] = i[104];
  assign o[53250] = i[104];
  assign o[53251] = i[104];
  assign o[53252] = i[104];
  assign o[53253] = i[104];
  assign o[53254] = i[104];
  assign o[53255] = i[104];
  assign o[53256] = i[104];
  assign o[53257] = i[104];
  assign o[53258] = i[104];
  assign o[53259] = i[104];
  assign o[53260] = i[104];
  assign o[53261] = i[104];
  assign o[53262] = i[104];
  assign o[53263] = i[104];
  assign o[53264] = i[104];
  assign o[53265] = i[104];
  assign o[53266] = i[104];
  assign o[53267] = i[104];
  assign o[53268] = i[104];
  assign o[53269] = i[104];
  assign o[53270] = i[104];
  assign o[53271] = i[104];
  assign o[53272] = i[104];
  assign o[53273] = i[104];
  assign o[53274] = i[104];
  assign o[53275] = i[104];
  assign o[53276] = i[104];
  assign o[53277] = i[104];
  assign o[53278] = i[104];
  assign o[53279] = i[104];
  assign o[53280] = i[104];
  assign o[53281] = i[104];
  assign o[53282] = i[104];
  assign o[53283] = i[104];
  assign o[53284] = i[104];
  assign o[53285] = i[104];
  assign o[53286] = i[104];
  assign o[53287] = i[104];
  assign o[53288] = i[104];
  assign o[53289] = i[104];
  assign o[53290] = i[104];
  assign o[53291] = i[104];
  assign o[53292] = i[104];
  assign o[53293] = i[104];
  assign o[53294] = i[104];
  assign o[53295] = i[104];
  assign o[53296] = i[104];
  assign o[53297] = i[104];
  assign o[53298] = i[104];
  assign o[53299] = i[104];
  assign o[53300] = i[104];
  assign o[53301] = i[104];
  assign o[53302] = i[104];
  assign o[53303] = i[104];
  assign o[53304] = i[104];
  assign o[53305] = i[104];
  assign o[53306] = i[104];
  assign o[53307] = i[104];
  assign o[53308] = i[104];
  assign o[53309] = i[104];
  assign o[53310] = i[104];
  assign o[53311] = i[104];
  assign o[53312] = i[104];
  assign o[53313] = i[104];
  assign o[53314] = i[104];
  assign o[53315] = i[104];
  assign o[53316] = i[104];
  assign o[53317] = i[104];
  assign o[53318] = i[104];
  assign o[53319] = i[104];
  assign o[53320] = i[104];
  assign o[53321] = i[104];
  assign o[53322] = i[104];
  assign o[53323] = i[104];
  assign o[53324] = i[104];
  assign o[53325] = i[104];
  assign o[53326] = i[104];
  assign o[53327] = i[104];
  assign o[53328] = i[104];
  assign o[53329] = i[104];
  assign o[53330] = i[104];
  assign o[53331] = i[104];
  assign o[53332] = i[104];
  assign o[53333] = i[104];
  assign o[53334] = i[104];
  assign o[53335] = i[104];
  assign o[53336] = i[104];
  assign o[53337] = i[104];
  assign o[53338] = i[104];
  assign o[53339] = i[104];
  assign o[53340] = i[104];
  assign o[53341] = i[104];
  assign o[53342] = i[104];
  assign o[53343] = i[104];
  assign o[53344] = i[104];
  assign o[53345] = i[104];
  assign o[53346] = i[104];
  assign o[53347] = i[104];
  assign o[53348] = i[104];
  assign o[53349] = i[104];
  assign o[53350] = i[104];
  assign o[53351] = i[104];
  assign o[53352] = i[104];
  assign o[53353] = i[104];
  assign o[53354] = i[104];
  assign o[53355] = i[104];
  assign o[53356] = i[104];
  assign o[53357] = i[104];
  assign o[53358] = i[104];
  assign o[53359] = i[104];
  assign o[53360] = i[104];
  assign o[53361] = i[104];
  assign o[53362] = i[104];
  assign o[53363] = i[104];
  assign o[53364] = i[104];
  assign o[53365] = i[104];
  assign o[53366] = i[104];
  assign o[53367] = i[104];
  assign o[53368] = i[104];
  assign o[53369] = i[104];
  assign o[53370] = i[104];
  assign o[53371] = i[104];
  assign o[53372] = i[104];
  assign o[53373] = i[104];
  assign o[53374] = i[104];
  assign o[53375] = i[104];
  assign o[53376] = i[104];
  assign o[53377] = i[104];
  assign o[53378] = i[104];
  assign o[53379] = i[104];
  assign o[53380] = i[104];
  assign o[53381] = i[104];
  assign o[53382] = i[104];
  assign o[53383] = i[104];
  assign o[53384] = i[104];
  assign o[53385] = i[104];
  assign o[53386] = i[104];
  assign o[53387] = i[104];
  assign o[53388] = i[104];
  assign o[53389] = i[104];
  assign o[53390] = i[104];
  assign o[53391] = i[104];
  assign o[53392] = i[104];
  assign o[53393] = i[104];
  assign o[53394] = i[104];
  assign o[53395] = i[104];
  assign o[53396] = i[104];
  assign o[53397] = i[104];
  assign o[53398] = i[104];
  assign o[53399] = i[104];
  assign o[53400] = i[104];
  assign o[53401] = i[104];
  assign o[53402] = i[104];
  assign o[53403] = i[104];
  assign o[53404] = i[104];
  assign o[53405] = i[104];
  assign o[53406] = i[104];
  assign o[53407] = i[104];
  assign o[53408] = i[104];
  assign o[53409] = i[104];
  assign o[53410] = i[104];
  assign o[53411] = i[104];
  assign o[53412] = i[104];
  assign o[53413] = i[104];
  assign o[53414] = i[104];
  assign o[53415] = i[104];
  assign o[53416] = i[104];
  assign o[53417] = i[104];
  assign o[53418] = i[104];
  assign o[53419] = i[104];
  assign o[53420] = i[104];
  assign o[53421] = i[104];
  assign o[53422] = i[104];
  assign o[53423] = i[104];
  assign o[53424] = i[104];
  assign o[53425] = i[104];
  assign o[53426] = i[104];
  assign o[53427] = i[104];
  assign o[53428] = i[104];
  assign o[53429] = i[104];
  assign o[53430] = i[104];
  assign o[53431] = i[104];
  assign o[53432] = i[104];
  assign o[53433] = i[104];
  assign o[53434] = i[104];
  assign o[53435] = i[104];
  assign o[53436] = i[104];
  assign o[53437] = i[104];
  assign o[53438] = i[104];
  assign o[53439] = i[104];
  assign o[53440] = i[104];
  assign o[53441] = i[104];
  assign o[53442] = i[104];
  assign o[53443] = i[104];
  assign o[53444] = i[104];
  assign o[53445] = i[104];
  assign o[53446] = i[104];
  assign o[53447] = i[104];
  assign o[53448] = i[104];
  assign o[53449] = i[104];
  assign o[53450] = i[104];
  assign o[53451] = i[104];
  assign o[53452] = i[104];
  assign o[53453] = i[104];
  assign o[53454] = i[104];
  assign o[53455] = i[104];
  assign o[53456] = i[104];
  assign o[53457] = i[104];
  assign o[53458] = i[104];
  assign o[53459] = i[104];
  assign o[53460] = i[104];
  assign o[53461] = i[104];
  assign o[53462] = i[104];
  assign o[53463] = i[104];
  assign o[53464] = i[104];
  assign o[53465] = i[104];
  assign o[53466] = i[104];
  assign o[53467] = i[104];
  assign o[53468] = i[104];
  assign o[53469] = i[104];
  assign o[53470] = i[104];
  assign o[53471] = i[104];
  assign o[53472] = i[104];
  assign o[53473] = i[104];
  assign o[53474] = i[104];
  assign o[53475] = i[104];
  assign o[53476] = i[104];
  assign o[53477] = i[104];
  assign o[53478] = i[104];
  assign o[53479] = i[104];
  assign o[53480] = i[104];
  assign o[53481] = i[104];
  assign o[53482] = i[104];
  assign o[53483] = i[104];
  assign o[53484] = i[104];
  assign o[53485] = i[104];
  assign o[53486] = i[104];
  assign o[53487] = i[104];
  assign o[53488] = i[104];
  assign o[53489] = i[104];
  assign o[53490] = i[104];
  assign o[53491] = i[104];
  assign o[53492] = i[104];
  assign o[53493] = i[104];
  assign o[53494] = i[104];
  assign o[53495] = i[104];
  assign o[53496] = i[104];
  assign o[53497] = i[104];
  assign o[53498] = i[104];
  assign o[53499] = i[104];
  assign o[53500] = i[104];
  assign o[53501] = i[104];
  assign o[53502] = i[104];
  assign o[53503] = i[104];
  assign o[53504] = i[104];
  assign o[53505] = i[104];
  assign o[53506] = i[104];
  assign o[53507] = i[104];
  assign o[53508] = i[104];
  assign o[53509] = i[104];
  assign o[53510] = i[104];
  assign o[53511] = i[104];
  assign o[53512] = i[104];
  assign o[53513] = i[104];
  assign o[53514] = i[104];
  assign o[53515] = i[104];
  assign o[53516] = i[104];
  assign o[53517] = i[104];
  assign o[53518] = i[104];
  assign o[53519] = i[104];
  assign o[53520] = i[104];
  assign o[53521] = i[104];
  assign o[53522] = i[104];
  assign o[53523] = i[104];
  assign o[53524] = i[104];
  assign o[53525] = i[104];
  assign o[53526] = i[104];
  assign o[53527] = i[104];
  assign o[53528] = i[104];
  assign o[53529] = i[104];
  assign o[53530] = i[104];
  assign o[53531] = i[104];
  assign o[53532] = i[104];
  assign o[53533] = i[104];
  assign o[53534] = i[104];
  assign o[53535] = i[104];
  assign o[53536] = i[104];
  assign o[53537] = i[104];
  assign o[53538] = i[104];
  assign o[53539] = i[104];
  assign o[53540] = i[104];
  assign o[53541] = i[104];
  assign o[53542] = i[104];
  assign o[53543] = i[104];
  assign o[53544] = i[104];
  assign o[53545] = i[104];
  assign o[53546] = i[104];
  assign o[53547] = i[104];
  assign o[53548] = i[104];
  assign o[53549] = i[104];
  assign o[53550] = i[104];
  assign o[53551] = i[104];
  assign o[53552] = i[104];
  assign o[53553] = i[104];
  assign o[53554] = i[104];
  assign o[53555] = i[104];
  assign o[53556] = i[104];
  assign o[53557] = i[104];
  assign o[53558] = i[104];
  assign o[53559] = i[104];
  assign o[53560] = i[104];
  assign o[53561] = i[104];
  assign o[53562] = i[104];
  assign o[53563] = i[104];
  assign o[53564] = i[104];
  assign o[53565] = i[104];
  assign o[53566] = i[104];
  assign o[53567] = i[104];
  assign o[53568] = i[104];
  assign o[53569] = i[104];
  assign o[53570] = i[104];
  assign o[53571] = i[104];
  assign o[53572] = i[104];
  assign o[53573] = i[104];
  assign o[53574] = i[104];
  assign o[53575] = i[104];
  assign o[53576] = i[104];
  assign o[53577] = i[104];
  assign o[53578] = i[104];
  assign o[53579] = i[104];
  assign o[53580] = i[104];
  assign o[53581] = i[104];
  assign o[53582] = i[104];
  assign o[53583] = i[104];
  assign o[53584] = i[104];
  assign o[53585] = i[104];
  assign o[53586] = i[104];
  assign o[53587] = i[104];
  assign o[53588] = i[104];
  assign o[53589] = i[104];
  assign o[53590] = i[104];
  assign o[53591] = i[104];
  assign o[53592] = i[104];
  assign o[53593] = i[104];
  assign o[53594] = i[104];
  assign o[53595] = i[104];
  assign o[53596] = i[104];
  assign o[53597] = i[104];
  assign o[53598] = i[104];
  assign o[53599] = i[104];
  assign o[53600] = i[104];
  assign o[53601] = i[104];
  assign o[53602] = i[104];
  assign o[53603] = i[104];
  assign o[53604] = i[104];
  assign o[53605] = i[104];
  assign o[53606] = i[104];
  assign o[53607] = i[104];
  assign o[53608] = i[104];
  assign o[53609] = i[104];
  assign o[53610] = i[104];
  assign o[53611] = i[104];
  assign o[53612] = i[104];
  assign o[53613] = i[104];
  assign o[53614] = i[104];
  assign o[53615] = i[104];
  assign o[53616] = i[104];
  assign o[53617] = i[104];
  assign o[53618] = i[104];
  assign o[53619] = i[104];
  assign o[53620] = i[104];
  assign o[53621] = i[104];
  assign o[53622] = i[104];
  assign o[53623] = i[104];
  assign o[53624] = i[104];
  assign o[53625] = i[104];
  assign o[53626] = i[104];
  assign o[53627] = i[104];
  assign o[53628] = i[104];
  assign o[53629] = i[104];
  assign o[53630] = i[104];
  assign o[53631] = i[104];
  assign o[53632] = i[104];
  assign o[53633] = i[104];
  assign o[53634] = i[104];
  assign o[53635] = i[104];
  assign o[53636] = i[104];
  assign o[53637] = i[104];
  assign o[53638] = i[104];
  assign o[53639] = i[104];
  assign o[53640] = i[104];
  assign o[53641] = i[104];
  assign o[53642] = i[104];
  assign o[53643] = i[104];
  assign o[53644] = i[104];
  assign o[53645] = i[104];
  assign o[53646] = i[104];
  assign o[53647] = i[104];
  assign o[53648] = i[104];
  assign o[53649] = i[104];
  assign o[53650] = i[104];
  assign o[53651] = i[104];
  assign o[53652] = i[104];
  assign o[53653] = i[104];
  assign o[53654] = i[104];
  assign o[53655] = i[104];
  assign o[53656] = i[104];
  assign o[53657] = i[104];
  assign o[53658] = i[104];
  assign o[53659] = i[104];
  assign o[53660] = i[104];
  assign o[53661] = i[104];
  assign o[53662] = i[104];
  assign o[53663] = i[104];
  assign o[53664] = i[104];
  assign o[53665] = i[104];
  assign o[53666] = i[104];
  assign o[53667] = i[104];
  assign o[53668] = i[104];
  assign o[53669] = i[104];
  assign o[53670] = i[104];
  assign o[53671] = i[104];
  assign o[53672] = i[104];
  assign o[53673] = i[104];
  assign o[53674] = i[104];
  assign o[53675] = i[104];
  assign o[53676] = i[104];
  assign o[53677] = i[104];
  assign o[53678] = i[104];
  assign o[53679] = i[104];
  assign o[53680] = i[104];
  assign o[53681] = i[104];
  assign o[53682] = i[104];
  assign o[53683] = i[104];
  assign o[53684] = i[104];
  assign o[53685] = i[104];
  assign o[53686] = i[104];
  assign o[53687] = i[104];
  assign o[53688] = i[104];
  assign o[53689] = i[104];
  assign o[53690] = i[104];
  assign o[53691] = i[104];
  assign o[53692] = i[104];
  assign o[53693] = i[104];
  assign o[53694] = i[104];
  assign o[53695] = i[104];
  assign o[53696] = i[104];
  assign o[53697] = i[104];
  assign o[53698] = i[104];
  assign o[53699] = i[104];
  assign o[53700] = i[104];
  assign o[53701] = i[104];
  assign o[53702] = i[104];
  assign o[53703] = i[104];
  assign o[53704] = i[104];
  assign o[53705] = i[104];
  assign o[53706] = i[104];
  assign o[53707] = i[104];
  assign o[53708] = i[104];
  assign o[53709] = i[104];
  assign o[53710] = i[104];
  assign o[53711] = i[104];
  assign o[53712] = i[104];
  assign o[53713] = i[104];
  assign o[53714] = i[104];
  assign o[53715] = i[104];
  assign o[53716] = i[104];
  assign o[53717] = i[104];
  assign o[53718] = i[104];
  assign o[53719] = i[104];
  assign o[53720] = i[104];
  assign o[53721] = i[104];
  assign o[53722] = i[104];
  assign o[53723] = i[104];
  assign o[53724] = i[104];
  assign o[53725] = i[104];
  assign o[53726] = i[104];
  assign o[53727] = i[104];
  assign o[53728] = i[104];
  assign o[53729] = i[104];
  assign o[53730] = i[104];
  assign o[53731] = i[104];
  assign o[53732] = i[104];
  assign o[53733] = i[104];
  assign o[53734] = i[104];
  assign o[53735] = i[104];
  assign o[53736] = i[104];
  assign o[53737] = i[104];
  assign o[53738] = i[104];
  assign o[53739] = i[104];
  assign o[53740] = i[104];
  assign o[53741] = i[104];
  assign o[53742] = i[104];
  assign o[53743] = i[104];
  assign o[53744] = i[104];
  assign o[53745] = i[104];
  assign o[53746] = i[104];
  assign o[53747] = i[104];
  assign o[53748] = i[104];
  assign o[53749] = i[104];
  assign o[53750] = i[104];
  assign o[53751] = i[104];
  assign o[53752] = i[104];
  assign o[53753] = i[104];
  assign o[53754] = i[104];
  assign o[53755] = i[104];
  assign o[53756] = i[104];
  assign o[53757] = i[104];
  assign o[53758] = i[104];
  assign o[53759] = i[104];
  assign o[52736] = i[103];
  assign o[52737] = i[103];
  assign o[52738] = i[103];
  assign o[52739] = i[103];
  assign o[52740] = i[103];
  assign o[52741] = i[103];
  assign o[52742] = i[103];
  assign o[52743] = i[103];
  assign o[52744] = i[103];
  assign o[52745] = i[103];
  assign o[52746] = i[103];
  assign o[52747] = i[103];
  assign o[52748] = i[103];
  assign o[52749] = i[103];
  assign o[52750] = i[103];
  assign o[52751] = i[103];
  assign o[52752] = i[103];
  assign o[52753] = i[103];
  assign o[52754] = i[103];
  assign o[52755] = i[103];
  assign o[52756] = i[103];
  assign o[52757] = i[103];
  assign o[52758] = i[103];
  assign o[52759] = i[103];
  assign o[52760] = i[103];
  assign o[52761] = i[103];
  assign o[52762] = i[103];
  assign o[52763] = i[103];
  assign o[52764] = i[103];
  assign o[52765] = i[103];
  assign o[52766] = i[103];
  assign o[52767] = i[103];
  assign o[52768] = i[103];
  assign o[52769] = i[103];
  assign o[52770] = i[103];
  assign o[52771] = i[103];
  assign o[52772] = i[103];
  assign o[52773] = i[103];
  assign o[52774] = i[103];
  assign o[52775] = i[103];
  assign o[52776] = i[103];
  assign o[52777] = i[103];
  assign o[52778] = i[103];
  assign o[52779] = i[103];
  assign o[52780] = i[103];
  assign o[52781] = i[103];
  assign o[52782] = i[103];
  assign o[52783] = i[103];
  assign o[52784] = i[103];
  assign o[52785] = i[103];
  assign o[52786] = i[103];
  assign o[52787] = i[103];
  assign o[52788] = i[103];
  assign o[52789] = i[103];
  assign o[52790] = i[103];
  assign o[52791] = i[103];
  assign o[52792] = i[103];
  assign o[52793] = i[103];
  assign o[52794] = i[103];
  assign o[52795] = i[103];
  assign o[52796] = i[103];
  assign o[52797] = i[103];
  assign o[52798] = i[103];
  assign o[52799] = i[103];
  assign o[52800] = i[103];
  assign o[52801] = i[103];
  assign o[52802] = i[103];
  assign o[52803] = i[103];
  assign o[52804] = i[103];
  assign o[52805] = i[103];
  assign o[52806] = i[103];
  assign o[52807] = i[103];
  assign o[52808] = i[103];
  assign o[52809] = i[103];
  assign o[52810] = i[103];
  assign o[52811] = i[103];
  assign o[52812] = i[103];
  assign o[52813] = i[103];
  assign o[52814] = i[103];
  assign o[52815] = i[103];
  assign o[52816] = i[103];
  assign o[52817] = i[103];
  assign o[52818] = i[103];
  assign o[52819] = i[103];
  assign o[52820] = i[103];
  assign o[52821] = i[103];
  assign o[52822] = i[103];
  assign o[52823] = i[103];
  assign o[52824] = i[103];
  assign o[52825] = i[103];
  assign o[52826] = i[103];
  assign o[52827] = i[103];
  assign o[52828] = i[103];
  assign o[52829] = i[103];
  assign o[52830] = i[103];
  assign o[52831] = i[103];
  assign o[52832] = i[103];
  assign o[52833] = i[103];
  assign o[52834] = i[103];
  assign o[52835] = i[103];
  assign o[52836] = i[103];
  assign o[52837] = i[103];
  assign o[52838] = i[103];
  assign o[52839] = i[103];
  assign o[52840] = i[103];
  assign o[52841] = i[103];
  assign o[52842] = i[103];
  assign o[52843] = i[103];
  assign o[52844] = i[103];
  assign o[52845] = i[103];
  assign o[52846] = i[103];
  assign o[52847] = i[103];
  assign o[52848] = i[103];
  assign o[52849] = i[103];
  assign o[52850] = i[103];
  assign o[52851] = i[103];
  assign o[52852] = i[103];
  assign o[52853] = i[103];
  assign o[52854] = i[103];
  assign o[52855] = i[103];
  assign o[52856] = i[103];
  assign o[52857] = i[103];
  assign o[52858] = i[103];
  assign o[52859] = i[103];
  assign o[52860] = i[103];
  assign o[52861] = i[103];
  assign o[52862] = i[103];
  assign o[52863] = i[103];
  assign o[52864] = i[103];
  assign o[52865] = i[103];
  assign o[52866] = i[103];
  assign o[52867] = i[103];
  assign o[52868] = i[103];
  assign o[52869] = i[103];
  assign o[52870] = i[103];
  assign o[52871] = i[103];
  assign o[52872] = i[103];
  assign o[52873] = i[103];
  assign o[52874] = i[103];
  assign o[52875] = i[103];
  assign o[52876] = i[103];
  assign o[52877] = i[103];
  assign o[52878] = i[103];
  assign o[52879] = i[103];
  assign o[52880] = i[103];
  assign o[52881] = i[103];
  assign o[52882] = i[103];
  assign o[52883] = i[103];
  assign o[52884] = i[103];
  assign o[52885] = i[103];
  assign o[52886] = i[103];
  assign o[52887] = i[103];
  assign o[52888] = i[103];
  assign o[52889] = i[103];
  assign o[52890] = i[103];
  assign o[52891] = i[103];
  assign o[52892] = i[103];
  assign o[52893] = i[103];
  assign o[52894] = i[103];
  assign o[52895] = i[103];
  assign o[52896] = i[103];
  assign o[52897] = i[103];
  assign o[52898] = i[103];
  assign o[52899] = i[103];
  assign o[52900] = i[103];
  assign o[52901] = i[103];
  assign o[52902] = i[103];
  assign o[52903] = i[103];
  assign o[52904] = i[103];
  assign o[52905] = i[103];
  assign o[52906] = i[103];
  assign o[52907] = i[103];
  assign o[52908] = i[103];
  assign o[52909] = i[103];
  assign o[52910] = i[103];
  assign o[52911] = i[103];
  assign o[52912] = i[103];
  assign o[52913] = i[103];
  assign o[52914] = i[103];
  assign o[52915] = i[103];
  assign o[52916] = i[103];
  assign o[52917] = i[103];
  assign o[52918] = i[103];
  assign o[52919] = i[103];
  assign o[52920] = i[103];
  assign o[52921] = i[103];
  assign o[52922] = i[103];
  assign o[52923] = i[103];
  assign o[52924] = i[103];
  assign o[52925] = i[103];
  assign o[52926] = i[103];
  assign o[52927] = i[103];
  assign o[52928] = i[103];
  assign o[52929] = i[103];
  assign o[52930] = i[103];
  assign o[52931] = i[103];
  assign o[52932] = i[103];
  assign o[52933] = i[103];
  assign o[52934] = i[103];
  assign o[52935] = i[103];
  assign o[52936] = i[103];
  assign o[52937] = i[103];
  assign o[52938] = i[103];
  assign o[52939] = i[103];
  assign o[52940] = i[103];
  assign o[52941] = i[103];
  assign o[52942] = i[103];
  assign o[52943] = i[103];
  assign o[52944] = i[103];
  assign o[52945] = i[103];
  assign o[52946] = i[103];
  assign o[52947] = i[103];
  assign o[52948] = i[103];
  assign o[52949] = i[103];
  assign o[52950] = i[103];
  assign o[52951] = i[103];
  assign o[52952] = i[103];
  assign o[52953] = i[103];
  assign o[52954] = i[103];
  assign o[52955] = i[103];
  assign o[52956] = i[103];
  assign o[52957] = i[103];
  assign o[52958] = i[103];
  assign o[52959] = i[103];
  assign o[52960] = i[103];
  assign o[52961] = i[103];
  assign o[52962] = i[103];
  assign o[52963] = i[103];
  assign o[52964] = i[103];
  assign o[52965] = i[103];
  assign o[52966] = i[103];
  assign o[52967] = i[103];
  assign o[52968] = i[103];
  assign o[52969] = i[103];
  assign o[52970] = i[103];
  assign o[52971] = i[103];
  assign o[52972] = i[103];
  assign o[52973] = i[103];
  assign o[52974] = i[103];
  assign o[52975] = i[103];
  assign o[52976] = i[103];
  assign o[52977] = i[103];
  assign o[52978] = i[103];
  assign o[52979] = i[103];
  assign o[52980] = i[103];
  assign o[52981] = i[103];
  assign o[52982] = i[103];
  assign o[52983] = i[103];
  assign o[52984] = i[103];
  assign o[52985] = i[103];
  assign o[52986] = i[103];
  assign o[52987] = i[103];
  assign o[52988] = i[103];
  assign o[52989] = i[103];
  assign o[52990] = i[103];
  assign o[52991] = i[103];
  assign o[52992] = i[103];
  assign o[52993] = i[103];
  assign o[52994] = i[103];
  assign o[52995] = i[103];
  assign o[52996] = i[103];
  assign o[52997] = i[103];
  assign o[52998] = i[103];
  assign o[52999] = i[103];
  assign o[53000] = i[103];
  assign o[53001] = i[103];
  assign o[53002] = i[103];
  assign o[53003] = i[103];
  assign o[53004] = i[103];
  assign o[53005] = i[103];
  assign o[53006] = i[103];
  assign o[53007] = i[103];
  assign o[53008] = i[103];
  assign o[53009] = i[103];
  assign o[53010] = i[103];
  assign o[53011] = i[103];
  assign o[53012] = i[103];
  assign o[53013] = i[103];
  assign o[53014] = i[103];
  assign o[53015] = i[103];
  assign o[53016] = i[103];
  assign o[53017] = i[103];
  assign o[53018] = i[103];
  assign o[53019] = i[103];
  assign o[53020] = i[103];
  assign o[53021] = i[103];
  assign o[53022] = i[103];
  assign o[53023] = i[103];
  assign o[53024] = i[103];
  assign o[53025] = i[103];
  assign o[53026] = i[103];
  assign o[53027] = i[103];
  assign o[53028] = i[103];
  assign o[53029] = i[103];
  assign o[53030] = i[103];
  assign o[53031] = i[103];
  assign o[53032] = i[103];
  assign o[53033] = i[103];
  assign o[53034] = i[103];
  assign o[53035] = i[103];
  assign o[53036] = i[103];
  assign o[53037] = i[103];
  assign o[53038] = i[103];
  assign o[53039] = i[103];
  assign o[53040] = i[103];
  assign o[53041] = i[103];
  assign o[53042] = i[103];
  assign o[53043] = i[103];
  assign o[53044] = i[103];
  assign o[53045] = i[103];
  assign o[53046] = i[103];
  assign o[53047] = i[103];
  assign o[53048] = i[103];
  assign o[53049] = i[103];
  assign o[53050] = i[103];
  assign o[53051] = i[103];
  assign o[53052] = i[103];
  assign o[53053] = i[103];
  assign o[53054] = i[103];
  assign o[53055] = i[103];
  assign o[53056] = i[103];
  assign o[53057] = i[103];
  assign o[53058] = i[103];
  assign o[53059] = i[103];
  assign o[53060] = i[103];
  assign o[53061] = i[103];
  assign o[53062] = i[103];
  assign o[53063] = i[103];
  assign o[53064] = i[103];
  assign o[53065] = i[103];
  assign o[53066] = i[103];
  assign o[53067] = i[103];
  assign o[53068] = i[103];
  assign o[53069] = i[103];
  assign o[53070] = i[103];
  assign o[53071] = i[103];
  assign o[53072] = i[103];
  assign o[53073] = i[103];
  assign o[53074] = i[103];
  assign o[53075] = i[103];
  assign o[53076] = i[103];
  assign o[53077] = i[103];
  assign o[53078] = i[103];
  assign o[53079] = i[103];
  assign o[53080] = i[103];
  assign o[53081] = i[103];
  assign o[53082] = i[103];
  assign o[53083] = i[103];
  assign o[53084] = i[103];
  assign o[53085] = i[103];
  assign o[53086] = i[103];
  assign o[53087] = i[103];
  assign o[53088] = i[103];
  assign o[53089] = i[103];
  assign o[53090] = i[103];
  assign o[53091] = i[103];
  assign o[53092] = i[103];
  assign o[53093] = i[103];
  assign o[53094] = i[103];
  assign o[53095] = i[103];
  assign o[53096] = i[103];
  assign o[53097] = i[103];
  assign o[53098] = i[103];
  assign o[53099] = i[103];
  assign o[53100] = i[103];
  assign o[53101] = i[103];
  assign o[53102] = i[103];
  assign o[53103] = i[103];
  assign o[53104] = i[103];
  assign o[53105] = i[103];
  assign o[53106] = i[103];
  assign o[53107] = i[103];
  assign o[53108] = i[103];
  assign o[53109] = i[103];
  assign o[53110] = i[103];
  assign o[53111] = i[103];
  assign o[53112] = i[103];
  assign o[53113] = i[103];
  assign o[53114] = i[103];
  assign o[53115] = i[103];
  assign o[53116] = i[103];
  assign o[53117] = i[103];
  assign o[53118] = i[103];
  assign o[53119] = i[103];
  assign o[53120] = i[103];
  assign o[53121] = i[103];
  assign o[53122] = i[103];
  assign o[53123] = i[103];
  assign o[53124] = i[103];
  assign o[53125] = i[103];
  assign o[53126] = i[103];
  assign o[53127] = i[103];
  assign o[53128] = i[103];
  assign o[53129] = i[103];
  assign o[53130] = i[103];
  assign o[53131] = i[103];
  assign o[53132] = i[103];
  assign o[53133] = i[103];
  assign o[53134] = i[103];
  assign o[53135] = i[103];
  assign o[53136] = i[103];
  assign o[53137] = i[103];
  assign o[53138] = i[103];
  assign o[53139] = i[103];
  assign o[53140] = i[103];
  assign o[53141] = i[103];
  assign o[53142] = i[103];
  assign o[53143] = i[103];
  assign o[53144] = i[103];
  assign o[53145] = i[103];
  assign o[53146] = i[103];
  assign o[53147] = i[103];
  assign o[53148] = i[103];
  assign o[53149] = i[103];
  assign o[53150] = i[103];
  assign o[53151] = i[103];
  assign o[53152] = i[103];
  assign o[53153] = i[103];
  assign o[53154] = i[103];
  assign o[53155] = i[103];
  assign o[53156] = i[103];
  assign o[53157] = i[103];
  assign o[53158] = i[103];
  assign o[53159] = i[103];
  assign o[53160] = i[103];
  assign o[53161] = i[103];
  assign o[53162] = i[103];
  assign o[53163] = i[103];
  assign o[53164] = i[103];
  assign o[53165] = i[103];
  assign o[53166] = i[103];
  assign o[53167] = i[103];
  assign o[53168] = i[103];
  assign o[53169] = i[103];
  assign o[53170] = i[103];
  assign o[53171] = i[103];
  assign o[53172] = i[103];
  assign o[53173] = i[103];
  assign o[53174] = i[103];
  assign o[53175] = i[103];
  assign o[53176] = i[103];
  assign o[53177] = i[103];
  assign o[53178] = i[103];
  assign o[53179] = i[103];
  assign o[53180] = i[103];
  assign o[53181] = i[103];
  assign o[53182] = i[103];
  assign o[53183] = i[103];
  assign o[53184] = i[103];
  assign o[53185] = i[103];
  assign o[53186] = i[103];
  assign o[53187] = i[103];
  assign o[53188] = i[103];
  assign o[53189] = i[103];
  assign o[53190] = i[103];
  assign o[53191] = i[103];
  assign o[53192] = i[103];
  assign o[53193] = i[103];
  assign o[53194] = i[103];
  assign o[53195] = i[103];
  assign o[53196] = i[103];
  assign o[53197] = i[103];
  assign o[53198] = i[103];
  assign o[53199] = i[103];
  assign o[53200] = i[103];
  assign o[53201] = i[103];
  assign o[53202] = i[103];
  assign o[53203] = i[103];
  assign o[53204] = i[103];
  assign o[53205] = i[103];
  assign o[53206] = i[103];
  assign o[53207] = i[103];
  assign o[53208] = i[103];
  assign o[53209] = i[103];
  assign o[53210] = i[103];
  assign o[53211] = i[103];
  assign o[53212] = i[103];
  assign o[53213] = i[103];
  assign o[53214] = i[103];
  assign o[53215] = i[103];
  assign o[53216] = i[103];
  assign o[53217] = i[103];
  assign o[53218] = i[103];
  assign o[53219] = i[103];
  assign o[53220] = i[103];
  assign o[53221] = i[103];
  assign o[53222] = i[103];
  assign o[53223] = i[103];
  assign o[53224] = i[103];
  assign o[53225] = i[103];
  assign o[53226] = i[103];
  assign o[53227] = i[103];
  assign o[53228] = i[103];
  assign o[53229] = i[103];
  assign o[53230] = i[103];
  assign o[53231] = i[103];
  assign o[53232] = i[103];
  assign o[53233] = i[103];
  assign o[53234] = i[103];
  assign o[53235] = i[103];
  assign o[53236] = i[103];
  assign o[53237] = i[103];
  assign o[53238] = i[103];
  assign o[53239] = i[103];
  assign o[53240] = i[103];
  assign o[53241] = i[103];
  assign o[53242] = i[103];
  assign o[53243] = i[103];
  assign o[53244] = i[103];
  assign o[53245] = i[103];
  assign o[53246] = i[103];
  assign o[53247] = i[103];
  assign o[52224] = i[102];
  assign o[52225] = i[102];
  assign o[52226] = i[102];
  assign o[52227] = i[102];
  assign o[52228] = i[102];
  assign o[52229] = i[102];
  assign o[52230] = i[102];
  assign o[52231] = i[102];
  assign o[52232] = i[102];
  assign o[52233] = i[102];
  assign o[52234] = i[102];
  assign o[52235] = i[102];
  assign o[52236] = i[102];
  assign o[52237] = i[102];
  assign o[52238] = i[102];
  assign o[52239] = i[102];
  assign o[52240] = i[102];
  assign o[52241] = i[102];
  assign o[52242] = i[102];
  assign o[52243] = i[102];
  assign o[52244] = i[102];
  assign o[52245] = i[102];
  assign o[52246] = i[102];
  assign o[52247] = i[102];
  assign o[52248] = i[102];
  assign o[52249] = i[102];
  assign o[52250] = i[102];
  assign o[52251] = i[102];
  assign o[52252] = i[102];
  assign o[52253] = i[102];
  assign o[52254] = i[102];
  assign o[52255] = i[102];
  assign o[52256] = i[102];
  assign o[52257] = i[102];
  assign o[52258] = i[102];
  assign o[52259] = i[102];
  assign o[52260] = i[102];
  assign o[52261] = i[102];
  assign o[52262] = i[102];
  assign o[52263] = i[102];
  assign o[52264] = i[102];
  assign o[52265] = i[102];
  assign o[52266] = i[102];
  assign o[52267] = i[102];
  assign o[52268] = i[102];
  assign o[52269] = i[102];
  assign o[52270] = i[102];
  assign o[52271] = i[102];
  assign o[52272] = i[102];
  assign o[52273] = i[102];
  assign o[52274] = i[102];
  assign o[52275] = i[102];
  assign o[52276] = i[102];
  assign o[52277] = i[102];
  assign o[52278] = i[102];
  assign o[52279] = i[102];
  assign o[52280] = i[102];
  assign o[52281] = i[102];
  assign o[52282] = i[102];
  assign o[52283] = i[102];
  assign o[52284] = i[102];
  assign o[52285] = i[102];
  assign o[52286] = i[102];
  assign o[52287] = i[102];
  assign o[52288] = i[102];
  assign o[52289] = i[102];
  assign o[52290] = i[102];
  assign o[52291] = i[102];
  assign o[52292] = i[102];
  assign o[52293] = i[102];
  assign o[52294] = i[102];
  assign o[52295] = i[102];
  assign o[52296] = i[102];
  assign o[52297] = i[102];
  assign o[52298] = i[102];
  assign o[52299] = i[102];
  assign o[52300] = i[102];
  assign o[52301] = i[102];
  assign o[52302] = i[102];
  assign o[52303] = i[102];
  assign o[52304] = i[102];
  assign o[52305] = i[102];
  assign o[52306] = i[102];
  assign o[52307] = i[102];
  assign o[52308] = i[102];
  assign o[52309] = i[102];
  assign o[52310] = i[102];
  assign o[52311] = i[102];
  assign o[52312] = i[102];
  assign o[52313] = i[102];
  assign o[52314] = i[102];
  assign o[52315] = i[102];
  assign o[52316] = i[102];
  assign o[52317] = i[102];
  assign o[52318] = i[102];
  assign o[52319] = i[102];
  assign o[52320] = i[102];
  assign o[52321] = i[102];
  assign o[52322] = i[102];
  assign o[52323] = i[102];
  assign o[52324] = i[102];
  assign o[52325] = i[102];
  assign o[52326] = i[102];
  assign o[52327] = i[102];
  assign o[52328] = i[102];
  assign o[52329] = i[102];
  assign o[52330] = i[102];
  assign o[52331] = i[102];
  assign o[52332] = i[102];
  assign o[52333] = i[102];
  assign o[52334] = i[102];
  assign o[52335] = i[102];
  assign o[52336] = i[102];
  assign o[52337] = i[102];
  assign o[52338] = i[102];
  assign o[52339] = i[102];
  assign o[52340] = i[102];
  assign o[52341] = i[102];
  assign o[52342] = i[102];
  assign o[52343] = i[102];
  assign o[52344] = i[102];
  assign o[52345] = i[102];
  assign o[52346] = i[102];
  assign o[52347] = i[102];
  assign o[52348] = i[102];
  assign o[52349] = i[102];
  assign o[52350] = i[102];
  assign o[52351] = i[102];
  assign o[52352] = i[102];
  assign o[52353] = i[102];
  assign o[52354] = i[102];
  assign o[52355] = i[102];
  assign o[52356] = i[102];
  assign o[52357] = i[102];
  assign o[52358] = i[102];
  assign o[52359] = i[102];
  assign o[52360] = i[102];
  assign o[52361] = i[102];
  assign o[52362] = i[102];
  assign o[52363] = i[102];
  assign o[52364] = i[102];
  assign o[52365] = i[102];
  assign o[52366] = i[102];
  assign o[52367] = i[102];
  assign o[52368] = i[102];
  assign o[52369] = i[102];
  assign o[52370] = i[102];
  assign o[52371] = i[102];
  assign o[52372] = i[102];
  assign o[52373] = i[102];
  assign o[52374] = i[102];
  assign o[52375] = i[102];
  assign o[52376] = i[102];
  assign o[52377] = i[102];
  assign o[52378] = i[102];
  assign o[52379] = i[102];
  assign o[52380] = i[102];
  assign o[52381] = i[102];
  assign o[52382] = i[102];
  assign o[52383] = i[102];
  assign o[52384] = i[102];
  assign o[52385] = i[102];
  assign o[52386] = i[102];
  assign o[52387] = i[102];
  assign o[52388] = i[102];
  assign o[52389] = i[102];
  assign o[52390] = i[102];
  assign o[52391] = i[102];
  assign o[52392] = i[102];
  assign o[52393] = i[102];
  assign o[52394] = i[102];
  assign o[52395] = i[102];
  assign o[52396] = i[102];
  assign o[52397] = i[102];
  assign o[52398] = i[102];
  assign o[52399] = i[102];
  assign o[52400] = i[102];
  assign o[52401] = i[102];
  assign o[52402] = i[102];
  assign o[52403] = i[102];
  assign o[52404] = i[102];
  assign o[52405] = i[102];
  assign o[52406] = i[102];
  assign o[52407] = i[102];
  assign o[52408] = i[102];
  assign o[52409] = i[102];
  assign o[52410] = i[102];
  assign o[52411] = i[102];
  assign o[52412] = i[102];
  assign o[52413] = i[102];
  assign o[52414] = i[102];
  assign o[52415] = i[102];
  assign o[52416] = i[102];
  assign o[52417] = i[102];
  assign o[52418] = i[102];
  assign o[52419] = i[102];
  assign o[52420] = i[102];
  assign o[52421] = i[102];
  assign o[52422] = i[102];
  assign o[52423] = i[102];
  assign o[52424] = i[102];
  assign o[52425] = i[102];
  assign o[52426] = i[102];
  assign o[52427] = i[102];
  assign o[52428] = i[102];
  assign o[52429] = i[102];
  assign o[52430] = i[102];
  assign o[52431] = i[102];
  assign o[52432] = i[102];
  assign o[52433] = i[102];
  assign o[52434] = i[102];
  assign o[52435] = i[102];
  assign o[52436] = i[102];
  assign o[52437] = i[102];
  assign o[52438] = i[102];
  assign o[52439] = i[102];
  assign o[52440] = i[102];
  assign o[52441] = i[102];
  assign o[52442] = i[102];
  assign o[52443] = i[102];
  assign o[52444] = i[102];
  assign o[52445] = i[102];
  assign o[52446] = i[102];
  assign o[52447] = i[102];
  assign o[52448] = i[102];
  assign o[52449] = i[102];
  assign o[52450] = i[102];
  assign o[52451] = i[102];
  assign o[52452] = i[102];
  assign o[52453] = i[102];
  assign o[52454] = i[102];
  assign o[52455] = i[102];
  assign o[52456] = i[102];
  assign o[52457] = i[102];
  assign o[52458] = i[102];
  assign o[52459] = i[102];
  assign o[52460] = i[102];
  assign o[52461] = i[102];
  assign o[52462] = i[102];
  assign o[52463] = i[102];
  assign o[52464] = i[102];
  assign o[52465] = i[102];
  assign o[52466] = i[102];
  assign o[52467] = i[102];
  assign o[52468] = i[102];
  assign o[52469] = i[102];
  assign o[52470] = i[102];
  assign o[52471] = i[102];
  assign o[52472] = i[102];
  assign o[52473] = i[102];
  assign o[52474] = i[102];
  assign o[52475] = i[102];
  assign o[52476] = i[102];
  assign o[52477] = i[102];
  assign o[52478] = i[102];
  assign o[52479] = i[102];
  assign o[52480] = i[102];
  assign o[52481] = i[102];
  assign o[52482] = i[102];
  assign o[52483] = i[102];
  assign o[52484] = i[102];
  assign o[52485] = i[102];
  assign o[52486] = i[102];
  assign o[52487] = i[102];
  assign o[52488] = i[102];
  assign o[52489] = i[102];
  assign o[52490] = i[102];
  assign o[52491] = i[102];
  assign o[52492] = i[102];
  assign o[52493] = i[102];
  assign o[52494] = i[102];
  assign o[52495] = i[102];
  assign o[52496] = i[102];
  assign o[52497] = i[102];
  assign o[52498] = i[102];
  assign o[52499] = i[102];
  assign o[52500] = i[102];
  assign o[52501] = i[102];
  assign o[52502] = i[102];
  assign o[52503] = i[102];
  assign o[52504] = i[102];
  assign o[52505] = i[102];
  assign o[52506] = i[102];
  assign o[52507] = i[102];
  assign o[52508] = i[102];
  assign o[52509] = i[102];
  assign o[52510] = i[102];
  assign o[52511] = i[102];
  assign o[52512] = i[102];
  assign o[52513] = i[102];
  assign o[52514] = i[102];
  assign o[52515] = i[102];
  assign o[52516] = i[102];
  assign o[52517] = i[102];
  assign o[52518] = i[102];
  assign o[52519] = i[102];
  assign o[52520] = i[102];
  assign o[52521] = i[102];
  assign o[52522] = i[102];
  assign o[52523] = i[102];
  assign o[52524] = i[102];
  assign o[52525] = i[102];
  assign o[52526] = i[102];
  assign o[52527] = i[102];
  assign o[52528] = i[102];
  assign o[52529] = i[102];
  assign o[52530] = i[102];
  assign o[52531] = i[102];
  assign o[52532] = i[102];
  assign o[52533] = i[102];
  assign o[52534] = i[102];
  assign o[52535] = i[102];
  assign o[52536] = i[102];
  assign o[52537] = i[102];
  assign o[52538] = i[102];
  assign o[52539] = i[102];
  assign o[52540] = i[102];
  assign o[52541] = i[102];
  assign o[52542] = i[102];
  assign o[52543] = i[102];
  assign o[52544] = i[102];
  assign o[52545] = i[102];
  assign o[52546] = i[102];
  assign o[52547] = i[102];
  assign o[52548] = i[102];
  assign o[52549] = i[102];
  assign o[52550] = i[102];
  assign o[52551] = i[102];
  assign o[52552] = i[102];
  assign o[52553] = i[102];
  assign o[52554] = i[102];
  assign o[52555] = i[102];
  assign o[52556] = i[102];
  assign o[52557] = i[102];
  assign o[52558] = i[102];
  assign o[52559] = i[102];
  assign o[52560] = i[102];
  assign o[52561] = i[102];
  assign o[52562] = i[102];
  assign o[52563] = i[102];
  assign o[52564] = i[102];
  assign o[52565] = i[102];
  assign o[52566] = i[102];
  assign o[52567] = i[102];
  assign o[52568] = i[102];
  assign o[52569] = i[102];
  assign o[52570] = i[102];
  assign o[52571] = i[102];
  assign o[52572] = i[102];
  assign o[52573] = i[102];
  assign o[52574] = i[102];
  assign o[52575] = i[102];
  assign o[52576] = i[102];
  assign o[52577] = i[102];
  assign o[52578] = i[102];
  assign o[52579] = i[102];
  assign o[52580] = i[102];
  assign o[52581] = i[102];
  assign o[52582] = i[102];
  assign o[52583] = i[102];
  assign o[52584] = i[102];
  assign o[52585] = i[102];
  assign o[52586] = i[102];
  assign o[52587] = i[102];
  assign o[52588] = i[102];
  assign o[52589] = i[102];
  assign o[52590] = i[102];
  assign o[52591] = i[102];
  assign o[52592] = i[102];
  assign o[52593] = i[102];
  assign o[52594] = i[102];
  assign o[52595] = i[102];
  assign o[52596] = i[102];
  assign o[52597] = i[102];
  assign o[52598] = i[102];
  assign o[52599] = i[102];
  assign o[52600] = i[102];
  assign o[52601] = i[102];
  assign o[52602] = i[102];
  assign o[52603] = i[102];
  assign o[52604] = i[102];
  assign o[52605] = i[102];
  assign o[52606] = i[102];
  assign o[52607] = i[102];
  assign o[52608] = i[102];
  assign o[52609] = i[102];
  assign o[52610] = i[102];
  assign o[52611] = i[102];
  assign o[52612] = i[102];
  assign o[52613] = i[102];
  assign o[52614] = i[102];
  assign o[52615] = i[102];
  assign o[52616] = i[102];
  assign o[52617] = i[102];
  assign o[52618] = i[102];
  assign o[52619] = i[102];
  assign o[52620] = i[102];
  assign o[52621] = i[102];
  assign o[52622] = i[102];
  assign o[52623] = i[102];
  assign o[52624] = i[102];
  assign o[52625] = i[102];
  assign o[52626] = i[102];
  assign o[52627] = i[102];
  assign o[52628] = i[102];
  assign o[52629] = i[102];
  assign o[52630] = i[102];
  assign o[52631] = i[102];
  assign o[52632] = i[102];
  assign o[52633] = i[102];
  assign o[52634] = i[102];
  assign o[52635] = i[102];
  assign o[52636] = i[102];
  assign o[52637] = i[102];
  assign o[52638] = i[102];
  assign o[52639] = i[102];
  assign o[52640] = i[102];
  assign o[52641] = i[102];
  assign o[52642] = i[102];
  assign o[52643] = i[102];
  assign o[52644] = i[102];
  assign o[52645] = i[102];
  assign o[52646] = i[102];
  assign o[52647] = i[102];
  assign o[52648] = i[102];
  assign o[52649] = i[102];
  assign o[52650] = i[102];
  assign o[52651] = i[102];
  assign o[52652] = i[102];
  assign o[52653] = i[102];
  assign o[52654] = i[102];
  assign o[52655] = i[102];
  assign o[52656] = i[102];
  assign o[52657] = i[102];
  assign o[52658] = i[102];
  assign o[52659] = i[102];
  assign o[52660] = i[102];
  assign o[52661] = i[102];
  assign o[52662] = i[102];
  assign o[52663] = i[102];
  assign o[52664] = i[102];
  assign o[52665] = i[102];
  assign o[52666] = i[102];
  assign o[52667] = i[102];
  assign o[52668] = i[102];
  assign o[52669] = i[102];
  assign o[52670] = i[102];
  assign o[52671] = i[102];
  assign o[52672] = i[102];
  assign o[52673] = i[102];
  assign o[52674] = i[102];
  assign o[52675] = i[102];
  assign o[52676] = i[102];
  assign o[52677] = i[102];
  assign o[52678] = i[102];
  assign o[52679] = i[102];
  assign o[52680] = i[102];
  assign o[52681] = i[102];
  assign o[52682] = i[102];
  assign o[52683] = i[102];
  assign o[52684] = i[102];
  assign o[52685] = i[102];
  assign o[52686] = i[102];
  assign o[52687] = i[102];
  assign o[52688] = i[102];
  assign o[52689] = i[102];
  assign o[52690] = i[102];
  assign o[52691] = i[102];
  assign o[52692] = i[102];
  assign o[52693] = i[102];
  assign o[52694] = i[102];
  assign o[52695] = i[102];
  assign o[52696] = i[102];
  assign o[52697] = i[102];
  assign o[52698] = i[102];
  assign o[52699] = i[102];
  assign o[52700] = i[102];
  assign o[52701] = i[102];
  assign o[52702] = i[102];
  assign o[52703] = i[102];
  assign o[52704] = i[102];
  assign o[52705] = i[102];
  assign o[52706] = i[102];
  assign o[52707] = i[102];
  assign o[52708] = i[102];
  assign o[52709] = i[102];
  assign o[52710] = i[102];
  assign o[52711] = i[102];
  assign o[52712] = i[102];
  assign o[52713] = i[102];
  assign o[52714] = i[102];
  assign o[52715] = i[102];
  assign o[52716] = i[102];
  assign o[52717] = i[102];
  assign o[52718] = i[102];
  assign o[52719] = i[102];
  assign o[52720] = i[102];
  assign o[52721] = i[102];
  assign o[52722] = i[102];
  assign o[52723] = i[102];
  assign o[52724] = i[102];
  assign o[52725] = i[102];
  assign o[52726] = i[102];
  assign o[52727] = i[102];
  assign o[52728] = i[102];
  assign o[52729] = i[102];
  assign o[52730] = i[102];
  assign o[52731] = i[102];
  assign o[52732] = i[102];
  assign o[52733] = i[102];
  assign o[52734] = i[102];
  assign o[52735] = i[102];
  assign o[51712] = i[101];
  assign o[51713] = i[101];
  assign o[51714] = i[101];
  assign o[51715] = i[101];
  assign o[51716] = i[101];
  assign o[51717] = i[101];
  assign o[51718] = i[101];
  assign o[51719] = i[101];
  assign o[51720] = i[101];
  assign o[51721] = i[101];
  assign o[51722] = i[101];
  assign o[51723] = i[101];
  assign o[51724] = i[101];
  assign o[51725] = i[101];
  assign o[51726] = i[101];
  assign o[51727] = i[101];
  assign o[51728] = i[101];
  assign o[51729] = i[101];
  assign o[51730] = i[101];
  assign o[51731] = i[101];
  assign o[51732] = i[101];
  assign o[51733] = i[101];
  assign o[51734] = i[101];
  assign o[51735] = i[101];
  assign o[51736] = i[101];
  assign o[51737] = i[101];
  assign o[51738] = i[101];
  assign o[51739] = i[101];
  assign o[51740] = i[101];
  assign o[51741] = i[101];
  assign o[51742] = i[101];
  assign o[51743] = i[101];
  assign o[51744] = i[101];
  assign o[51745] = i[101];
  assign o[51746] = i[101];
  assign o[51747] = i[101];
  assign o[51748] = i[101];
  assign o[51749] = i[101];
  assign o[51750] = i[101];
  assign o[51751] = i[101];
  assign o[51752] = i[101];
  assign o[51753] = i[101];
  assign o[51754] = i[101];
  assign o[51755] = i[101];
  assign o[51756] = i[101];
  assign o[51757] = i[101];
  assign o[51758] = i[101];
  assign o[51759] = i[101];
  assign o[51760] = i[101];
  assign o[51761] = i[101];
  assign o[51762] = i[101];
  assign o[51763] = i[101];
  assign o[51764] = i[101];
  assign o[51765] = i[101];
  assign o[51766] = i[101];
  assign o[51767] = i[101];
  assign o[51768] = i[101];
  assign o[51769] = i[101];
  assign o[51770] = i[101];
  assign o[51771] = i[101];
  assign o[51772] = i[101];
  assign o[51773] = i[101];
  assign o[51774] = i[101];
  assign o[51775] = i[101];
  assign o[51776] = i[101];
  assign o[51777] = i[101];
  assign o[51778] = i[101];
  assign o[51779] = i[101];
  assign o[51780] = i[101];
  assign o[51781] = i[101];
  assign o[51782] = i[101];
  assign o[51783] = i[101];
  assign o[51784] = i[101];
  assign o[51785] = i[101];
  assign o[51786] = i[101];
  assign o[51787] = i[101];
  assign o[51788] = i[101];
  assign o[51789] = i[101];
  assign o[51790] = i[101];
  assign o[51791] = i[101];
  assign o[51792] = i[101];
  assign o[51793] = i[101];
  assign o[51794] = i[101];
  assign o[51795] = i[101];
  assign o[51796] = i[101];
  assign o[51797] = i[101];
  assign o[51798] = i[101];
  assign o[51799] = i[101];
  assign o[51800] = i[101];
  assign o[51801] = i[101];
  assign o[51802] = i[101];
  assign o[51803] = i[101];
  assign o[51804] = i[101];
  assign o[51805] = i[101];
  assign o[51806] = i[101];
  assign o[51807] = i[101];
  assign o[51808] = i[101];
  assign o[51809] = i[101];
  assign o[51810] = i[101];
  assign o[51811] = i[101];
  assign o[51812] = i[101];
  assign o[51813] = i[101];
  assign o[51814] = i[101];
  assign o[51815] = i[101];
  assign o[51816] = i[101];
  assign o[51817] = i[101];
  assign o[51818] = i[101];
  assign o[51819] = i[101];
  assign o[51820] = i[101];
  assign o[51821] = i[101];
  assign o[51822] = i[101];
  assign o[51823] = i[101];
  assign o[51824] = i[101];
  assign o[51825] = i[101];
  assign o[51826] = i[101];
  assign o[51827] = i[101];
  assign o[51828] = i[101];
  assign o[51829] = i[101];
  assign o[51830] = i[101];
  assign o[51831] = i[101];
  assign o[51832] = i[101];
  assign o[51833] = i[101];
  assign o[51834] = i[101];
  assign o[51835] = i[101];
  assign o[51836] = i[101];
  assign o[51837] = i[101];
  assign o[51838] = i[101];
  assign o[51839] = i[101];
  assign o[51840] = i[101];
  assign o[51841] = i[101];
  assign o[51842] = i[101];
  assign o[51843] = i[101];
  assign o[51844] = i[101];
  assign o[51845] = i[101];
  assign o[51846] = i[101];
  assign o[51847] = i[101];
  assign o[51848] = i[101];
  assign o[51849] = i[101];
  assign o[51850] = i[101];
  assign o[51851] = i[101];
  assign o[51852] = i[101];
  assign o[51853] = i[101];
  assign o[51854] = i[101];
  assign o[51855] = i[101];
  assign o[51856] = i[101];
  assign o[51857] = i[101];
  assign o[51858] = i[101];
  assign o[51859] = i[101];
  assign o[51860] = i[101];
  assign o[51861] = i[101];
  assign o[51862] = i[101];
  assign o[51863] = i[101];
  assign o[51864] = i[101];
  assign o[51865] = i[101];
  assign o[51866] = i[101];
  assign o[51867] = i[101];
  assign o[51868] = i[101];
  assign o[51869] = i[101];
  assign o[51870] = i[101];
  assign o[51871] = i[101];
  assign o[51872] = i[101];
  assign o[51873] = i[101];
  assign o[51874] = i[101];
  assign o[51875] = i[101];
  assign o[51876] = i[101];
  assign o[51877] = i[101];
  assign o[51878] = i[101];
  assign o[51879] = i[101];
  assign o[51880] = i[101];
  assign o[51881] = i[101];
  assign o[51882] = i[101];
  assign o[51883] = i[101];
  assign o[51884] = i[101];
  assign o[51885] = i[101];
  assign o[51886] = i[101];
  assign o[51887] = i[101];
  assign o[51888] = i[101];
  assign o[51889] = i[101];
  assign o[51890] = i[101];
  assign o[51891] = i[101];
  assign o[51892] = i[101];
  assign o[51893] = i[101];
  assign o[51894] = i[101];
  assign o[51895] = i[101];
  assign o[51896] = i[101];
  assign o[51897] = i[101];
  assign o[51898] = i[101];
  assign o[51899] = i[101];
  assign o[51900] = i[101];
  assign o[51901] = i[101];
  assign o[51902] = i[101];
  assign o[51903] = i[101];
  assign o[51904] = i[101];
  assign o[51905] = i[101];
  assign o[51906] = i[101];
  assign o[51907] = i[101];
  assign o[51908] = i[101];
  assign o[51909] = i[101];
  assign o[51910] = i[101];
  assign o[51911] = i[101];
  assign o[51912] = i[101];
  assign o[51913] = i[101];
  assign o[51914] = i[101];
  assign o[51915] = i[101];
  assign o[51916] = i[101];
  assign o[51917] = i[101];
  assign o[51918] = i[101];
  assign o[51919] = i[101];
  assign o[51920] = i[101];
  assign o[51921] = i[101];
  assign o[51922] = i[101];
  assign o[51923] = i[101];
  assign o[51924] = i[101];
  assign o[51925] = i[101];
  assign o[51926] = i[101];
  assign o[51927] = i[101];
  assign o[51928] = i[101];
  assign o[51929] = i[101];
  assign o[51930] = i[101];
  assign o[51931] = i[101];
  assign o[51932] = i[101];
  assign o[51933] = i[101];
  assign o[51934] = i[101];
  assign o[51935] = i[101];
  assign o[51936] = i[101];
  assign o[51937] = i[101];
  assign o[51938] = i[101];
  assign o[51939] = i[101];
  assign o[51940] = i[101];
  assign o[51941] = i[101];
  assign o[51942] = i[101];
  assign o[51943] = i[101];
  assign o[51944] = i[101];
  assign o[51945] = i[101];
  assign o[51946] = i[101];
  assign o[51947] = i[101];
  assign o[51948] = i[101];
  assign o[51949] = i[101];
  assign o[51950] = i[101];
  assign o[51951] = i[101];
  assign o[51952] = i[101];
  assign o[51953] = i[101];
  assign o[51954] = i[101];
  assign o[51955] = i[101];
  assign o[51956] = i[101];
  assign o[51957] = i[101];
  assign o[51958] = i[101];
  assign o[51959] = i[101];
  assign o[51960] = i[101];
  assign o[51961] = i[101];
  assign o[51962] = i[101];
  assign o[51963] = i[101];
  assign o[51964] = i[101];
  assign o[51965] = i[101];
  assign o[51966] = i[101];
  assign o[51967] = i[101];
  assign o[51968] = i[101];
  assign o[51969] = i[101];
  assign o[51970] = i[101];
  assign o[51971] = i[101];
  assign o[51972] = i[101];
  assign o[51973] = i[101];
  assign o[51974] = i[101];
  assign o[51975] = i[101];
  assign o[51976] = i[101];
  assign o[51977] = i[101];
  assign o[51978] = i[101];
  assign o[51979] = i[101];
  assign o[51980] = i[101];
  assign o[51981] = i[101];
  assign o[51982] = i[101];
  assign o[51983] = i[101];
  assign o[51984] = i[101];
  assign o[51985] = i[101];
  assign o[51986] = i[101];
  assign o[51987] = i[101];
  assign o[51988] = i[101];
  assign o[51989] = i[101];
  assign o[51990] = i[101];
  assign o[51991] = i[101];
  assign o[51992] = i[101];
  assign o[51993] = i[101];
  assign o[51994] = i[101];
  assign o[51995] = i[101];
  assign o[51996] = i[101];
  assign o[51997] = i[101];
  assign o[51998] = i[101];
  assign o[51999] = i[101];
  assign o[52000] = i[101];
  assign o[52001] = i[101];
  assign o[52002] = i[101];
  assign o[52003] = i[101];
  assign o[52004] = i[101];
  assign o[52005] = i[101];
  assign o[52006] = i[101];
  assign o[52007] = i[101];
  assign o[52008] = i[101];
  assign o[52009] = i[101];
  assign o[52010] = i[101];
  assign o[52011] = i[101];
  assign o[52012] = i[101];
  assign o[52013] = i[101];
  assign o[52014] = i[101];
  assign o[52015] = i[101];
  assign o[52016] = i[101];
  assign o[52017] = i[101];
  assign o[52018] = i[101];
  assign o[52019] = i[101];
  assign o[52020] = i[101];
  assign o[52021] = i[101];
  assign o[52022] = i[101];
  assign o[52023] = i[101];
  assign o[52024] = i[101];
  assign o[52025] = i[101];
  assign o[52026] = i[101];
  assign o[52027] = i[101];
  assign o[52028] = i[101];
  assign o[52029] = i[101];
  assign o[52030] = i[101];
  assign o[52031] = i[101];
  assign o[52032] = i[101];
  assign o[52033] = i[101];
  assign o[52034] = i[101];
  assign o[52035] = i[101];
  assign o[52036] = i[101];
  assign o[52037] = i[101];
  assign o[52038] = i[101];
  assign o[52039] = i[101];
  assign o[52040] = i[101];
  assign o[52041] = i[101];
  assign o[52042] = i[101];
  assign o[52043] = i[101];
  assign o[52044] = i[101];
  assign o[52045] = i[101];
  assign o[52046] = i[101];
  assign o[52047] = i[101];
  assign o[52048] = i[101];
  assign o[52049] = i[101];
  assign o[52050] = i[101];
  assign o[52051] = i[101];
  assign o[52052] = i[101];
  assign o[52053] = i[101];
  assign o[52054] = i[101];
  assign o[52055] = i[101];
  assign o[52056] = i[101];
  assign o[52057] = i[101];
  assign o[52058] = i[101];
  assign o[52059] = i[101];
  assign o[52060] = i[101];
  assign o[52061] = i[101];
  assign o[52062] = i[101];
  assign o[52063] = i[101];
  assign o[52064] = i[101];
  assign o[52065] = i[101];
  assign o[52066] = i[101];
  assign o[52067] = i[101];
  assign o[52068] = i[101];
  assign o[52069] = i[101];
  assign o[52070] = i[101];
  assign o[52071] = i[101];
  assign o[52072] = i[101];
  assign o[52073] = i[101];
  assign o[52074] = i[101];
  assign o[52075] = i[101];
  assign o[52076] = i[101];
  assign o[52077] = i[101];
  assign o[52078] = i[101];
  assign o[52079] = i[101];
  assign o[52080] = i[101];
  assign o[52081] = i[101];
  assign o[52082] = i[101];
  assign o[52083] = i[101];
  assign o[52084] = i[101];
  assign o[52085] = i[101];
  assign o[52086] = i[101];
  assign o[52087] = i[101];
  assign o[52088] = i[101];
  assign o[52089] = i[101];
  assign o[52090] = i[101];
  assign o[52091] = i[101];
  assign o[52092] = i[101];
  assign o[52093] = i[101];
  assign o[52094] = i[101];
  assign o[52095] = i[101];
  assign o[52096] = i[101];
  assign o[52097] = i[101];
  assign o[52098] = i[101];
  assign o[52099] = i[101];
  assign o[52100] = i[101];
  assign o[52101] = i[101];
  assign o[52102] = i[101];
  assign o[52103] = i[101];
  assign o[52104] = i[101];
  assign o[52105] = i[101];
  assign o[52106] = i[101];
  assign o[52107] = i[101];
  assign o[52108] = i[101];
  assign o[52109] = i[101];
  assign o[52110] = i[101];
  assign o[52111] = i[101];
  assign o[52112] = i[101];
  assign o[52113] = i[101];
  assign o[52114] = i[101];
  assign o[52115] = i[101];
  assign o[52116] = i[101];
  assign o[52117] = i[101];
  assign o[52118] = i[101];
  assign o[52119] = i[101];
  assign o[52120] = i[101];
  assign o[52121] = i[101];
  assign o[52122] = i[101];
  assign o[52123] = i[101];
  assign o[52124] = i[101];
  assign o[52125] = i[101];
  assign o[52126] = i[101];
  assign o[52127] = i[101];
  assign o[52128] = i[101];
  assign o[52129] = i[101];
  assign o[52130] = i[101];
  assign o[52131] = i[101];
  assign o[52132] = i[101];
  assign o[52133] = i[101];
  assign o[52134] = i[101];
  assign o[52135] = i[101];
  assign o[52136] = i[101];
  assign o[52137] = i[101];
  assign o[52138] = i[101];
  assign o[52139] = i[101];
  assign o[52140] = i[101];
  assign o[52141] = i[101];
  assign o[52142] = i[101];
  assign o[52143] = i[101];
  assign o[52144] = i[101];
  assign o[52145] = i[101];
  assign o[52146] = i[101];
  assign o[52147] = i[101];
  assign o[52148] = i[101];
  assign o[52149] = i[101];
  assign o[52150] = i[101];
  assign o[52151] = i[101];
  assign o[52152] = i[101];
  assign o[52153] = i[101];
  assign o[52154] = i[101];
  assign o[52155] = i[101];
  assign o[52156] = i[101];
  assign o[52157] = i[101];
  assign o[52158] = i[101];
  assign o[52159] = i[101];
  assign o[52160] = i[101];
  assign o[52161] = i[101];
  assign o[52162] = i[101];
  assign o[52163] = i[101];
  assign o[52164] = i[101];
  assign o[52165] = i[101];
  assign o[52166] = i[101];
  assign o[52167] = i[101];
  assign o[52168] = i[101];
  assign o[52169] = i[101];
  assign o[52170] = i[101];
  assign o[52171] = i[101];
  assign o[52172] = i[101];
  assign o[52173] = i[101];
  assign o[52174] = i[101];
  assign o[52175] = i[101];
  assign o[52176] = i[101];
  assign o[52177] = i[101];
  assign o[52178] = i[101];
  assign o[52179] = i[101];
  assign o[52180] = i[101];
  assign o[52181] = i[101];
  assign o[52182] = i[101];
  assign o[52183] = i[101];
  assign o[52184] = i[101];
  assign o[52185] = i[101];
  assign o[52186] = i[101];
  assign o[52187] = i[101];
  assign o[52188] = i[101];
  assign o[52189] = i[101];
  assign o[52190] = i[101];
  assign o[52191] = i[101];
  assign o[52192] = i[101];
  assign o[52193] = i[101];
  assign o[52194] = i[101];
  assign o[52195] = i[101];
  assign o[52196] = i[101];
  assign o[52197] = i[101];
  assign o[52198] = i[101];
  assign o[52199] = i[101];
  assign o[52200] = i[101];
  assign o[52201] = i[101];
  assign o[52202] = i[101];
  assign o[52203] = i[101];
  assign o[52204] = i[101];
  assign o[52205] = i[101];
  assign o[52206] = i[101];
  assign o[52207] = i[101];
  assign o[52208] = i[101];
  assign o[52209] = i[101];
  assign o[52210] = i[101];
  assign o[52211] = i[101];
  assign o[52212] = i[101];
  assign o[52213] = i[101];
  assign o[52214] = i[101];
  assign o[52215] = i[101];
  assign o[52216] = i[101];
  assign o[52217] = i[101];
  assign o[52218] = i[101];
  assign o[52219] = i[101];
  assign o[52220] = i[101];
  assign o[52221] = i[101];
  assign o[52222] = i[101];
  assign o[52223] = i[101];
  assign o[51200] = i[100];
  assign o[51201] = i[100];
  assign o[51202] = i[100];
  assign o[51203] = i[100];
  assign o[51204] = i[100];
  assign o[51205] = i[100];
  assign o[51206] = i[100];
  assign o[51207] = i[100];
  assign o[51208] = i[100];
  assign o[51209] = i[100];
  assign o[51210] = i[100];
  assign o[51211] = i[100];
  assign o[51212] = i[100];
  assign o[51213] = i[100];
  assign o[51214] = i[100];
  assign o[51215] = i[100];
  assign o[51216] = i[100];
  assign o[51217] = i[100];
  assign o[51218] = i[100];
  assign o[51219] = i[100];
  assign o[51220] = i[100];
  assign o[51221] = i[100];
  assign o[51222] = i[100];
  assign o[51223] = i[100];
  assign o[51224] = i[100];
  assign o[51225] = i[100];
  assign o[51226] = i[100];
  assign o[51227] = i[100];
  assign o[51228] = i[100];
  assign o[51229] = i[100];
  assign o[51230] = i[100];
  assign o[51231] = i[100];
  assign o[51232] = i[100];
  assign o[51233] = i[100];
  assign o[51234] = i[100];
  assign o[51235] = i[100];
  assign o[51236] = i[100];
  assign o[51237] = i[100];
  assign o[51238] = i[100];
  assign o[51239] = i[100];
  assign o[51240] = i[100];
  assign o[51241] = i[100];
  assign o[51242] = i[100];
  assign o[51243] = i[100];
  assign o[51244] = i[100];
  assign o[51245] = i[100];
  assign o[51246] = i[100];
  assign o[51247] = i[100];
  assign o[51248] = i[100];
  assign o[51249] = i[100];
  assign o[51250] = i[100];
  assign o[51251] = i[100];
  assign o[51252] = i[100];
  assign o[51253] = i[100];
  assign o[51254] = i[100];
  assign o[51255] = i[100];
  assign o[51256] = i[100];
  assign o[51257] = i[100];
  assign o[51258] = i[100];
  assign o[51259] = i[100];
  assign o[51260] = i[100];
  assign o[51261] = i[100];
  assign o[51262] = i[100];
  assign o[51263] = i[100];
  assign o[51264] = i[100];
  assign o[51265] = i[100];
  assign o[51266] = i[100];
  assign o[51267] = i[100];
  assign o[51268] = i[100];
  assign o[51269] = i[100];
  assign o[51270] = i[100];
  assign o[51271] = i[100];
  assign o[51272] = i[100];
  assign o[51273] = i[100];
  assign o[51274] = i[100];
  assign o[51275] = i[100];
  assign o[51276] = i[100];
  assign o[51277] = i[100];
  assign o[51278] = i[100];
  assign o[51279] = i[100];
  assign o[51280] = i[100];
  assign o[51281] = i[100];
  assign o[51282] = i[100];
  assign o[51283] = i[100];
  assign o[51284] = i[100];
  assign o[51285] = i[100];
  assign o[51286] = i[100];
  assign o[51287] = i[100];
  assign o[51288] = i[100];
  assign o[51289] = i[100];
  assign o[51290] = i[100];
  assign o[51291] = i[100];
  assign o[51292] = i[100];
  assign o[51293] = i[100];
  assign o[51294] = i[100];
  assign o[51295] = i[100];
  assign o[51296] = i[100];
  assign o[51297] = i[100];
  assign o[51298] = i[100];
  assign o[51299] = i[100];
  assign o[51300] = i[100];
  assign o[51301] = i[100];
  assign o[51302] = i[100];
  assign o[51303] = i[100];
  assign o[51304] = i[100];
  assign o[51305] = i[100];
  assign o[51306] = i[100];
  assign o[51307] = i[100];
  assign o[51308] = i[100];
  assign o[51309] = i[100];
  assign o[51310] = i[100];
  assign o[51311] = i[100];
  assign o[51312] = i[100];
  assign o[51313] = i[100];
  assign o[51314] = i[100];
  assign o[51315] = i[100];
  assign o[51316] = i[100];
  assign o[51317] = i[100];
  assign o[51318] = i[100];
  assign o[51319] = i[100];
  assign o[51320] = i[100];
  assign o[51321] = i[100];
  assign o[51322] = i[100];
  assign o[51323] = i[100];
  assign o[51324] = i[100];
  assign o[51325] = i[100];
  assign o[51326] = i[100];
  assign o[51327] = i[100];
  assign o[51328] = i[100];
  assign o[51329] = i[100];
  assign o[51330] = i[100];
  assign o[51331] = i[100];
  assign o[51332] = i[100];
  assign o[51333] = i[100];
  assign o[51334] = i[100];
  assign o[51335] = i[100];
  assign o[51336] = i[100];
  assign o[51337] = i[100];
  assign o[51338] = i[100];
  assign o[51339] = i[100];
  assign o[51340] = i[100];
  assign o[51341] = i[100];
  assign o[51342] = i[100];
  assign o[51343] = i[100];
  assign o[51344] = i[100];
  assign o[51345] = i[100];
  assign o[51346] = i[100];
  assign o[51347] = i[100];
  assign o[51348] = i[100];
  assign o[51349] = i[100];
  assign o[51350] = i[100];
  assign o[51351] = i[100];
  assign o[51352] = i[100];
  assign o[51353] = i[100];
  assign o[51354] = i[100];
  assign o[51355] = i[100];
  assign o[51356] = i[100];
  assign o[51357] = i[100];
  assign o[51358] = i[100];
  assign o[51359] = i[100];
  assign o[51360] = i[100];
  assign o[51361] = i[100];
  assign o[51362] = i[100];
  assign o[51363] = i[100];
  assign o[51364] = i[100];
  assign o[51365] = i[100];
  assign o[51366] = i[100];
  assign o[51367] = i[100];
  assign o[51368] = i[100];
  assign o[51369] = i[100];
  assign o[51370] = i[100];
  assign o[51371] = i[100];
  assign o[51372] = i[100];
  assign o[51373] = i[100];
  assign o[51374] = i[100];
  assign o[51375] = i[100];
  assign o[51376] = i[100];
  assign o[51377] = i[100];
  assign o[51378] = i[100];
  assign o[51379] = i[100];
  assign o[51380] = i[100];
  assign o[51381] = i[100];
  assign o[51382] = i[100];
  assign o[51383] = i[100];
  assign o[51384] = i[100];
  assign o[51385] = i[100];
  assign o[51386] = i[100];
  assign o[51387] = i[100];
  assign o[51388] = i[100];
  assign o[51389] = i[100];
  assign o[51390] = i[100];
  assign o[51391] = i[100];
  assign o[51392] = i[100];
  assign o[51393] = i[100];
  assign o[51394] = i[100];
  assign o[51395] = i[100];
  assign o[51396] = i[100];
  assign o[51397] = i[100];
  assign o[51398] = i[100];
  assign o[51399] = i[100];
  assign o[51400] = i[100];
  assign o[51401] = i[100];
  assign o[51402] = i[100];
  assign o[51403] = i[100];
  assign o[51404] = i[100];
  assign o[51405] = i[100];
  assign o[51406] = i[100];
  assign o[51407] = i[100];
  assign o[51408] = i[100];
  assign o[51409] = i[100];
  assign o[51410] = i[100];
  assign o[51411] = i[100];
  assign o[51412] = i[100];
  assign o[51413] = i[100];
  assign o[51414] = i[100];
  assign o[51415] = i[100];
  assign o[51416] = i[100];
  assign o[51417] = i[100];
  assign o[51418] = i[100];
  assign o[51419] = i[100];
  assign o[51420] = i[100];
  assign o[51421] = i[100];
  assign o[51422] = i[100];
  assign o[51423] = i[100];
  assign o[51424] = i[100];
  assign o[51425] = i[100];
  assign o[51426] = i[100];
  assign o[51427] = i[100];
  assign o[51428] = i[100];
  assign o[51429] = i[100];
  assign o[51430] = i[100];
  assign o[51431] = i[100];
  assign o[51432] = i[100];
  assign o[51433] = i[100];
  assign o[51434] = i[100];
  assign o[51435] = i[100];
  assign o[51436] = i[100];
  assign o[51437] = i[100];
  assign o[51438] = i[100];
  assign o[51439] = i[100];
  assign o[51440] = i[100];
  assign o[51441] = i[100];
  assign o[51442] = i[100];
  assign o[51443] = i[100];
  assign o[51444] = i[100];
  assign o[51445] = i[100];
  assign o[51446] = i[100];
  assign o[51447] = i[100];
  assign o[51448] = i[100];
  assign o[51449] = i[100];
  assign o[51450] = i[100];
  assign o[51451] = i[100];
  assign o[51452] = i[100];
  assign o[51453] = i[100];
  assign o[51454] = i[100];
  assign o[51455] = i[100];
  assign o[51456] = i[100];
  assign o[51457] = i[100];
  assign o[51458] = i[100];
  assign o[51459] = i[100];
  assign o[51460] = i[100];
  assign o[51461] = i[100];
  assign o[51462] = i[100];
  assign o[51463] = i[100];
  assign o[51464] = i[100];
  assign o[51465] = i[100];
  assign o[51466] = i[100];
  assign o[51467] = i[100];
  assign o[51468] = i[100];
  assign o[51469] = i[100];
  assign o[51470] = i[100];
  assign o[51471] = i[100];
  assign o[51472] = i[100];
  assign o[51473] = i[100];
  assign o[51474] = i[100];
  assign o[51475] = i[100];
  assign o[51476] = i[100];
  assign o[51477] = i[100];
  assign o[51478] = i[100];
  assign o[51479] = i[100];
  assign o[51480] = i[100];
  assign o[51481] = i[100];
  assign o[51482] = i[100];
  assign o[51483] = i[100];
  assign o[51484] = i[100];
  assign o[51485] = i[100];
  assign o[51486] = i[100];
  assign o[51487] = i[100];
  assign o[51488] = i[100];
  assign o[51489] = i[100];
  assign o[51490] = i[100];
  assign o[51491] = i[100];
  assign o[51492] = i[100];
  assign o[51493] = i[100];
  assign o[51494] = i[100];
  assign o[51495] = i[100];
  assign o[51496] = i[100];
  assign o[51497] = i[100];
  assign o[51498] = i[100];
  assign o[51499] = i[100];
  assign o[51500] = i[100];
  assign o[51501] = i[100];
  assign o[51502] = i[100];
  assign o[51503] = i[100];
  assign o[51504] = i[100];
  assign o[51505] = i[100];
  assign o[51506] = i[100];
  assign o[51507] = i[100];
  assign o[51508] = i[100];
  assign o[51509] = i[100];
  assign o[51510] = i[100];
  assign o[51511] = i[100];
  assign o[51512] = i[100];
  assign o[51513] = i[100];
  assign o[51514] = i[100];
  assign o[51515] = i[100];
  assign o[51516] = i[100];
  assign o[51517] = i[100];
  assign o[51518] = i[100];
  assign o[51519] = i[100];
  assign o[51520] = i[100];
  assign o[51521] = i[100];
  assign o[51522] = i[100];
  assign o[51523] = i[100];
  assign o[51524] = i[100];
  assign o[51525] = i[100];
  assign o[51526] = i[100];
  assign o[51527] = i[100];
  assign o[51528] = i[100];
  assign o[51529] = i[100];
  assign o[51530] = i[100];
  assign o[51531] = i[100];
  assign o[51532] = i[100];
  assign o[51533] = i[100];
  assign o[51534] = i[100];
  assign o[51535] = i[100];
  assign o[51536] = i[100];
  assign o[51537] = i[100];
  assign o[51538] = i[100];
  assign o[51539] = i[100];
  assign o[51540] = i[100];
  assign o[51541] = i[100];
  assign o[51542] = i[100];
  assign o[51543] = i[100];
  assign o[51544] = i[100];
  assign o[51545] = i[100];
  assign o[51546] = i[100];
  assign o[51547] = i[100];
  assign o[51548] = i[100];
  assign o[51549] = i[100];
  assign o[51550] = i[100];
  assign o[51551] = i[100];
  assign o[51552] = i[100];
  assign o[51553] = i[100];
  assign o[51554] = i[100];
  assign o[51555] = i[100];
  assign o[51556] = i[100];
  assign o[51557] = i[100];
  assign o[51558] = i[100];
  assign o[51559] = i[100];
  assign o[51560] = i[100];
  assign o[51561] = i[100];
  assign o[51562] = i[100];
  assign o[51563] = i[100];
  assign o[51564] = i[100];
  assign o[51565] = i[100];
  assign o[51566] = i[100];
  assign o[51567] = i[100];
  assign o[51568] = i[100];
  assign o[51569] = i[100];
  assign o[51570] = i[100];
  assign o[51571] = i[100];
  assign o[51572] = i[100];
  assign o[51573] = i[100];
  assign o[51574] = i[100];
  assign o[51575] = i[100];
  assign o[51576] = i[100];
  assign o[51577] = i[100];
  assign o[51578] = i[100];
  assign o[51579] = i[100];
  assign o[51580] = i[100];
  assign o[51581] = i[100];
  assign o[51582] = i[100];
  assign o[51583] = i[100];
  assign o[51584] = i[100];
  assign o[51585] = i[100];
  assign o[51586] = i[100];
  assign o[51587] = i[100];
  assign o[51588] = i[100];
  assign o[51589] = i[100];
  assign o[51590] = i[100];
  assign o[51591] = i[100];
  assign o[51592] = i[100];
  assign o[51593] = i[100];
  assign o[51594] = i[100];
  assign o[51595] = i[100];
  assign o[51596] = i[100];
  assign o[51597] = i[100];
  assign o[51598] = i[100];
  assign o[51599] = i[100];
  assign o[51600] = i[100];
  assign o[51601] = i[100];
  assign o[51602] = i[100];
  assign o[51603] = i[100];
  assign o[51604] = i[100];
  assign o[51605] = i[100];
  assign o[51606] = i[100];
  assign o[51607] = i[100];
  assign o[51608] = i[100];
  assign o[51609] = i[100];
  assign o[51610] = i[100];
  assign o[51611] = i[100];
  assign o[51612] = i[100];
  assign o[51613] = i[100];
  assign o[51614] = i[100];
  assign o[51615] = i[100];
  assign o[51616] = i[100];
  assign o[51617] = i[100];
  assign o[51618] = i[100];
  assign o[51619] = i[100];
  assign o[51620] = i[100];
  assign o[51621] = i[100];
  assign o[51622] = i[100];
  assign o[51623] = i[100];
  assign o[51624] = i[100];
  assign o[51625] = i[100];
  assign o[51626] = i[100];
  assign o[51627] = i[100];
  assign o[51628] = i[100];
  assign o[51629] = i[100];
  assign o[51630] = i[100];
  assign o[51631] = i[100];
  assign o[51632] = i[100];
  assign o[51633] = i[100];
  assign o[51634] = i[100];
  assign o[51635] = i[100];
  assign o[51636] = i[100];
  assign o[51637] = i[100];
  assign o[51638] = i[100];
  assign o[51639] = i[100];
  assign o[51640] = i[100];
  assign o[51641] = i[100];
  assign o[51642] = i[100];
  assign o[51643] = i[100];
  assign o[51644] = i[100];
  assign o[51645] = i[100];
  assign o[51646] = i[100];
  assign o[51647] = i[100];
  assign o[51648] = i[100];
  assign o[51649] = i[100];
  assign o[51650] = i[100];
  assign o[51651] = i[100];
  assign o[51652] = i[100];
  assign o[51653] = i[100];
  assign o[51654] = i[100];
  assign o[51655] = i[100];
  assign o[51656] = i[100];
  assign o[51657] = i[100];
  assign o[51658] = i[100];
  assign o[51659] = i[100];
  assign o[51660] = i[100];
  assign o[51661] = i[100];
  assign o[51662] = i[100];
  assign o[51663] = i[100];
  assign o[51664] = i[100];
  assign o[51665] = i[100];
  assign o[51666] = i[100];
  assign o[51667] = i[100];
  assign o[51668] = i[100];
  assign o[51669] = i[100];
  assign o[51670] = i[100];
  assign o[51671] = i[100];
  assign o[51672] = i[100];
  assign o[51673] = i[100];
  assign o[51674] = i[100];
  assign o[51675] = i[100];
  assign o[51676] = i[100];
  assign o[51677] = i[100];
  assign o[51678] = i[100];
  assign o[51679] = i[100];
  assign o[51680] = i[100];
  assign o[51681] = i[100];
  assign o[51682] = i[100];
  assign o[51683] = i[100];
  assign o[51684] = i[100];
  assign o[51685] = i[100];
  assign o[51686] = i[100];
  assign o[51687] = i[100];
  assign o[51688] = i[100];
  assign o[51689] = i[100];
  assign o[51690] = i[100];
  assign o[51691] = i[100];
  assign o[51692] = i[100];
  assign o[51693] = i[100];
  assign o[51694] = i[100];
  assign o[51695] = i[100];
  assign o[51696] = i[100];
  assign o[51697] = i[100];
  assign o[51698] = i[100];
  assign o[51699] = i[100];
  assign o[51700] = i[100];
  assign o[51701] = i[100];
  assign o[51702] = i[100];
  assign o[51703] = i[100];
  assign o[51704] = i[100];
  assign o[51705] = i[100];
  assign o[51706] = i[100];
  assign o[51707] = i[100];
  assign o[51708] = i[100];
  assign o[51709] = i[100];
  assign o[51710] = i[100];
  assign o[51711] = i[100];
  assign o[50688] = i[99];
  assign o[50689] = i[99];
  assign o[50690] = i[99];
  assign o[50691] = i[99];
  assign o[50692] = i[99];
  assign o[50693] = i[99];
  assign o[50694] = i[99];
  assign o[50695] = i[99];
  assign o[50696] = i[99];
  assign o[50697] = i[99];
  assign o[50698] = i[99];
  assign o[50699] = i[99];
  assign o[50700] = i[99];
  assign o[50701] = i[99];
  assign o[50702] = i[99];
  assign o[50703] = i[99];
  assign o[50704] = i[99];
  assign o[50705] = i[99];
  assign o[50706] = i[99];
  assign o[50707] = i[99];
  assign o[50708] = i[99];
  assign o[50709] = i[99];
  assign o[50710] = i[99];
  assign o[50711] = i[99];
  assign o[50712] = i[99];
  assign o[50713] = i[99];
  assign o[50714] = i[99];
  assign o[50715] = i[99];
  assign o[50716] = i[99];
  assign o[50717] = i[99];
  assign o[50718] = i[99];
  assign o[50719] = i[99];
  assign o[50720] = i[99];
  assign o[50721] = i[99];
  assign o[50722] = i[99];
  assign o[50723] = i[99];
  assign o[50724] = i[99];
  assign o[50725] = i[99];
  assign o[50726] = i[99];
  assign o[50727] = i[99];
  assign o[50728] = i[99];
  assign o[50729] = i[99];
  assign o[50730] = i[99];
  assign o[50731] = i[99];
  assign o[50732] = i[99];
  assign o[50733] = i[99];
  assign o[50734] = i[99];
  assign o[50735] = i[99];
  assign o[50736] = i[99];
  assign o[50737] = i[99];
  assign o[50738] = i[99];
  assign o[50739] = i[99];
  assign o[50740] = i[99];
  assign o[50741] = i[99];
  assign o[50742] = i[99];
  assign o[50743] = i[99];
  assign o[50744] = i[99];
  assign o[50745] = i[99];
  assign o[50746] = i[99];
  assign o[50747] = i[99];
  assign o[50748] = i[99];
  assign o[50749] = i[99];
  assign o[50750] = i[99];
  assign o[50751] = i[99];
  assign o[50752] = i[99];
  assign o[50753] = i[99];
  assign o[50754] = i[99];
  assign o[50755] = i[99];
  assign o[50756] = i[99];
  assign o[50757] = i[99];
  assign o[50758] = i[99];
  assign o[50759] = i[99];
  assign o[50760] = i[99];
  assign o[50761] = i[99];
  assign o[50762] = i[99];
  assign o[50763] = i[99];
  assign o[50764] = i[99];
  assign o[50765] = i[99];
  assign o[50766] = i[99];
  assign o[50767] = i[99];
  assign o[50768] = i[99];
  assign o[50769] = i[99];
  assign o[50770] = i[99];
  assign o[50771] = i[99];
  assign o[50772] = i[99];
  assign o[50773] = i[99];
  assign o[50774] = i[99];
  assign o[50775] = i[99];
  assign o[50776] = i[99];
  assign o[50777] = i[99];
  assign o[50778] = i[99];
  assign o[50779] = i[99];
  assign o[50780] = i[99];
  assign o[50781] = i[99];
  assign o[50782] = i[99];
  assign o[50783] = i[99];
  assign o[50784] = i[99];
  assign o[50785] = i[99];
  assign o[50786] = i[99];
  assign o[50787] = i[99];
  assign o[50788] = i[99];
  assign o[50789] = i[99];
  assign o[50790] = i[99];
  assign o[50791] = i[99];
  assign o[50792] = i[99];
  assign o[50793] = i[99];
  assign o[50794] = i[99];
  assign o[50795] = i[99];
  assign o[50796] = i[99];
  assign o[50797] = i[99];
  assign o[50798] = i[99];
  assign o[50799] = i[99];
  assign o[50800] = i[99];
  assign o[50801] = i[99];
  assign o[50802] = i[99];
  assign o[50803] = i[99];
  assign o[50804] = i[99];
  assign o[50805] = i[99];
  assign o[50806] = i[99];
  assign o[50807] = i[99];
  assign o[50808] = i[99];
  assign o[50809] = i[99];
  assign o[50810] = i[99];
  assign o[50811] = i[99];
  assign o[50812] = i[99];
  assign o[50813] = i[99];
  assign o[50814] = i[99];
  assign o[50815] = i[99];
  assign o[50816] = i[99];
  assign o[50817] = i[99];
  assign o[50818] = i[99];
  assign o[50819] = i[99];
  assign o[50820] = i[99];
  assign o[50821] = i[99];
  assign o[50822] = i[99];
  assign o[50823] = i[99];
  assign o[50824] = i[99];
  assign o[50825] = i[99];
  assign o[50826] = i[99];
  assign o[50827] = i[99];
  assign o[50828] = i[99];
  assign o[50829] = i[99];
  assign o[50830] = i[99];
  assign o[50831] = i[99];
  assign o[50832] = i[99];
  assign o[50833] = i[99];
  assign o[50834] = i[99];
  assign o[50835] = i[99];
  assign o[50836] = i[99];
  assign o[50837] = i[99];
  assign o[50838] = i[99];
  assign o[50839] = i[99];
  assign o[50840] = i[99];
  assign o[50841] = i[99];
  assign o[50842] = i[99];
  assign o[50843] = i[99];
  assign o[50844] = i[99];
  assign o[50845] = i[99];
  assign o[50846] = i[99];
  assign o[50847] = i[99];
  assign o[50848] = i[99];
  assign o[50849] = i[99];
  assign o[50850] = i[99];
  assign o[50851] = i[99];
  assign o[50852] = i[99];
  assign o[50853] = i[99];
  assign o[50854] = i[99];
  assign o[50855] = i[99];
  assign o[50856] = i[99];
  assign o[50857] = i[99];
  assign o[50858] = i[99];
  assign o[50859] = i[99];
  assign o[50860] = i[99];
  assign o[50861] = i[99];
  assign o[50862] = i[99];
  assign o[50863] = i[99];
  assign o[50864] = i[99];
  assign o[50865] = i[99];
  assign o[50866] = i[99];
  assign o[50867] = i[99];
  assign o[50868] = i[99];
  assign o[50869] = i[99];
  assign o[50870] = i[99];
  assign o[50871] = i[99];
  assign o[50872] = i[99];
  assign o[50873] = i[99];
  assign o[50874] = i[99];
  assign o[50875] = i[99];
  assign o[50876] = i[99];
  assign o[50877] = i[99];
  assign o[50878] = i[99];
  assign o[50879] = i[99];
  assign o[50880] = i[99];
  assign o[50881] = i[99];
  assign o[50882] = i[99];
  assign o[50883] = i[99];
  assign o[50884] = i[99];
  assign o[50885] = i[99];
  assign o[50886] = i[99];
  assign o[50887] = i[99];
  assign o[50888] = i[99];
  assign o[50889] = i[99];
  assign o[50890] = i[99];
  assign o[50891] = i[99];
  assign o[50892] = i[99];
  assign o[50893] = i[99];
  assign o[50894] = i[99];
  assign o[50895] = i[99];
  assign o[50896] = i[99];
  assign o[50897] = i[99];
  assign o[50898] = i[99];
  assign o[50899] = i[99];
  assign o[50900] = i[99];
  assign o[50901] = i[99];
  assign o[50902] = i[99];
  assign o[50903] = i[99];
  assign o[50904] = i[99];
  assign o[50905] = i[99];
  assign o[50906] = i[99];
  assign o[50907] = i[99];
  assign o[50908] = i[99];
  assign o[50909] = i[99];
  assign o[50910] = i[99];
  assign o[50911] = i[99];
  assign o[50912] = i[99];
  assign o[50913] = i[99];
  assign o[50914] = i[99];
  assign o[50915] = i[99];
  assign o[50916] = i[99];
  assign o[50917] = i[99];
  assign o[50918] = i[99];
  assign o[50919] = i[99];
  assign o[50920] = i[99];
  assign o[50921] = i[99];
  assign o[50922] = i[99];
  assign o[50923] = i[99];
  assign o[50924] = i[99];
  assign o[50925] = i[99];
  assign o[50926] = i[99];
  assign o[50927] = i[99];
  assign o[50928] = i[99];
  assign o[50929] = i[99];
  assign o[50930] = i[99];
  assign o[50931] = i[99];
  assign o[50932] = i[99];
  assign o[50933] = i[99];
  assign o[50934] = i[99];
  assign o[50935] = i[99];
  assign o[50936] = i[99];
  assign o[50937] = i[99];
  assign o[50938] = i[99];
  assign o[50939] = i[99];
  assign o[50940] = i[99];
  assign o[50941] = i[99];
  assign o[50942] = i[99];
  assign o[50943] = i[99];
  assign o[50944] = i[99];
  assign o[50945] = i[99];
  assign o[50946] = i[99];
  assign o[50947] = i[99];
  assign o[50948] = i[99];
  assign o[50949] = i[99];
  assign o[50950] = i[99];
  assign o[50951] = i[99];
  assign o[50952] = i[99];
  assign o[50953] = i[99];
  assign o[50954] = i[99];
  assign o[50955] = i[99];
  assign o[50956] = i[99];
  assign o[50957] = i[99];
  assign o[50958] = i[99];
  assign o[50959] = i[99];
  assign o[50960] = i[99];
  assign o[50961] = i[99];
  assign o[50962] = i[99];
  assign o[50963] = i[99];
  assign o[50964] = i[99];
  assign o[50965] = i[99];
  assign o[50966] = i[99];
  assign o[50967] = i[99];
  assign o[50968] = i[99];
  assign o[50969] = i[99];
  assign o[50970] = i[99];
  assign o[50971] = i[99];
  assign o[50972] = i[99];
  assign o[50973] = i[99];
  assign o[50974] = i[99];
  assign o[50975] = i[99];
  assign o[50976] = i[99];
  assign o[50977] = i[99];
  assign o[50978] = i[99];
  assign o[50979] = i[99];
  assign o[50980] = i[99];
  assign o[50981] = i[99];
  assign o[50982] = i[99];
  assign o[50983] = i[99];
  assign o[50984] = i[99];
  assign o[50985] = i[99];
  assign o[50986] = i[99];
  assign o[50987] = i[99];
  assign o[50988] = i[99];
  assign o[50989] = i[99];
  assign o[50990] = i[99];
  assign o[50991] = i[99];
  assign o[50992] = i[99];
  assign o[50993] = i[99];
  assign o[50994] = i[99];
  assign o[50995] = i[99];
  assign o[50996] = i[99];
  assign o[50997] = i[99];
  assign o[50998] = i[99];
  assign o[50999] = i[99];
  assign o[51000] = i[99];
  assign o[51001] = i[99];
  assign o[51002] = i[99];
  assign o[51003] = i[99];
  assign o[51004] = i[99];
  assign o[51005] = i[99];
  assign o[51006] = i[99];
  assign o[51007] = i[99];
  assign o[51008] = i[99];
  assign o[51009] = i[99];
  assign o[51010] = i[99];
  assign o[51011] = i[99];
  assign o[51012] = i[99];
  assign o[51013] = i[99];
  assign o[51014] = i[99];
  assign o[51015] = i[99];
  assign o[51016] = i[99];
  assign o[51017] = i[99];
  assign o[51018] = i[99];
  assign o[51019] = i[99];
  assign o[51020] = i[99];
  assign o[51021] = i[99];
  assign o[51022] = i[99];
  assign o[51023] = i[99];
  assign o[51024] = i[99];
  assign o[51025] = i[99];
  assign o[51026] = i[99];
  assign o[51027] = i[99];
  assign o[51028] = i[99];
  assign o[51029] = i[99];
  assign o[51030] = i[99];
  assign o[51031] = i[99];
  assign o[51032] = i[99];
  assign o[51033] = i[99];
  assign o[51034] = i[99];
  assign o[51035] = i[99];
  assign o[51036] = i[99];
  assign o[51037] = i[99];
  assign o[51038] = i[99];
  assign o[51039] = i[99];
  assign o[51040] = i[99];
  assign o[51041] = i[99];
  assign o[51042] = i[99];
  assign o[51043] = i[99];
  assign o[51044] = i[99];
  assign o[51045] = i[99];
  assign o[51046] = i[99];
  assign o[51047] = i[99];
  assign o[51048] = i[99];
  assign o[51049] = i[99];
  assign o[51050] = i[99];
  assign o[51051] = i[99];
  assign o[51052] = i[99];
  assign o[51053] = i[99];
  assign o[51054] = i[99];
  assign o[51055] = i[99];
  assign o[51056] = i[99];
  assign o[51057] = i[99];
  assign o[51058] = i[99];
  assign o[51059] = i[99];
  assign o[51060] = i[99];
  assign o[51061] = i[99];
  assign o[51062] = i[99];
  assign o[51063] = i[99];
  assign o[51064] = i[99];
  assign o[51065] = i[99];
  assign o[51066] = i[99];
  assign o[51067] = i[99];
  assign o[51068] = i[99];
  assign o[51069] = i[99];
  assign o[51070] = i[99];
  assign o[51071] = i[99];
  assign o[51072] = i[99];
  assign o[51073] = i[99];
  assign o[51074] = i[99];
  assign o[51075] = i[99];
  assign o[51076] = i[99];
  assign o[51077] = i[99];
  assign o[51078] = i[99];
  assign o[51079] = i[99];
  assign o[51080] = i[99];
  assign o[51081] = i[99];
  assign o[51082] = i[99];
  assign o[51083] = i[99];
  assign o[51084] = i[99];
  assign o[51085] = i[99];
  assign o[51086] = i[99];
  assign o[51087] = i[99];
  assign o[51088] = i[99];
  assign o[51089] = i[99];
  assign o[51090] = i[99];
  assign o[51091] = i[99];
  assign o[51092] = i[99];
  assign o[51093] = i[99];
  assign o[51094] = i[99];
  assign o[51095] = i[99];
  assign o[51096] = i[99];
  assign o[51097] = i[99];
  assign o[51098] = i[99];
  assign o[51099] = i[99];
  assign o[51100] = i[99];
  assign o[51101] = i[99];
  assign o[51102] = i[99];
  assign o[51103] = i[99];
  assign o[51104] = i[99];
  assign o[51105] = i[99];
  assign o[51106] = i[99];
  assign o[51107] = i[99];
  assign o[51108] = i[99];
  assign o[51109] = i[99];
  assign o[51110] = i[99];
  assign o[51111] = i[99];
  assign o[51112] = i[99];
  assign o[51113] = i[99];
  assign o[51114] = i[99];
  assign o[51115] = i[99];
  assign o[51116] = i[99];
  assign o[51117] = i[99];
  assign o[51118] = i[99];
  assign o[51119] = i[99];
  assign o[51120] = i[99];
  assign o[51121] = i[99];
  assign o[51122] = i[99];
  assign o[51123] = i[99];
  assign o[51124] = i[99];
  assign o[51125] = i[99];
  assign o[51126] = i[99];
  assign o[51127] = i[99];
  assign o[51128] = i[99];
  assign o[51129] = i[99];
  assign o[51130] = i[99];
  assign o[51131] = i[99];
  assign o[51132] = i[99];
  assign o[51133] = i[99];
  assign o[51134] = i[99];
  assign o[51135] = i[99];
  assign o[51136] = i[99];
  assign o[51137] = i[99];
  assign o[51138] = i[99];
  assign o[51139] = i[99];
  assign o[51140] = i[99];
  assign o[51141] = i[99];
  assign o[51142] = i[99];
  assign o[51143] = i[99];
  assign o[51144] = i[99];
  assign o[51145] = i[99];
  assign o[51146] = i[99];
  assign o[51147] = i[99];
  assign o[51148] = i[99];
  assign o[51149] = i[99];
  assign o[51150] = i[99];
  assign o[51151] = i[99];
  assign o[51152] = i[99];
  assign o[51153] = i[99];
  assign o[51154] = i[99];
  assign o[51155] = i[99];
  assign o[51156] = i[99];
  assign o[51157] = i[99];
  assign o[51158] = i[99];
  assign o[51159] = i[99];
  assign o[51160] = i[99];
  assign o[51161] = i[99];
  assign o[51162] = i[99];
  assign o[51163] = i[99];
  assign o[51164] = i[99];
  assign o[51165] = i[99];
  assign o[51166] = i[99];
  assign o[51167] = i[99];
  assign o[51168] = i[99];
  assign o[51169] = i[99];
  assign o[51170] = i[99];
  assign o[51171] = i[99];
  assign o[51172] = i[99];
  assign o[51173] = i[99];
  assign o[51174] = i[99];
  assign o[51175] = i[99];
  assign o[51176] = i[99];
  assign o[51177] = i[99];
  assign o[51178] = i[99];
  assign o[51179] = i[99];
  assign o[51180] = i[99];
  assign o[51181] = i[99];
  assign o[51182] = i[99];
  assign o[51183] = i[99];
  assign o[51184] = i[99];
  assign o[51185] = i[99];
  assign o[51186] = i[99];
  assign o[51187] = i[99];
  assign o[51188] = i[99];
  assign o[51189] = i[99];
  assign o[51190] = i[99];
  assign o[51191] = i[99];
  assign o[51192] = i[99];
  assign o[51193] = i[99];
  assign o[51194] = i[99];
  assign o[51195] = i[99];
  assign o[51196] = i[99];
  assign o[51197] = i[99];
  assign o[51198] = i[99];
  assign o[51199] = i[99];
  assign o[50176] = i[98];
  assign o[50177] = i[98];
  assign o[50178] = i[98];
  assign o[50179] = i[98];
  assign o[50180] = i[98];
  assign o[50181] = i[98];
  assign o[50182] = i[98];
  assign o[50183] = i[98];
  assign o[50184] = i[98];
  assign o[50185] = i[98];
  assign o[50186] = i[98];
  assign o[50187] = i[98];
  assign o[50188] = i[98];
  assign o[50189] = i[98];
  assign o[50190] = i[98];
  assign o[50191] = i[98];
  assign o[50192] = i[98];
  assign o[50193] = i[98];
  assign o[50194] = i[98];
  assign o[50195] = i[98];
  assign o[50196] = i[98];
  assign o[50197] = i[98];
  assign o[50198] = i[98];
  assign o[50199] = i[98];
  assign o[50200] = i[98];
  assign o[50201] = i[98];
  assign o[50202] = i[98];
  assign o[50203] = i[98];
  assign o[50204] = i[98];
  assign o[50205] = i[98];
  assign o[50206] = i[98];
  assign o[50207] = i[98];
  assign o[50208] = i[98];
  assign o[50209] = i[98];
  assign o[50210] = i[98];
  assign o[50211] = i[98];
  assign o[50212] = i[98];
  assign o[50213] = i[98];
  assign o[50214] = i[98];
  assign o[50215] = i[98];
  assign o[50216] = i[98];
  assign o[50217] = i[98];
  assign o[50218] = i[98];
  assign o[50219] = i[98];
  assign o[50220] = i[98];
  assign o[50221] = i[98];
  assign o[50222] = i[98];
  assign o[50223] = i[98];
  assign o[50224] = i[98];
  assign o[50225] = i[98];
  assign o[50226] = i[98];
  assign o[50227] = i[98];
  assign o[50228] = i[98];
  assign o[50229] = i[98];
  assign o[50230] = i[98];
  assign o[50231] = i[98];
  assign o[50232] = i[98];
  assign o[50233] = i[98];
  assign o[50234] = i[98];
  assign o[50235] = i[98];
  assign o[50236] = i[98];
  assign o[50237] = i[98];
  assign o[50238] = i[98];
  assign o[50239] = i[98];
  assign o[50240] = i[98];
  assign o[50241] = i[98];
  assign o[50242] = i[98];
  assign o[50243] = i[98];
  assign o[50244] = i[98];
  assign o[50245] = i[98];
  assign o[50246] = i[98];
  assign o[50247] = i[98];
  assign o[50248] = i[98];
  assign o[50249] = i[98];
  assign o[50250] = i[98];
  assign o[50251] = i[98];
  assign o[50252] = i[98];
  assign o[50253] = i[98];
  assign o[50254] = i[98];
  assign o[50255] = i[98];
  assign o[50256] = i[98];
  assign o[50257] = i[98];
  assign o[50258] = i[98];
  assign o[50259] = i[98];
  assign o[50260] = i[98];
  assign o[50261] = i[98];
  assign o[50262] = i[98];
  assign o[50263] = i[98];
  assign o[50264] = i[98];
  assign o[50265] = i[98];
  assign o[50266] = i[98];
  assign o[50267] = i[98];
  assign o[50268] = i[98];
  assign o[50269] = i[98];
  assign o[50270] = i[98];
  assign o[50271] = i[98];
  assign o[50272] = i[98];
  assign o[50273] = i[98];
  assign o[50274] = i[98];
  assign o[50275] = i[98];
  assign o[50276] = i[98];
  assign o[50277] = i[98];
  assign o[50278] = i[98];
  assign o[50279] = i[98];
  assign o[50280] = i[98];
  assign o[50281] = i[98];
  assign o[50282] = i[98];
  assign o[50283] = i[98];
  assign o[50284] = i[98];
  assign o[50285] = i[98];
  assign o[50286] = i[98];
  assign o[50287] = i[98];
  assign o[50288] = i[98];
  assign o[50289] = i[98];
  assign o[50290] = i[98];
  assign o[50291] = i[98];
  assign o[50292] = i[98];
  assign o[50293] = i[98];
  assign o[50294] = i[98];
  assign o[50295] = i[98];
  assign o[50296] = i[98];
  assign o[50297] = i[98];
  assign o[50298] = i[98];
  assign o[50299] = i[98];
  assign o[50300] = i[98];
  assign o[50301] = i[98];
  assign o[50302] = i[98];
  assign o[50303] = i[98];
  assign o[50304] = i[98];
  assign o[50305] = i[98];
  assign o[50306] = i[98];
  assign o[50307] = i[98];
  assign o[50308] = i[98];
  assign o[50309] = i[98];
  assign o[50310] = i[98];
  assign o[50311] = i[98];
  assign o[50312] = i[98];
  assign o[50313] = i[98];
  assign o[50314] = i[98];
  assign o[50315] = i[98];
  assign o[50316] = i[98];
  assign o[50317] = i[98];
  assign o[50318] = i[98];
  assign o[50319] = i[98];
  assign o[50320] = i[98];
  assign o[50321] = i[98];
  assign o[50322] = i[98];
  assign o[50323] = i[98];
  assign o[50324] = i[98];
  assign o[50325] = i[98];
  assign o[50326] = i[98];
  assign o[50327] = i[98];
  assign o[50328] = i[98];
  assign o[50329] = i[98];
  assign o[50330] = i[98];
  assign o[50331] = i[98];
  assign o[50332] = i[98];
  assign o[50333] = i[98];
  assign o[50334] = i[98];
  assign o[50335] = i[98];
  assign o[50336] = i[98];
  assign o[50337] = i[98];
  assign o[50338] = i[98];
  assign o[50339] = i[98];
  assign o[50340] = i[98];
  assign o[50341] = i[98];
  assign o[50342] = i[98];
  assign o[50343] = i[98];
  assign o[50344] = i[98];
  assign o[50345] = i[98];
  assign o[50346] = i[98];
  assign o[50347] = i[98];
  assign o[50348] = i[98];
  assign o[50349] = i[98];
  assign o[50350] = i[98];
  assign o[50351] = i[98];
  assign o[50352] = i[98];
  assign o[50353] = i[98];
  assign o[50354] = i[98];
  assign o[50355] = i[98];
  assign o[50356] = i[98];
  assign o[50357] = i[98];
  assign o[50358] = i[98];
  assign o[50359] = i[98];
  assign o[50360] = i[98];
  assign o[50361] = i[98];
  assign o[50362] = i[98];
  assign o[50363] = i[98];
  assign o[50364] = i[98];
  assign o[50365] = i[98];
  assign o[50366] = i[98];
  assign o[50367] = i[98];
  assign o[50368] = i[98];
  assign o[50369] = i[98];
  assign o[50370] = i[98];
  assign o[50371] = i[98];
  assign o[50372] = i[98];
  assign o[50373] = i[98];
  assign o[50374] = i[98];
  assign o[50375] = i[98];
  assign o[50376] = i[98];
  assign o[50377] = i[98];
  assign o[50378] = i[98];
  assign o[50379] = i[98];
  assign o[50380] = i[98];
  assign o[50381] = i[98];
  assign o[50382] = i[98];
  assign o[50383] = i[98];
  assign o[50384] = i[98];
  assign o[50385] = i[98];
  assign o[50386] = i[98];
  assign o[50387] = i[98];
  assign o[50388] = i[98];
  assign o[50389] = i[98];
  assign o[50390] = i[98];
  assign o[50391] = i[98];
  assign o[50392] = i[98];
  assign o[50393] = i[98];
  assign o[50394] = i[98];
  assign o[50395] = i[98];
  assign o[50396] = i[98];
  assign o[50397] = i[98];
  assign o[50398] = i[98];
  assign o[50399] = i[98];
  assign o[50400] = i[98];
  assign o[50401] = i[98];
  assign o[50402] = i[98];
  assign o[50403] = i[98];
  assign o[50404] = i[98];
  assign o[50405] = i[98];
  assign o[50406] = i[98];
  assign o[50407] = i[98];
  assign o[50408] = i[98];
  assign o[50409] = i[98];
  assign o[50410] = i[98];
  assign o[50411] = i[98];
  assign o[50412] = i[98];
  assign o[50413] = i[98];
  assign o[50414] = i[98];
  assign o[50415] = i[98];
  assign o[50416] = i[98];
  assign o[50417] = i[98];
  assign o[50418] = i[98];
  assign o[50419] = i[98];
  assign o[50420] = i[98];
  assign o[50421] = i[98];
  assign o[50422] = i[98];
  assign o[50423] = i[98];
  assign o[50424] = i[98];
  assign o[50425] = i[98];
  assign o[50426] = i[98];
  assign o[50427] = i[98];
  assign o[50428] = i[98];
  assign o[50429] = i[98];
  assign o[50430] = i[98];
  assign o[50431] = i[98];
  assign o[50432] = i[98];
  assign o[50433] = i[98];
  assign o[50434] = i[98];
  assign o[50435] = i[98];
  assign o[50436] = i[98];
  assign o[50437] = i[98];
  assign o[50438] = i[98];
  assign o[50439] = i[98];
  assign o[50440] = i[98];
  assign o[50441] = i[98];
  assign o[50442] = i[98];
  assign o[50443] = i[98];
  assign o[50444] = i[98];
  assign o[50445] = i[98];
  assign o[50446] = i[98];
  assign o[50447] = i[98];
  assign o[50448] = i[98];
  assign o[50449] = i[98];
  assign o[50450] = i[98];
  assign o[50451] = i[98];
  assign o[50452] = i[98];
  assign o[50453] = i[98];
  assign o[50454] = i[98];
  assign o[50455] = i[98];
  assign o[50456] = i[98];
  assign o[50457] = i[98];
  assign o[50458] = i[98];
  assign o[50459] = i[98];
  assign o[50460] = i[98];
  assign o[50461] = i[98];
  assign o[50462] = i[98];
  assign o[50463] = i[98];
  assign o[50464] = i[98];
  assign o[50465] = i[98];
  assign o[50466] = i[98];
  assign o[50467] = i[98];
  assign o[50468] = i[98];
  assign o[50469] = i[98];
  assign o[50470] = i[98];
  assign o[50471] = i[98];
  assign o[50472] = i[98];
  assign o[50473] = i[98];
  assign o[50474] = i[98];
  assign o[50475] = i[98];
  assign o[50476] = i[98];
  assign o[50477] = i[98];
  assign o[50478] = i[98];
  assign o[50479] = i[98];
  assign o[50480] = i[98];
  assign o[50481] = i[98];
  assign o[50482] = i[98];
  assign o[50483] = i[98];
  assign o[50484] = i[98];
  assign o[50485] = i[98];
  assign o[50486] = i[98];
  assign o[50487] = i[98];
  assign o[50488] = i[98];
  assign o[50489] = i[98];
  assign o[50490] = i[98];
  assign o[50491] = i[98];
  assign o[50492] = i[98];
  assign o[50493] = i[98];
  assign o[50494] = i[98];
  assign o[50495] = i[98];
  assign o[50496] = i[98];
  assign o[50497] = i[98];
  assign o[50498] = i[98];
  assign o[50499] = i[98];
  assign o[50500] = i[98];
  assign o[50501] = i[98];
  assign o[50502] = i[98];
  assign o[50503] = i[98];
  assign o[50504] = i[98];
  assign o[50505] = i[98];
  assign o[50506] = i[98];
  assign o[50507] = i[98];
  assign o[50508] = i[98];
  assign o[50509] = i[98];
  assign o[50510] = i[98];
  assign o[50511] = i[98];
  assign o[50512] = i[98];
  assign o[50513] = i[98];
  assign o[50514] = i[98];
  assign o[50515] = i[98];
  assign o[50516] = i[98];
  assign o[50517] = i[98];
  assign o[50518] = i[98];
  assign o[50519] = i[98];
  assign o[50520] = i[98];
  assign o[50521] = i[98];
  assign o[50522] = i[98];
  assign o[50523] = i[98];
  assign o[50524] = i[98];
  assign o[50525] = i[98];
  assign o[50526] = i[98];
  assign o[50527] = i[98];
  assign o[50528] = i[98];
  assign o[50529] = i[98];
  assign o[50530] = i[98];
  assign o[50531] = i[98];
  assign o[50532] = i[98];
  assign o[50533] = i[98];
  assign o[50534] = i[98];
  assign o[50535] = i[98];
  assign o[50536] = i[98];
  assign o[50537] = i[98];
  assign o[50538] = i[98];
  assign o[50539] = i[98];
  assign o[50540] = i[98];
  assign o[50541] = i[98];
  assign o[50542] = i[98];
  assign o[50543] = i[98];
  assign o[50544] = i[98];
  assign o[50545] = i[98];
  assign o[50546] = i[98];
  assign o[50547] = i[98];
  assign o[50548] = i[98];
  assign o[50549] = i[98];
  assign o[50550] = i[98];
  assign o[50551] = i[98];
  assign o[50552] = i[98];
  assign o[50553] = i[98];
  assign o[50554] = i[98];
  assign o[50555] = i[98];
  assign o[50556] = i[98];
  assign o[50557] = i[98];
  assign o[50558] = i[98];
  assign o[50559] = i[98];
  assign o[50560] = i[98];
  assign o[50561] = i[98];
  assign o[50562] = i[98];
  assign o[50563] = i[98];
  assign o[50564] = i[98];
  assign o[50565] = i[98];
  assign o[50566] = i[98];
  assign o[50567] = i[98];
  assign o[50568] = i[98];
  assign o[50569] = i[98];
  assign o[50570] = i[98];
  assign o[50571] = i[98];
  assign o[50572] = i[98];
  assign o[50573] = i[98];
  assign o[50574] = i[98];
  assign o[50575] = i[98];
  assign o[50576] = i[98];
  assign o[50577] = i[98];
  assign o[50578] = i[98];
  assign o[50579] = i[98];
  assign o[50580] = i[98];
  assign o[50581] = i[98];
  assign o[50582] = i[98];
  assign o[50583] = i[98];
  assign o[50584] = i[98];
  assign o[50585] = i[98];
  assign o[50586] = i[98];
  assign o[50587] = i[98];
  assign o[50588] = i[98];
  assign o[50589] = i[98];
  assign o[50590] = i[98];
  assign o[50591] = i[98];
  assign o[50592] = i[98];
  assign o[50593] = i[98];
  assign o[50594] = i[98];
  assign o[50595] = i[98];
  assign o[50596] = i[98];
  assign o[50597] = i[98];
  assign o[50598] = i[98];
  assign o[50599] = i[98];
  assign o[50600] = i[98];
  assign o[50601] = i[98];
  assign o[50602] = i[98];
  assign o[50603] = i[98];
  assign o[50604] = i[98];
  assign o[50605] = i[98];
  assign o[50606] = i[98];
  assign o[50607] = i[98];
  assign o[50608] = i[98];
  assign o[50609] = i[98];
  assign o[50610] = i[98];
  assign o[50611] = i[98];
  assign o[50612] = i[98];
  assign o[50613] = i[98];
  assign o[50614] = i[98];
  assign o[50615] = i[98];
  assign o[50616] = i[98];
  assign o[50617] = i[98];
  assign o[50618] = i[98];
  assign o[50619] = i[98];
  assign o[50620] = i[98];
  assign o[50621] = i[98];
  assign o[50622] = i[98];
  assign o[50623] = i[98];
  assign o[50624] = i[98];
  assign o[50625] = i[98];
  assign o[50626] = i[98];
  assign o[50627] = i[98];
  assign o[50628] = i[98];
  assign o[50629] = i[98];
  assign o[50630] = i[98];
  assign o[50631] = i[98];
  assign o[50632] = i[98];
  assign o[50633] = i[98];
  assign o[50634] = i[98];
  assign o[50635] = i[98];
  assign o[50636] = i[98];
  assign o[50637] = i[98];
  assign o[50638] = i[98];
  assign o[50639] = i[98];
  assign o[50640] = i[98];
  assign o[50641] = i[98];
  assign o[50642] = i[98];
  assign o[50643] = i[98];
  assign o[50644] = i[98];
  assign o[50645] = i[98];
  assign o[50646] = i[98];
  assign o[50647] = i[98];
  assign o[50648] = i[98];
  assign o[50649] = i[98];
  assign o[50650] = i[98];
  assign o[50651] = i[98];
  assign o[50652] = i[98];
  assign o[50653] = i[98];
  assign o[50654] = i[98];
  assign o[50655] = i[98];
  assign o[50656] = i[98];
  assign o[50657] = i[98];
  assign o[50658] = i[98];
  assign o[50659] = i[98];
  assign o[50660] = i[98];
  assign o[50661] = i[98];
  assign o[50662] = i[98];
  assign o[50663] = i[98];
  assign o[50664] = i[98];
  assign o[50665] = i[98];
  assign o[50666] = i[98];
  assign o[50667] = i[98];
  assign o[50668] = i[98];
  assign o[50669] = i[98];
  assign o[50670] = i[98];
  assign o[50671] = i[98];
  assign o[50672] = i[98];
  assign o[50673] = i[98];
  assign o[50674] = i[98];
  assign o[50675] = i[98];
  assign o[50676] = i[98];
  assign o[50677] = i[98];
  assign o[50678] = i[98];
  assign o[50679] = i[98];
  assign o[50680] = i[98];
  assign o[50681] = i[98];
  assign o[50682] = i[98];
  assign o[50683] = i[98];
  assign o[50684] = i[98];
  assign o[50685] = i[98];
  assign o[50686] = i[98];
  assign o[50687] = i[98];
  assign o[49664] = i[97];
  assign o[49665] = i[97];
  assign o[49666] = i[97];
  assign o[49667] = i[97];
  assign o[49668] = i[97];
  assign o[49669] = i[97];
  assign o[49670] = i[97];
  assign o[49671] = i[97];
  assign o[49672] = i[97];
  assign o[49673] = i[97];
  assign o[49674] = i[97];
  assign o[49675] = i[97];
  assign o[49676] = i[97];
  assign o[49677] = i[97];
  assign o[49678] = i[97];
  assign o[49679] = i[97];
  assign o[49680] = i[97];
  assign o[49681] = i[97];
  assign o[49682] = i[97];
  assign o[49683] = i[97];
  assign o[49684] = i[97];
  assign o[49685] = i[97];
  assign o[49686] = i[97];
  assign o[49687] = i[97];
  assign o[49688] = i[97];
  assign o[49689] = i[97];
  assign o[49690] = i[97];
  assign o[49691] = i[97];
  assign o[49692] = i[97];
  assign o[49693] = i[97];
  assign o[49694] = i[97];
  assign o[49695] = i[97];
  assign o[49696] = i[97];
  assign o[49697] = i[97];
  assign o[49698] = i[97];
  assign o[49699] = i[97];
  assign o[49700] = i[97];
  assign o[49701] = i[97];
  assign o[49702] = i[97];
  assign o[49703] = i[97];
  assign o[49704] = i[97];
  assign o[49705] = i[97];
  assign o[49706] = i[97];
  assign o[49707] = i[97];
  assign o[49708] = i[97];
  assign o[49709] = i[97];
  assign o[49710] = i[97];
  assign o[49711] = i[97];
  assign o[49712] = i[97];
  assign o[49713] = i[97];
  assign o[49714] = i[97];
  assign o[49715] = i[97];
  assign o[49716] = i[97];
  assign o[49717] = i[97];
  assign o[49718] = i[97];
  assign o[49719] = i[97];
  assign o[49720] = i[97];
  assign o[49721] = i[97];
  assign o[49722] = i[97];
  assign o[49723] = i[97];
  assign o[49724] = i[97];
  assign o[49725] = i[97];
  assign o[49726] = i[97];
  assign o[49727] = i[97];
  assign o[49728] = i[97];
  assign o[49729] = i[97];
  assign o[49730] = i[97];
  assign o[49731] = i[97];
  assign o[49732] = i[97];
  assign o[49733] = i[97];
  assign o[49734] = i[97];
  assign o[49735] = i[97];
  assign o[49736] = i[97];
  assign o[49737] = i[97];
  assign o[49738] = i[97];
  assign o[49739] = i[97];
  assign o[49740] = i[97];
  assign o[49741] = i[97];
  assign o[49742] = i[97];
  assign o[49743] = i[97];
  assign o[49744] = i[97];
  assign o[49745] = i[97];
  assign o[49746] = i[97];
  assign o[49747] = i[97];
  assign o[49748] = i[97];
  assign o[49749] = i[97];
  assign o[49750] = i[97];
  assign o[49751] = i[97];
  assign o[49752] = i[97];
  assign o[49753] = i[97];
  assign o[49754] = i[97];
  assign o[49755] = i[97];
  assign o[49756] = i[97];
  assign o[49757] = i[97];
  assign o[49758] = i[97];
  assign o[49759] = i[97];
  assign o[49760] = i[97];
  assign o[49761] = i[97];
  assign o[49762] = i[97];
  assign o[49763] = i[97];
  assign o[49764] = i[97];
  assign o[49765] = i[97];
  assign o[49766] = i[97];
  assign o[49767] = i[97];
  assign o[49768] = i[97];
  assign o[49769] = i[97];
  assign o[49770] = i[97];
  assign o[49771] = i[97];
  assign o[49772] = i[97];
  assign o[49773] = i[97];
  assign o[49774] = i[97];
  assign o[49775] = i[97];
  assign o[49776] = i[97];
  assign o[49777] = i[97];
  assign o[49778] = i[97];
  assign o[49779] = i[97];
  assign o[49780] = i[97];
  assign o[49781] = i[97];
  assign o[49782] = i[97];
  assign o[49783] = i[97];
  assign o[49784] = i[97];
  assign o[49785] = i[97];
  assign o[49786] = i[97];
  assign o[49787] = i[97];
  assign o[49788] = i[97];
  assign o[49789] = i[97];
  assign o[49790] = i[97];
  assign o[49791] = i[97];
  assign o[49792] = i[97];
  assign o[49793] = i[97];
  assign o[49794] = i[97];
  assign o[49795] = i[97];
  assign o[49796] = i[97];
  assign o[49797] = i[97];
  assign o[49798] = i[97];
  assign o[49799] = i[97];
  assign o[49800] = i[97];
  assign o[49801] = i[97];
  assign o[49802] = i[97];
  assign o[49803] = i[97];
  assign o[49804] = i[97];
  assign o[49805] = i[97];
  assign o[49806] = i[97];
  assign o[49807] = i[97];
  assign o[49808] = i[97];
  assign o[49809] = i[97];
  assign o[49810] = i[97];
  assign o[49811] = i[97];
  assign o[49812] = i[97];
  assign o[49813] = i[97];
  assign o[49814] = i[97];
  assign o[49815] = i[97];
  assign o[49816] = i[97];
  assign o[49817] = i[97];
  assign o[49818] = i[97];
  assign o[49819] = i[97];
  assign o[49820] = i[97];
  assign o[49821] = i[97];
  assign o[49822] = i[97];
  assign o[49823] = i[97];
  assign o[49824] = i[97];
  assign o[49825] = i[97];
  assign o[49826] = i[97];
  assign o[49827] = i[97];
  assign o[49828] = i[97];
  assign o[49829] = i[97];
  assign o[49830] = i[97];
  assign o[49831] = i[97];
  assign o[49832] = i[97];
  assign o[49833] = i[97];
  assign o[49834] = i[97];
  assign o[49835] = i[97];
  assign o[49836] = i[97];
  assign o[49837] = i[97];
  assign o[49838] = i[97];
  assign o[49839] = i[97];
  assign o[49840] = i[97];
  assign o[49841] = i[97];
  assign o[49842] = i[97];
  assign o[49843] = i[97];
  assign o[49844] = i[97];
  assign o[49845] = i[97];
  assign o[49846] = i[97];
  assign o[49847] = i[97];
  assign o[49848] = i[97];
  assign o[49849] = i[97];
  assign o[49850] = i[97];
  assign o[49851] = i[97];
  assign o[49852] = i[97];
  assign o[49853] = i[97];
  assign o[49854] = i[97];
  assign o[49855] = i[97];
  assign o[49856] = i[97];
  assign o[49857] = i[97];
  assign o[49858] = i[97];
  assign o[49859] = i[97];
  assign o[49860] = i[97];
  assign o[49861] = i[97];
  assign o[49862] = i[97];
  assign o[49863] = i[97];
  assign o[49864] = i[97];
  assign o[49865] = i[97];
  assign o[49866] = i[97];
  assign o[49867] = i[97];
  assign o[49868] = i[97];
  assign o[49869] = i[97];
  assign o[49870] = i[97];
  assign o[49871] = i[97];
  assign o[49872] = i[97];
  assign o[49873] = i[97];
  assign o[49874] = i[97];
  assign o[49875] = i[97];
  assign o[49876] = i[97];
  assign o[49877] = i[97];
  assign o[49878] = i[97];
  assign o[49879] = i[97];
  assign o[49880] = i[97];
  assign o[49881] = i[97];
  assign o[49882] = i[97];
  assign o[49883] = i[97];
  assign o[49884] = i[97];
  assign o[49885] = i[97];
  assign o[49886] = i[97];
  assign o[49887] = i[97];
  assign o[49888] = i[97];
  assign o[49889] = i[97];
  assign o[49890] = i[97];
  assign o[49891] = i[97];
  assign o[49892] = i[97];
  assign o[49893] = i[97];
  assign o[49894] = i[97];
  assign o[49895] = i[97];
  assign o[49896] = i[97];
  assign o[49897] = i[97];
  assign o[49898] = i[97];
  assign o[49899] = i[97];
  assign o[49900] = i[97];
  assign o[49901] = i[97];
  assign o[49902] = i[97];
  assign o[49903] = i[97];
  assign o[49904] = i[97];
  assign o[49905] = i[97];
  assign o[49906] = i[97];
  assign o[49907] = i[97];
  assign o[49908] = i[97];
  assign o[49909] = i[97];
  assign o[49910] = i[97];
  assign o[49911] = i[97];
  assign o[49912] = i[97];
  assign o[49913] = i[97];
  assign o[49914] = i[97];
  assign o[49915] = i[97];
  assign o[49916] = i[97];
  assign o[49917] = i[97];
  assign o[49918] = i[97];
  assign o[49919] = i[97];
  assign o[49920] = i[97];
  assign o[49921] = i[97];
  assign o[49922] = i[97];
  assign o[49923] = i[97];
  assign o[49924] = i[97];
  assign o[49925] = i[97];
  assign o[49926] = i[97];
  assign o[49927] = i[97];
  assign o[49928] = i[97];
  assign o[49929] = i[97];
  assign o[49930] = i[97];
  assign o[49931] = i[97];
  assign o[49932] = i[97];
  assign o[49933] = i[97];
  assign o[49934] = i[97];
  assign o[49935] = i[97];
  assign o[49936] = i[97];
  assign o[49937] = i[97];
  assign o[49938] = i[97];
  assign o[49939] = i[97];
  assign o[49940] = i[97];
  assign o[49941] = i[97];
  assign o[49942] = i[97];
  assign o[49943] = i[97];
  assign o[49944] = i[97];
  assign o[49945] = i[97];
  assign o[49946] = i[97];
  assign o[49947] = i[97];
  assign o[49948] = i[97];
  assign o[49949] = i[97];
  assign o[49950] = i[97];
  assign o[49951] = i[97];
  assign o[49952] = i[97];
  assign o[49953] = i[97];
  assign o[49954] = i[97];
  assign o[49955] = i[97];
  assign o[49956] = i[97];
  assign o[49957] = i[97];
  assign o[49958] = i[97];
  assign o[49959] = i[97];
  assign o[49960] = i[97];
  assign o[49961] = i[97];
  assign o[49962] = i[97];
  assign o[49963] = i[97];
  assign o[49964] = i[97];
  assign o[49965] = i[97];
  assign o[49966] = i[97];
  assign o[49967] = i[97];
  assign o[49968] = i[97];
  assign o[49969] = i[97];
  assign o[49970] = i[97];
  assign o[49971] = i[97];
  assign o[49972] = i[97];
  assign o[49973] = i[97];
  assign o[49974] = i[97];
  assign o[49975] = i[97];
  assign o[49976] = i[97];
  assign o[49977] = i[97];
  assign o[49978] = i[97];
  assign o[49979] = i[97];
  assign o[49980] = i[97];
  assign o[49981] = i[97];
  assign o[49982] = i[97];
  assign o[49983] = i[97];
  assign o[49984] = i[97];
  assign o[49985] = i[97];
  assign o[49986] = i[97];
  assign o[49987] = i[97];
  assign o[49988] = i[97];
  assign o[49989] = i[97];
  assign o[49990] = i[97];
  assign o[49991] = i[97];
  assign o[49992] = i[97];
  assign o[49993] = i[97];
  assign o[49994] = i[97];
  assign o[49995] = i[97];
  assign o[49996] = i[97];
  assign o[49997] = i[97];
  assign o[49998] = i[97];
  assign o[49999] = i[97];
  assign o[50000] = i[97];
  assign o[50001] = i[97];
  assign o[50002] = i[97];
  assign o[50003] = i[97];
  assign o[50004] = i[97];
  assign o[50005] = i[97];
  assign o[50006] = i[97];
  assign o[50007] = i[97];
  assign o[50008] = i[97];
  assign o[50009] = i[97];
  assign o[50010] = i[97];
  assign o[50011] = i[97];
  assign o[50012] = i[97];
  assign o[50013] = i[97];
  assign o[50014] = i[97];
  assign o[50015] = i[97];
  assign o[50016] = i[97];
  assign o[50017] = i[97];
  assign o[50018] = i[97];
  assign o[50019] = i[97];
  assign o[50020] = i[97];
  assign o[50021] = i[97];
  assign o[50022] = i[97];
  assign o[50023] = i[97];
  assign o[50024] = i[97];
  assign o[50025] = i[97];
  assign o[50026] = i[97];
  assign o[50027] = i[97];
  assign o[50028] = i[97];
  assign o[50029] = i[97];
  assign o[50030] = i[97];
  assign o[50031] = i[97];
  assign o[50032] = i[97];
  assign o[50033] = i[97];
  assign o[50034] = i[97];
  assign o[50035] = i[97];
  assign o[50036] = i[97];
  assign o[50037] = i[97];
  assign o[50038] = i[97];
  assign o[50039] = i[97];
  assign o[50040] = i[97];
  assign o[50041] = i[97];
  assign o[50042] = i[97];
  assign o[50043] = i[97];
  assign o[50044] = i[97];
  assign o[50045] = i[97];
  assign o[50046] = i[97];
  assign o[50047] = i[97];
  assign o[50048] = i[97];
  assign o[50049] = i[97];
  assign o[50050] = i[97];
  assign o[50051] = i[97];
  assign o[50052] = i[97];
  assign o[50053] = i[97];
  assign o[50054] = i[97];
  assign o[50055] = i[97];
  assign o[50056] = i[97];
  assign o[50057] = i[97];
  assign o[50058] = i[97];
  assign o[50059] = i[97];
  assign o[50060] = i[97];
  assign o[50061] = i[97];
  assign o[50062] = i[97];
  assign o[50063] = i[97];
  assign o[50064] = i[97];
  assign o[50065] = i[97];
  assign o[50066] = i[97];
  assign o[50067] = i[97];
  assign o[50068] = i[97];
  assign o[50069] = i[97];
  assign o[50070] = i[97];
  assign o[50071] = i[97];
  assign o[50072] = i[97];
  assign o[50073] = i[97];
  assign o[50074] = i[97];
  assign o[50075] = i[97];
  assign o[50076] = i[97];
  assign o[50077] = i[97];
  assign o[50078] = i[97];
  assign o[50079] = i[97];
  assign o[50080] = i[97];
  assign o[50081] = i[97];
  assign o[50082] = i[97];
  assign o[50083] = i[97];
  assign o[50084] = i[97];
  assign o[50085] = i[97];
  assign o[50086] = i[97];
  assign o[50087] = i[97];
  assign o[50088] = i[97];
  assign o[50089] = i[97];
  assign o[50090] = i[97];
  assign o[50091] = i[97];
  assign o[50092] = i[97];
  assign o[50093] = i[97];
  assign o[50094] = i[97];
  assign o[50095] = i[97];
  assign o[50096] = i[97];
  assign o[50097] = i[97];
  assign o[50098] = i[97];
  assign o[50099] = i[97];
  assign o[50100] = i[97];
  assign o[50101] = i[97];
  assign o[50102] = i[97];
  assign o[50103] = i[97];
  assign o[50104] = i[97];
  assign o[50105] = i[97];
  assign o[50106] = i[97];
  assign o[50107] = i[97];
  assign o[50108] = i[97];
  assign o[50109] = i[97];
  assign o[50110] = i[97];
  assign o[50111] = i[97];
  assign o[50112] = i[97];
  assign o[50113] = i[97];
  assign o[50114] = i[97];
  assign o[50115] = i[97];
  assign o[50116] = i[97];
  assign o[50117] = i[97];
  assign o[50118] = i[97];
  assign o[50119] = i[97];
  assign o[50120] = i[97];
  assign o[50121] = i[97];
  assign o[50122] = i[97];
  assign o[50123] = i[97];
  assign o[50124] = i[97];
  assign o[50125] = i[97];
  assign o[50126] = i[97];
  assign o[50127] = i[97];
  assign o[50128] = i[97];
  assign o[50129] = i[97];
  assign o[50130] = i[97];
  assign o[50131] = i[97];
  assign o[50132] = i[97];
  assign o[50133] = i[97];
  assign o[50134] = i[97];
  assign o[50135] = i[97];
  assign o[50136] = i[97];
  assign o[50137] = i[97];
  assign o[50138] = i[97];
  assign o[50139] = i[97];
  assign o[50140] = i[97];
  assign o[50141] = i[97];
  assign o[50142] = i[97];
  assign o[50143] = i[97];
  assign o[50144] = i[97];
  assign o[50145] = i[97];
  assign o[50146] = i[97];
  assign o[50147] = i[97];
  assign o[50148] = i[97];
  assign o[50149] = i[97];
  assign o[50150] = i[97];
  assign o[50151] = i[97];
  assign o[50152] = i[97];
  assign o[50153] = i[97];
  assign o[50154] = i[97];
  assign o[50155] = i[97];
  assign o[50156] = i[97];
  assign o[50157] = i[97];
  assign o[50158] = i[97];
  assign o[50159] = i[97];
  assign o[50160] = i[97];
  assign o[50161] = i[97];
  assign o[50162] = i[97];
  assign o[50163] = i[97];
  assign o[50164] = i[97];
  assign o[50165] = i[97];
  assign o[50166] = i[97];
  assign o[50167] = i[97];
  assign o[50168] = i[97];
  assign o[50169] = i[97];
  assign o[50170] = i[97];
  assign o[50171] = i[97];
  assign o[50172] = i[97];
  assign o[50173] = i[97];
  assign o[50174] = i[97];
  assign o[50175] = i[97];
  assign o[49152] = i[96];
  assign o[49153] = i[96];
  assign o[49154] = i[96];
  assign o[49155] = i[96];
  assign o[49156] = i[96];
  assign o[49157] = i[96];
  assign o[49158] = i[96];
  assign o[49159] = i[96];
  assign o[49160] = i[96];
  assign o[49161] = i[96];
  assign o[49162] = i[96];
  assign o[49163] = i[96];
  assign o[49164] = i[96];
  assign o[49165] = i[96];
  assign o[49166] = i[96];
  assign o[49167] = i[96];
  assign o[49168] = i[96];
  assign o[49169] = i[96];
  assign o[49170] = i[96];
  assign o[49171] = i[96];
  assign o[49172] = i[96];
  assign o[49173] = i[96];
  assign o[49174] = i[96];
  assign o[49175] = i[96];
  assign o[49176] = i[96];
  assign o[49177] = i[96];
  assign o[49178] = i[96];
  assign o[49179] = i[96];
  assign o[49180] = i[96];
  assign o[49181] = i[96];
  assign o[49182] = i[96];
  assign o[49183] = i[96];
  assign o[49184] = i[96];
  assign o[49185] = i[96];
  assign o[49186] = i[96];
  assign o[49187] = i[96];
  assign o[49188] = i[96];
  assign o[49189] = i[96];
  assign o[49190] = i[96];
  assign o[49191] = i[96];
  assign o[49192] = i[96];
  assign o[49193] = i[96];
  assign o[49194] = i[96];
  assign o[49195] = i[96];
  assign o[49196] = i[96];
  assign o[49197] = i[96];
  assign o[49198] = i[96];
  assign o[49199] = i[96];
  assign o[49200] = i[96];
  assign o[49201] = i[96];
  assign o[49202] = i[96];
  assign o[49203] = i[96];
  assign o[49204] = i[96];
  assign o[49205] = i[96];
  assign o[49206] = i[96];
  assign o[49207] = i[96];
  assign o[49208] = i[96];
  assign o[49209] = i[96];
  assign o[49210] = i[96];
  assign o[49211] = i[96];
  assign o[49212] = i[96];
  assign o[49213] = i[96];
  assign o[49214] = i[96];
  assign o[49215] = i[96];
  assign o[49216] = i[96];
  assign o[49217] = i[96];
  assign o[49218] = i[96];
  assign o[49219] = i[96];
  assign o[49220] = i[96];
  assign o[49221] = i[96];
  assign o[49222] = i[96];
  assign o[49223] = i[96];
  assign o[49224] = i[96];
  assign o[49225] = i[96];
  assign o[49226] = i[96];
  assign o[49227] = i[96];
  assign o[49228] = i[96];
  assign o[49229] = i[96];
  assign o[49230] = i[96];
  assign o[49231] = i[96];
  assign o[49232] = i[96];
  assign o[49233] = i[96];
  assign o[49234] = i[96];
  assign o[49235] = i[96];
  assign o[49236] = i[96];
  assign o[49237] = i[96];
  assign o[49238] = i[96];
  assign o[49239] = i[96];
  assign o[49240] = i[96];
  assign o[49241] = i[96];
  assign o[49242] = i[96];
  assign o[49243] = i[96];
  assign o[49244] = i[96];
  assign o[49245] = i[96];
  assign o[49246] = i[96];
  assign o[49247] = i[96];
  assign o[49248] = i[96];
  assign o[49249] = i[96];
  assign o[49250] = i[96];
  assign o[49251] = i[96];
  assign o[49252] = i[96];
  assign o[49253] = i[96];
  assign o[49254] = i[96];
  assign o[49255] = i[96];
  assign o[49256] = i[96];
  assign o[49257] = i[96];
  assign o[49258] = i[96];
  assign o[49259] = i[96];
  assign o[49260] = i[96];
  assign o[49261] = i[96];
  assign o[49262] = i[96];
  assign o[49263] = i[96];
  assign o[49264] = i[96];
  assign o[49265] = i[96];
  assign o[49266] = i[96];
  assign o[49267] = i[96];
  assign o[49268] = i[96];
  assign o[49269] = i[96];
  assign o[49270] = i[96];
  assign o[49271] = i[96];
  assign o[49272] = i[96];
  assign o[49273] = i[96];
  assign o[49274] = i[96];
  assign o[49275] = i[96];
  assign o[49276] = i[96];
  assign o[49277] = i[96];
  assign o[49278] = i[96];
  assign o[49279] = i[96];
  assign o[49280] = i[96];
  assign o[49281] = i[96];
  assign o[49282] = i[96];
  assign o[49283] = i[96];
  assign o[49284] = i[96];
  assign o[49285] = i[96];
  assign o[49286] = i[96];
  assign o[49287] = i[96];
  assign o[49288] = i[96];
  assign o[49289] = i[96];
  assign o[49290] = i[96];
  assign o[49291] = i[96];
  assign o[49292] = i[96];
  assign o[49293] = i[96];
  assign o[49294] = i[96];
  assign o[49295] = i[96];
  assign o[49296] = i[96];
  assign o[49297] = i[96];
  assign o[49298] = i[96];
  assign o[49299] = i[96];
  assign o[49300] = i[96];
  assign o[49301] = i[96];
  assign o[49302] = i[96];
  assign o[49303] = i[96];
  assign o[49304] = i[96];
  assign o[49305] = i[96];
  assign o[49306] = i[96];
  assign o[49307] = i[96];
  assign o[49308] = i[96];
  assign o[49309] = i[96];
  assign o[49310] = i[96];
  assign o[49311] = i[96];
  assign o[49312] = i[96];
  assign o[49313] = i[96];
  assign o[49314] = i[96];
  assign o[49315] = i[96];
  assign o[49316] = i[96];
  assign o[49317] = i[96];
  assign o[49318] = i[96];
  assign o[49319] = i[96];
  assign o[49320] = i[96];
  assign o[49321] = i[96];
  assign o[49322] = i[96];
  assign o[49323] = i[96];
  assign o[49324] = i[96];
  assign o[49325] = i[96];
  assign o[49326] = i[96];
  assign o[49327] = i[96];
  assign o[49328] = i[96];
  assign o[49329] = i[96];
  assign o[49330] = i[96];
  assign o[49331] = i[96];
  assign o[49332] = i[96];
  assign o[49333] = i[96];
  assign o[49334] = i[96];
  assign o[49335] = i[96];
  assign o[49336] = i[96];
  assign o[49337] = i[96];
  assign o[49338] = i[96];
  assign o[49339] = i[96];
  assign o[49340] = i[96];
  assign o[49341] = i[96];
  assign o[49342] = i[96];
  assign o[49343] = i[96];
  assign o[49344] = i[96];
  assign o[49345] = i[96];
  assign o[49346] = i[96];
  assign o[49347] = i[96];
  assign o[49348] = i[96];
  assign o[49349] = i[96];
  assign o[49350] = i[96];
  assign o[49351] = i[96];
  assign o[49352] = i[96];
  assign o[49353] = i[96];
  assign o[49354] = i[96];
  assign o[49355] = i[96];
  assign o[49356] = i[96];
  assign o[49357] = i[96];
  assign o[49358] = i[96];
  assign o[49359] = i[96];
  assign o[49360] = i[96];
  assign o[49361] = i[96];
  assign o[49362] = i[96];
  assign o[49363] = i[96];
  assign o[49364] = i[96];
  assign o[49365] = i[96];
  assign o[49366] = i[96];
  assign o[49367] = i[96];
  assign o[49368] = i[96];
  assign o[49369] = i[96];
  assign o[49370] = i[96];
  assign o[49371] = i[96];
  assign o[49372] = i[96];
  assign o[49373] = i[96];
  assign o[49374] = i[96];
  assign o[49375] = i[96];
  assign o[49376] = i[96];
  assign o[49377] = i[96];
  assign o[49378] = i[96];
  assign o[49379] = i[96];
  assign o[49380] = i[96];
  assign o[49381] = i[96];
  assign o[49382] = i[96];
  assign o[49383] = i[96];
  assign o[49384] = i[96];
  assign o[49385] = i[96];
  assign o[49386] = i[96];
  assign o[49387] = i[96];
  assign o[49388] = i[96];
  assign o[49389] = i[96];
  assign o[49390] = i[96];
  assign o[49391] = i[96];
  assign o[49392] = i[96];
  assign o[49393] = i[96];
  assign o[49394] = i[96];
  assign o[49395] = i[96];
  assign o[49396] = i[96];
  assign o[49397] = i[96];
  assign o[49398] = i[96];
  assign o[49399] = i[96];
  assign o[49400] = i[96];
  assign o[49401] = i[96];
  assign o[49402] = i[96];
  assign o[49403] = i[96];
  assign o[49404] = i[96];
  assign o[49405] = i[96];
  assign o[49406] = i[96];
  assign o[49407] = i[96];
  assign o[49408] = i[96];
  assign o[49409] = i[96];
  assign o[49410] = i[96];
  assign o[49411] = i[96];
  assign o[49412] = i[96];
  assign o[49413] = i[96];
  assign o[49414] = i[96];
  assign o[49415] = i[96];
  assign o[49416] = i[96];
  assign o[49417] = i[96];
  assign o[49418] = i[96];
  assign o[49419] = i[96];
  assign o[49420] = i[96];
  assign o[49421] = i[96];
  assign o[49422] = i[96];
  assign o[49423] = i[96];
  assign o[49424] = i[96];
  assign o[49425] = i[96];
  assign o[49426] = i[96];
  assign o[49427] = i[96];
  assign o[49428] = i[96];
  assign o[49429] = i[96];
  assign o[49430] = i[96];
  assign o[49431] = i[96];
  assign o[49432] = i[96];
  assign o[49433] = i[96];
  assign o[49434] = i[96];
  assign o[49435] = i[96];
  assign o[49436] = i[96];
  assign o[49437] = i[96];
  assign o[49438] = i[96];
  assign o[49439] = i[96];
  assign o[49440] = i[96];
  assign o[49441] = i[96];
  assign o[49442] = i[96];
  assign o[49443] = i[96];
  assign o[49444] = i[96];
  assign o[49445] = i[96];
  assign o[49446] = i[96];
  assign o[49447] = i[96];
  assign o[49448] = i[96];
  assign o[49449] = i[96];
  assign o[49450] = i[96];
  assign o[49451] = i[96];
  assign o[49452] = i[96];
  assign o[49453] = i[96];
  assign o[49454] = i[96];
  assign o[49455] = i[96];
  assign o[49456] = i[96];
  assign o[49457] = i[96];
  assign o[49458] = i[96];
  assign o[49459] = i[96];
  assign o[49460] = i[96];
  assign o[49461] = i[96];
  assign o[49462] = i[96];
  assign o[49463] = i[96];
  assign o[49464] = i[96];
  assign o[49465] = i[96];
  assign o[49466] = i[96];
  assign o[49467] = i[96];
  assign o[49468] = i[96];
  assign o[49469] = i[96];
  assign o[49470] = i[96];
  assign o[49471] = i[96];
  assign o[49472] = i[96];
  assign o[49473] = i[96];
  assign o[49474] = i[96];
  assign o[49475] = i[96];
  assign o[49476] = i[96];
  assign o[49477] = i[96];
  assign o[49478] = i[96];
  assign o[49479] = i[96];
  assign o[49480] = i[96];
  assign o[49481] = i[96];
  assign o[49482] = i[96];
  assign o[49483] = i[96];
  assign o[49484] = i[96];
  assign o[49485] = i[96];
  assign o[49486] = i[96];
  assign o[49487] = i[96];
  assign o[49488] = i[96];
  assign o[49489] = i[96];
  assign o[49490] = i[96];
  assign o[49491] = i[96];
  assign o[49492] = i[96];
  assign o[49493] = i[96];
  assign o[49494] = i[96];
  assign o[49495] = i[96];
  assign o[49496] = i[96];
  assign o[49497] = i[96];
  assign o[49498] = i[96];
  assign o[49499] = i[96];
  assign o[49500] = i[96];
  assign o[49501] = i[96];
  assign o[49502] = i[96];
  assign o[49503] = i[96];
  assign o[49504] = i[96];
  assign o[49505] = i[96];
  assign o[49506] = i[96];
  assign o[49507] = i[96];
  assign o[49508] = i[96];
  assign o[49509] = i[96];
  assign o[49510] = i[96];
  assign o[49511] = i[96];
  assign o[49512] = i[96];
  assign o[49513] = i[96];
  assign o[49514] = i[96];
  assign o[49515] = i[96];
  assign o[49516] = i[96];
  assign o[49517] = i[96];
  assign o[49518] = i[96];
  assign o[49519] = i[96];
  assign o[49520] = i[96];
  assign o[49521] = i[96];
  assign o[49522] = i[96];
  assign o[49523] = i[96];
  assign o[49524] = i[96];
  assign o[49525] = i[96];
  assign o[49526] = i[96];
  assign o[49527] = i[96];
  assign o[49528] = i[96];
  assign o[49529] = i[96];
  assign o[49530] = i[96];
  assign o[49531] = i[96];
  assign o[49532] = i[96];
  assign o[49533] = i[96];
  assign o[49534] = i[96];
  assign o[49535] = i[96];
  assign o[49536] = i[96];
  assign o[49537] = i[96];
  assign o[49538] = i[96];
  assign o[49539] = i[96];
  assign o[49540] = i[96];
  assign o[49541] = i[96];
  assign o[49542] = i[96];
  assign o[49543] = i[96];
  assign o[49544] = i[96];
  assign o[49545] = i[96];
  assign o[49546] = i[96];
  assign o[49547] = i[96];
  assign o[49548] = i[96];
  assign o[49549] = i[96];
  assign o[49550] = i[96];
  assign o[49551] = i[96];
  assign o[49552] = i[96];
  assign o[49553] = i[96];
  assign o[49554] = i[96];
  assign o[49555] = i[96];
  assign o[49556] = i[96];
  assign o[49557] = i[96];
  assign o[49558] = i[96];
  assign o[49559] = i[96];
  assign o[49560] = i[96];
  assign o[49561] = i[96];
  assign o[49562] = i[96];
  assign o[49563] = i[96];
  assign o[49564] = i[96];
  assign o[49565] = i[96];
  assign o[49566] = i[96];
  assign o[49567] = i[96];
  assign o[49568] = i[96];
  assign o[49569] = i[96];
  assign o[49570] = i[96];
  assign o[49571] = i[96];
  assign o[49572] = i[96];
  assign o[49573] = i[96];
  assign o[49574] = i[96];
  assign o[49575] = i[96];
  assign o[49576] = i[96];
  assign o[49577] = i[96];
  assign o[49578] = i[96];
  assign o[49579] = i[96];
  assign o[49580] = i[96];
  assign o[49581] = i[96];
  assign o[49582] = i[96];
  assign o[49583] = i[96];
  assign o[49584] = i[96];
  assign o[49585] = i[96];
  assign o[49586] = i[96];
  assign o[49587] = i[96];
  assign o[49588] = i[96];
  assign o[49589] = i[96];
  assign o[49590] = i[96];
  assign o[49591] = i[96];
  assign o[49592] = i[96];
  assign o[49593] = i[96];
  assign o[49594] = i[96];
  assign o[49595] = i[96];
  assign o[49596] = i[96];
  assign o[49597] = i[96];
  assign o[49598] = i[96];
  assign o[49599] = i[96];
  assign o[49600] = i[96];
  assign o[49601] = i[96];
  assign o[49602] = i[96];
  assign o[49603] = i[96];
  assign o[49604] = i[96];
  assign o[49605] = i[96];
  assign o[49606] = i[96];
  assign o[49607] = i[96];
  assign o[49608] = i[96];
  assign o[49609] = i[96];
  assign o[49610] = i[96];
  assign o[49611] = i[96];
  assign o[49612] = i[96];
  assign o[49613] = i[96];
  assign o[49614] = i[96];
  assign o[49615] = i[96];
  assign o[49616] = i[96];
  assign o[49617] = i[96];
  assign o[49618] = i[96];
  assign o[49619] = i[96];
  assign o[49620] = i[96];
  assign o[49621] = i[96];
  assign o[49622] = i[96];
  assign o[49623] = i[96];
  assign o[49624] = i[96];
  assign o[49625] = i[96];
  assign o[49626] = i[96];
  assign o[49627] = i[96];
  assign o[49628] = i[96];
  assign o[49629] = i[96];
  assign o[49630] = i[96];
  assign o[49631] = i[96];
  assign o[49632] = i[96];
  assign o[49633] = i[96];
  assign o[49634] = i[96];
  assign o[49635] = i[96];
  assign o[49636] = i[96];
  assign o[49637] = i[96];
  assign o[49638] = i[96];
  assign o[49639] = i[96];
  assign o[49640] = i[96];
  assign o[49641] = i[96];
  assign o[49642] = i[96];
  assign o[49643] = i[96];
  assign o[49644] = i[96];
  assign o[49645] = i[96];
  assign o[49646] = i[96];
  assign o[49647] = i[96];
  assign o[49648] = i[96];
  assign o[49649] = i[96];
  assign o[49650] = i[96];
  assign o[49651] = i[96];
  assign o[49652] = i[96];
  assign o[49653] = i[96];
  assign o[49654] = i[96];
  assign o[49655] = i[96];
  assign o[49656] = i[96];
  assign o[49657] = i[96];
  assign o[49658] = i[96];
  assign o[49659] = i[96];
  assign o[49660] = i[96];
  assign o[49661] = i[96];
  assign o[49662] = i[96];
  assign o[49663] = i[96];
  assign o[48640] = i[95];
  assign o[48641] = i[95];
  assign o[48642] = i[95];
  assign o[48643] = i[95];
  assign o[48644] = i[95];
  assign o[48645] = i[95];
  assign o[48646] = i[95];
  assign o[48647] = i[95];
  assign o[48648] = i[95];
  assign o[48649] = i[95];
  assign o[48650] = i[95];
  assign o[48651] = i[95];
  assign o[48652] = i[95];
  assign o[48653] = i[95];
  assign o[48654] = i[95];
  assign o[48655] = i[95];
  assign o[48656] = i[95];
  assign o[48657] = i[95];
  assign o[48658] = i[95];
  assign o[48659] = i[95];
  assign o[48660] = i[95];
  assign o[48661] = i[95];
  assign o[48662] = i[95];
  assign o[48663] = i[95];
  assign o[48664] = i[95];
  assign o[48665] = i[95];
  assign o[48666] = i[95];
  assign o[48667] = i[95];
  assign o[48668] = i[95];
  assign o[48669] = i[95];
  assign o[48670] = i[95];
  assign o[48671] = i[95];
  assign o[48672] = i[95];
  assign o[48673] = i[95];
  assign o[48674] = i[95];
  assign o[48675] = i[95];
  assign o[48676] = i[95];
  assign o[48677] = i[95];
  assign o[48678] = i[95];
  assign o[48679] = i[95];
  assign o[48680] = i[95];
  assign o[48681] = i[95];
  assign o[48682] = i[95];
  assign o[48683] = i[95];
  assign o[48684] = i[95];
  assign o[48685] = i[95];
  assign o[48686] = i[95];
  assign o[48687] = i[95];
  assign o[48688] = i[95];
  assign o[48689] = i[95];
  assign o[48690] = i[95];
  assign o[48691] = i[95];
  assign o[48692] = i[95];
  assign o[48693] = i[95];
  assign o[48694] = i[95];
  assign o[48695] = i[95];
  assign o[48696] = i[95];
  assign o[48697] = i[95];
  assign o[48698] = i[95];
  assign o[48699] = i[95];
  assign o[48700] = i[95];
  assign o[48701] = i[95];
  assign o[48702] = i[95];
  assign o[48703] = i[95];
  assign o[48704] = i[95];
  assign o[48705] = i[95];
  assign o[48706] = i[95];
  assign o[48707] = i[95];
  assign o[48708] = i[95];
  assign o[48709] = i[95];
  assign o[48710] = i[95];
  assign o[48711] = i[95];
  assign o[48712] = i[95];
  assign o[48713] = i[95];
  assign o[48714] = i[95];
  assign o[48715] = i[95];
  assign o[48716] = i[95];
  assign o[48717] = i[95];
  assign o[48718] = i[95];
  assign o[48719] = i[95];
  assign o[48720] = i[95];
  assign o[48721] = i[95];
  assign o[48722] = i[95];
  assign o[48723] = i[95];
  assign o[48724] = i[95];
  assign o[48725] = i[95];
  assign o[48726] = i[95];
  assign o[48727] = i[95];
  assign o[48728] = i[95];
  assign o[48729] = i[95];
  assign o[48730] = i[95];
  assign o[48731] = i[95];
  assign o[48732] = i[95];
  assign o[48733] = i[95];
  assign o[48734] = i[95];
  assign o[48735] = i[95];
  assign o[48736] = i[95];
  assign o[48737] = i[95];
  assign o[48738] = i[95];
  assign o[48739] = i[95];
  assign o[48740] = i[95];
  assign o[48741] = i[95];
  assign o[48742] = i[95];
  assign o[48743] = i[95];
  assign o[48744] = i[95];
  assign o[48745] = i[95];
  assign o[48746] = i[95];
  assign o[48747] = i[95];
  assign o[48748] = i[95];
  assign o[48749] = i[95];
  assign o[48750] = i[95];
  assign o[48751] = i[95];
  assign o[48752] = i[95];
  assign o[48753] = i[95];
  assign o[48754] = i[95];
  assign o[48755] = i[95];
  assign o[48756] = i[95];
  assign o[48757] = i[95];
  assign o[48758] = i[95];
  assign o[48759] = i[95];
  assign o[48760] = i[95];
  assign o[48761] = i[95];
  assign o[48762] = i[95];
  assign o[48763] = i[95];
  assign o[48764] = i[95];
  assign o[48765] = i[95];
  assign o[48766] = i[95];
  assign o[48767] = i[95];
  assign o[48768] = i[95];
  assign o[48769] = i[95];
  assign o[48770] = i[95];
  assign o[48771] = i[95];
  assign o[48772] = i[95];
  assign o[48773] = i[95];
  assign o[48774] = i[95];
  assign o[48775] = i[95];
  assign o[48776] = i[95];
  assign o[48777] = i[95];
  assign o[48778] = i[95];
  assign o[48779] = i[95];
  assign o[48780] = i[95];
  assign o[48781] = i[95];
  assign o[48782] = i[95];
  assign o[48783] = i[95];
  assign o[48784] = i[95];
  assign o[48785] = i[95];
  assign o[48786] = i[95];
  assign o[48787] = i[95];
  assign o[48788] = i[95];
  assign o[48789] = i[95];
  assign o[48790] = i[95];
  assign o[48791] = i[95];
  assign o[48792] = i[95];
  assign o[48793] = i[95];
  assign o[48794] = i[95];
  assign o[48795] = i[95];
  assign o[48796] = i[95];
  assign o[48797] = i[95];
  assign o[48798] = i[95];
  assign o[48799] = i[95];
  assign o[48800] = i[95];
  assign o[48801] = i[95];
  assign o[48802] = i[95];
  assign o[48803] = i[95];
  assign o[48804] = i[95];
  assign o[48805] = i[95];
  assign o[48806] = i[95];
  assign o[48807] = i[95];
  assign o[48808] = i[95];
  assign o[48809] = i[95];
  assign o[48810] = i[95];
  assign o[48811] = i[95];
  assign o[48812] = i[95];
  assign o[48813] = i[95];
  assign o[48814] = i[95];
  assign o[48815] = i[95];
  assign o[48816] = i[95];
  assign o[48817] = i[95];
  assign o[48818] = i[95];
  assign o[48819] = i[95];
  assign o[48820] = i[95];
  assign o[48821] = i[95];
  assign o[48822] = i[95];
  assign o[48823] = i[95];
  assign o[48824] = i[95];
  assign o[48825] = i[95];
  assign o[48826] = i[95];
  assign o[48827] = i[95];
  assign o[48828] = i[95];
  assign o[48829] = i[95];
  assign o[48830] = i[95];
  assign o[48831] = i[95];
  assign o[48832] = i[95];
  assign o[48833] = i[95];
  assign o[48834] = i[95];
  assign o[48835] = i[95];
  assign o[48836] = i[95];
  assign o[48837] = i[95];
  assign o[48838] = i[95];
  assign o[48839] = i[95];
  assign o[48840] = i[95];
  assign o[48841] = i[95];
  assign o[48842] = i[95];
  assign o[48843] = i[95];
  assign o[48844] = i[95];
  assign o[48845] = i[95];
  assign o[48846] = i[95];
  assign o[48847] = i[95];
  assign o[48848] = i[95];
  assign o[48849] = i[95];
  assign o[48850] = i[95];
  assign o[48851] = i[95];
  assign o[48852] = i[95];
  assign o[48853] = i[95];
  assign o[48854] = i[95];
  assign o[48855] = i[95];
  assign o[48856] = i[95];
  assign o[48857] = i[95];
  assign o[48858] = i[95];
  assign o[48859] = i[95];
  assign o[48860] = i[95];
  assign o[48861] = i[95];
  assign o[48862] = i[95];
  assign o[48863] = i[95];
  assign o[48864] = i[95];
  assign o[48865] = i[95];
  assign o[48866] = i[95];
  assign o[48867] = i[95];
  assign o[48868] = i[95];
  assign o[48869] = i[95];
  assign o[48870] = i[95];
  assign o[48871] = i[95];
  assign o[48872] = i[95];
  assign o[48873] = i[95];
  assign o[48874] = i[95];
  assign o[48875] = i[95];
  assign o[48876] = i[95];
  assign o[48877] = i[95];
  assign o[48878] = i[95];
  assign o[48879] = i[95];
  assign o[48880] = i[95];
  assign o[48881] = i[95];
  assign o[48882] = i[95];
  assign o[48883] = i[95];
  assign o[48884] = i[95];
  assign o[48885] = i[95];
  assign o[48886] = i[95];
  assign o[48887] = i[95];
  assign o[48888] = i[95];
  assign o[48889] = i[95];
  assign o[48890] = i[95];
  assign o[48891] = i[95];
  assign o[48892] = i[95];
  assign o[48893] = i[95];
  assign o[48894] = i[95];
  assign o[48895] = i[95];
  assign o[48896] = i[95];
  assign o[48897] = i[95];
  assign o[48898] = i[95];
  assign o[48899] = i[95];
  assign o[48900] = i[95];
  assign o[48901] = i[95];
  assign o[48902] = i[95];
  assign o[48903] = i[95];
  assign o[48904] = i[95];
  assign o[48905] = i[95];
  assign o[48906] = i[95];
  assign o[48907] = i[95];
  assign o[48908] = i[95];
  assign o[48909] = i[95];
  assign o[48910] = i[95];
  assign o[48911] = i[95];
  assign o[48912] = i[95];
  assign o[48913] = i[95];
  assign o[48914] = i[95];
  assign o[48915] = i[95];
  assign o[48916] = i[95];
  assign o[48917] = i[95];
  assign o[48918] = i[95];
  assign o[48919] = i[95];
  assign o[48920] = i[95];
  assign o[48921] = i[95];
  assign o[48922] = i[95];
  assign o[48923] = i[95];
  assign o[48924] = i[95];
  assign o[48925] = i[95];
  assign o[48926] = i[95];
  assign o[48927] = i[95];
  assign o[48928] = i[95];
  assign o[48929] = i[95];
  assign o[48930] = i[95];
  assign o[48931] = i[95];
  assign o[48932] = i[95];
  assign o[48933] = i[95];
  assign o[48934] = i[95];
  assign o[48935] = i[95];
  assign o[48936] = i[95];
  assign o[48937] = i[95];
  assign o[48938] = i[95];
  assign o[48939] = i[95];
  assign o[48940] = i[95];
  assign o[48941] = i[95];
  assign o[48942] = i[95];
  assign o[48943] = i[95];
  assign o[48944] = i[95];
  assign o[48945] = i[95];
  assign o[48946] = i[95];
  assign o[48947] = i[95];
  assign o[48948] = i[95];
  assign o[48949] = i[95];
  assign o[48950] = i[95];
  assign o[48951] = i[95];
  assign o[48952] = i[95];
  assign o[48953] = i[95];
  assign o[48954] = i[95];
  assign o[48955] = i[95];
  assign o[48956] = i[95];
  assign o[48957] = i[95];
  assign o[48958] = i[95];
  assign o[48959] = i[95];
  assign o[48960] = i[95];
  assign o[48961] = i[95];
  assign o[48962] = i[95];
  assign o[48963] = i[95];
  assign o[48964] = i[95];
  assign o[48965] = i[95];
  assign o[48966] = i[95];
  assign o[48967] = i[95];
  assign o[48968] = i[95];
  assign o[48969] = i[95];
  assign o[48970] = i[95];
  assign o[48971] = i[95];
  assign o[48972] = i[95];
  assign o[48973] = i[95];
  assign o[48974] = i[95];
  assign o[48975] = i[95];
  assign o[48976] = i[95];
  assign o[48977] = i[95];
  assign o[48978] = i[95];
  assign o[48979] = i[95];
  assign o[48980] = i[95];
  assign o[48981] = i[95];
  assign o[48982] = i[95];
  assign o[48983] = i[95];
  assign o[48984] = i[95];
  assign o[48985] = i[95];
  assign o[48986] = i[95];
  assign o[48987] = i[95];
  assign o[48988] = i[95];
  assign o[48989] = i[95];
  assign o[48990] = i[95];
  assign o[48991] = i[95];
  assign o[48992] = i[95];
  assign o[48993] = i[95];
  assign o[48994] = i[95];
  assign o[48995] = i[95];
  assign o[48996] = i[95];
  assign o[48997] = i[95];
  assign o[48998] = i[95];
  assign o[48999] = i[95];
  assign o[49000] = i[95];
  assign o[49001] = i[95];
  assign o[49002] = i[95];
  assign o[49003] = i[95];
  assign o[49004] = i[95];
  assign o[49005] = i[95];
  assign o[49006] = i[95];
  assign o[49007] = i[95];
  assign o[49008] = i[95];
  assign o[49009] = i[95];
  assign o[49010] = i[95];
  assign o[49011] = i[95];
  assign o[49012] = i[95];
  assign o[49013] = i[95];
  assign o[49014] = i[95];
  assign o[49015] = i[95];
  assign o[49016] = i[95];
  assign o[49017] = i[95];
  assign o[49018] = i[95];
  assign o[49019] = i[95];
  assign o[49020] = i[95];
  assign o[49021] = i[95];
  assign o[49022] = i[95];
  assign o[49023] = i[95];
  assign o[49024] = i[95];
  assign o[49025] = i[95];
  assign o[49026] = i[95];
  assign o[49027] = i[95];
  assign o[49028] = i[95];
  assign o[49029] = i[95];
  assign o[49030] = i[95];
  assign o[49031] = i[95];
  assign o[49032] = i[95];
  assign o[49033] = i[95];
  assign o[49034] = i[95];
  assign o[49035] = i[95];
  assign o[49036] = i[95];
  assign o[49037] = i[95];
  assign o[49038] = i[95];
  assign o[49039] = i[95];
  assign o[49040] = i[95];
  assign o[49041] = i[95];
  assign o[49042] = i[95];
  assign o[49043] = i[95];
  assign o[49044] = i[95];
  assign o[49045] = i[95];
  assign o[49046] = i[95];
  assign o[49047] = i[95];
  assign o[49048] = i[95];
  assign o[49049] = i[95];
  assign o[49050] = i[95];
  assign o[49051] = i[95];
  assign o[49052] = i[95];
  assign o[49053] = i[95];
  assign o[49054] = i[95];
  assign o[49055] = i[95];
  assign o[49056] = i[95];
  assign o[49057] = i[95];
  assign o[49058] = i[95];
  assign o[49059] = i[95];
  assign o[49060] = i[95];
  assign o[49061] = i[95];
  assign o[49062] = i[95];
  assign o[49063] = i[95];
  assign o[49064] = i[95];
  assign o[49065] = i[95];
  assign o[49066] = i[95];
  assign o[49067] = i[95];
  assign o[49068] = i[95];
  assign o[49069] = i[95];
  assign o[49070] = i[95];
  assign o[49071] = i[95];
  assign o[49072] = i[95];
  assign o[49073] = i[95];
  assign o[49074] = i[95];
  assign o[49075] = i[95];
  assign o[49076] = i[95];
  assign o[49077] = i[95];
  assign o[49078] = i[95];
  assign o[49079] = i[95];
  assign o[49080] = i[95];
  assign o[49081] = i[95];
  assign o[49082] = i[95];
  assign o[49083] = i[95];
  assign o[49084] = i[95];
  assign o[49085] = i[95];
  assign o[49086] = i[95];
  assign o[49087] = i[95];
  assign o[49088] = i[95];
  assign o[49089] = i[95];
  assign o[49090] = i[95];
  assign o[49091] = i[95];
  assign o[49092] = i[95];
  assign o[49093] = i[95];
  assign o[49094] = i[95];
  assign o[49095] = i[95];
  assign o[49096] = i[95];
  assign o[49097] = i[95];
  assign o[49098] = i[95];
  assign o[49099] = i[95];
  assign o[49100] = i[95];
  assign o[49101] = i[95];
  assign o[49102] = i[95];
  assign o[49103] = i[95];
  assign o[49104] = i[95];
  assign o[49105] = i[95];
  assign o[49106] = i[95];
  assign o[49107] = i[95];
  assign o[49108] = i[95];
  assign o[49109] = i[95];
  assign o[49110] = i[95];
  assign o[49111] = i[95];
  assign o[49112] = i[95];
  assign o[49113] = i[95];
  assign o[49114] = i[95];
  assign o[49115] = i[95];
  assign o[49116] = i[95];
  assign o[49117] = i[95];
  assign o[49118] = i[95];
  assign o[49119] = i[95];
  assign o[49120] = i[95];
  assign o[49121] = i[95];
  assign o[49122] = i[95];
  assign o[49123] = i[95];
  assign o[49124] = i[95];
  assign o[49125] = i[95];
  assign o[49126] = i[95];
  assign o[49127] = i[95];
  assign o[49128] = i[95];
  assign o[49129] = i[95];
  assign o[49130] = i[95];
  assign o[49131] = i[95];
  assign o[49132] = i[95];
  assign o[49133] = i[95];
  assign o[49134] = i[95];
  assign o[49135] = i[95];
  assign o[49136] = i[95];
  assign o[49137] = i[95];
  assign o[49138] = i[95];
  assign o[49139] = i[95];
  assign o[49140] = i[95];
  assign o[49141] = i[95];
  assign o[49142] = i[95];
  assign o[49143] = i[95];
  assign o[49144] = i[95];
  assign o[49145] = i[95];
  assign o[49146] = i[95];
  assign o[49147] = i[95];
  assign o[49148] = i[95];
  assign o[49149] = i[95];
  assign o[49150] = i[95];
  assign o[49151] = i[95];
  assign o[48128] = i[94];
  assign o[48129] = i[94];
  assign o[48130] = i[94];
  assign o[48131] = i[94];
  assign o[48132] = i[94];
  assign o[48133] = i[94];
  assign o[48134] = i[94];
  assign o[48135] = i[94];
  assign o[48136] = i[94];
  assign o[48137] = i[94];
  assign o[48138] = i[94];
  assign o[48139] = i[94];
  assign o[48140] = i[94];
  assign o[48141] = i[94];
  assign o[48142] = i[94];
  assign o[48143] = i[94];
  assign o[48144] = i[94];
  assign o[48145] = i[94];
  assign o[48146] = i[94];
  assign o[48147] = i[94];
  assign o[48148] = i[94];
  assign o[48149] = i[94];
  assign o[48150] = i[94];
  assign o[48151] = i[94];
  assign o[48152] = i[94];
  assign o[48153] = i[94];
  assign o[48154] = i[94];
  assign o[48155] = i[94];
  assign o[48156] = i[94];
  assign o[48157] = i[94];
  assign o[48158] = i[94];
  assign o[48159] = i[94];
  assign o[48160] = i[94];
  assign o[48161] = i[94];
  assign o[48162] = i[94];
  assign o[48163] = i[94];
  assign o[48164] = i[94];
  assign o[48165] = i[94];
  assign o[48166] = i[94];
  assign o[48167] = i[94];
  assign o[48168] = i[94];
  assign o[48169] = i[94];
  assign o[48170] = i[94];
  assign o[48171] = i[94];
  assign o[48172] = i[94];
  assign o[48173] = i[94];
  assign o[48174] = i[94];
  assign o[48175] = i[94];
  assign o[48176] = i[94];
  assign o[48177] = i[94];
  assign o[48178] = i[94];
  assign o[48179] = i[94];
  assign o[48180] = i[94];
  assign o[48181] = i[94];
  assign o[48182] = i[94];
  assign o[48183] = i[94];
  assign o[48184] = i[94];
  assign o[48185] = i[94];
  assign o[48186] = i[94];
  assign o[48187] = i[94];
  assign o[48188] = i[94];
  assign o[48189] = i[94];
  assign o[48190] = i[94];
  assign o[48191] = i[94];
  assign o[48192] = i[94];
  assign o[48193] = i[94];
  assign o[48194] = i[94];
  assign o[48195] = i[94];
  assign o[48196] = i[94];
  assign o[48197] = i[94];
  assign o[48198] = i[94];
  assign o[48199] = i[94];
  assign o[48200] = i[94];
  assign o[48201] = i[94];
  assign o[48202] = i[94];
  assign o[48203] = i[94];
  assign o[48204] = i[94];
  assign o[48205] = i[94];
  assign o[48206] = i[94];
  assign o[48207] = i[94];
  assign o[48208] = i[94];
  assign o[48209] = i[94];
  assign o[48210] = i[94];
  assign o[48211] = i[94];
  assign o[48212] = i[94];
  assign o[48213] = i[94];
  assign o[48214] = i[94];
  assign o[48215] = i[94];
  assign o[48216] = i[94];
  assign o[48217] = i[94];
  assign o[48218] = i[94];
  assign o[48219] = i[94];
  assign o[48220] = i[94];
  assign o[48221] = i[94];
  assign o[48222] = i[94];
  assign o[48223] = i[94];
  assign o[48224] = i[94];
  assign o[48225] = i[94];
  assign o[48226] = i[94];
  assign o[48227] = i[94];
  assign o[48228] = i[94];
  assign o[48229] = i[94];
  assign o[48230] = i[94];
  assign o[48231] = i[94];
  assign o[48232] = i[94];
  assign o[48233] = i[94];
  assign o[48234] = i[94];
  assign o[48235] = i[94];
  assign o[48236] = i[94];
  assign o[48237] = i[94];
  assign o[48238] = i[94];
  assign o[48239] = i[94];
  assign o[48240] = i[94];
  assign o[48241] = i[94];
  assign o[48242] = i[94];
  assign o[48243] = i[94];
  assign o[48244] = i[94];
  assign o[48245] = i[94];
  assign o[48246] = i[94];
  assign o[48247] = i[94];
  assign o[48248] = i[94];
  assign o[48249] = i[94];
  assign o[48250] = i[94];
  assign o[48251] = i[94];
  assign o[48252] = i[94];
  assign o[48253] = i[94];
  assign o[48254] = i[94];
  assign o[48255] = i[94];
  assign o[48256] = i[94];
  assign o[48257] = i[94];
  assign o[48258] = i[94];
  assign o[48259] = i[94];
  assign o[48260] = i[94];
  assign o[48261] = i[94];
  assign o[48262] = i[94];
  assign o[48263] = i[94];
  assign o[48264] = i[94];
  assign o[48265] = i[94];
  assign o[48266] = i[94];
  assign o[48267] = i[94];
  assign o[48268] = i[94];
  assign o[48269] = i[94];
  assign o[48270] = i[94];
  assign o[48271] = i[94];
  assign o[48272] = i[94];
  assign o[48273] = i[94];
  assign o[48274] = i[94];
  assign o[48275] = i[94];
  assign o[48276] = i[94];
  assign o[48277] = i[94];
  assign o[48278] = i[94];
  assign o[48279] = i[94];
  assign o[48280] = i[94];
  assign o[48281] = i[94];
  assign o[48282] = i[94];
  assign o[48283] = i[94];
  assign o[48284] = i[94];
  assign o[48285] = i[94];
  assign o[48286] = i[94];
  assign o[48287] = i[94];
  assign o[48288] = i[94];
  assign o[48289] = i[94];
  assign o[48290] = i[94];
  assign o[48291] = i[94];
  assign o[48292] = i[94];
  assign o[48293] = i[94];
  assign o[48294] = i[94];
  assign o[48295] = i[94];
  assign o[48296] = i[94];
  assign o[48297] = i[94];
  assign o[48298] = i[94];
  assign o[48299] = i[94];
  assign o[48300] = i[94];
  assign o[48301] = i[94];
  assign o[48302] = i[94];
  assign o[48303] = i[94];
  assign o[48304] = i[94];
  assign o[48305] = i[94];
  assign o[48306] = i[94];
  assign o[48307] = i[94];
  assign o[48308] = i[94];
  assign o[48309] = i[94];
  assign o[48310] = i[94];
  assign o[48311] = i[94];
  assign o[48312] = i[94];
  assign o[48313] = i[94];
  assign o[48314] = i[94];
  assign o[48315] = i[94];
  assign o[48316] = i[94];
  assign o[48317] = i[94];
  assign o[48318] = i[94];
  assign o[48319] = i[94];
  assign o[48320] = i[94];
  assign o[48321] = i[94];
  assign o[48322] = i[94];
  assign o[48323] = i[94];
  assign o[48324] = i[94];
  assign o[48325] = i[94];
  assign o[48326] = i[94];
  assign o[48327] = i[94];
  assign o[48328] = i[94];
  assign o[48329] = i[94];
  assign o[48330] = i[94];
  assign o[48331] = i[94];
  assign o[48332] = i[94];
  assign o[48333] = i[94];
  assign o[48334] = i[94];
  assign o[48335] = i[94];
  assign o[48336] = i[94];
  assign o[48337] = i[94];
  assign o[48338] = i[94];
  assign o[48339] = i[94];
  assign o[48340] = i[94];
  assign o[48341] = i[94];
  assign o[48342] = i[94];
  assign o[48343] = i[94];
  assign o[48344] = i[94];
  assign o[48345] = i[94];
  assign o[48346] = i[94];
  assign o[48347] = i[94];
  assign o[48348] = i[94];
  assign o[48349] = i[94];
  assign o[48350] = i[94];
  assign o[48351] = i[94];
  assign o[48352] = i[94];
  assign o[48353] = i[94];
  assign o[48354] = i[94];
  assign o[48355] = i[94];
  assign o[48356] = i[94];
  assign o[48357] = i[94];
  assign o[48358] = i[94];
  assign o[48359] = i[94];
  assign o[48360] = i[94];
  assign o[48361] = i[94];
  assign o[48362] = i[94];
  assign o[48363] = i[94];
  assign o[48364] = i[94];
  assign o[48365] = i[94];
  assign o[48366] = i[94];
  assign o[48367] = i[94];
  assign o[48368] = i[94];
  assign o[48369] = i[94];
  assign o[48370] = i[94];
  assign o[48371] = i[94];
  assign o[48372] = i[94];
  assign o[48373] = i[94];
  assign o[48374] = i[94];
  assign o[48375] = i[94];
  assign o[48376] = i[94];
  assign o[48377] = i[94];
  assign o[48378] = i[94];
  assign o[48379] = i[94];
  assign o[48380] = i[94];
  assign o[48381] = i[94];
  assign o[48382] = i[94];
  assign o[48383] = i[94];
  assign o[48384] = i[94];
  assign o[48385] = i[94];
  assign o[48386] = i[94];
  assign o[48387] = i[94];
  assign o[48388] = i[94];
  assign o[48389] = i[94];
  assign o[48390] = i[94];
  assign o[48391] = i[94];
  assign o[48392] = i[94];
  assign o[48393] = i[94];
  assign o[48394] = i[94];
  assign o[48395] = i[94];
  assign o[48396] = i[94];
  assign o[48397] = i[94];
  assign o[48398] = i[94];
  assign o[48399] = i[94];
  assign o[48400] = i[94];
  assign o[48401] = i[94];
  assign o[48402] = i[94];
  assign o[48403] = i[94];
  assign o[48404] = i[94];
  assign o[48405] = i[94];
  assign o[48406] = i[94];
  assign o[48407] = i[94];
  assign o[48408] = i[94];
  assign o[48409] = i[94];
  assign o[48410] = i[94];
  assign o[48411] = i[94];
  assign o[48412] = i[94];
  assign o[48413] = i[94];
  assign o[48414] = i[94];
  assign o[48415] = i[94];
  assign o[48416] = i[94];
  assign o[48417] = i[94];
  assign o[48418] = i[94];
  assign o[48419] = i[94];
  assign o[48420] = i[94];
  assign o[48421] = i[94];
  assign o[48422] = i[94];
  assign o[48423] = i[94];
  assign o[48424] = i[94];
  assign o[48425] = i[94];
  assign o[48426] = i[94];
  assign o[48427] = i[94];
  assign o[48428] = i[94];
  assign o[48429] = i[94];
  assign o[48430] = i[94];
  assign o[48431] = i[94];
  assign o[48432] = i[94];
  assign o[48433] = i[94];
  assign o[48434] = i[94];
  assign o[48435] = i[94];
  assign o[48436] = i[94];
  assign o[48437] = i[94];
  assign o[48438] = i[94];
  assign o[48439] = i[94];
  assign o[48440] = i[94];
  assign o[48441] = i[94];
  assign o[48442] = i[94];
  assign o[48443] = i[94];
  assign o[48444] = i[94];
  assign o[48445] = i[94];
  assign o[48446] = i[94];
  assign o[48447] = i[94];
  assign o[48448] = i[94];
  assign o[48449] = i[94];
  assign o[48450] = i[94];
  assign o[48451] = i[94];
  assign o[48452] = i[94];
  assign o[48453] = i[94];
  assign o[48454] = i[94];
  assign o[48455] = i[94];
  assign o[48456] = i[94];
  assign o[48457] = i[94];
  assign o[48458] = i[94];
  assign o[48459] = i[94];
  assign o[48460] = i[94];
  assign o[48461] = i[94];
  assign o[48462] = i[94];
  assign o[48463] = i[94];
  assign o[48464] = i[94];
  assign o[48465] = i[94];
  assign o[48466] = i[94];
  assign o[48467] = i[94];
  assign o[48468] = i[94];
  assign o[48469] = i[94];
  assign o[48470] = i[94];
  assign o[48471] = i[94];
  assign o[48472] = i[94];
  assign o[48473] = i[94];
  assign o[48474] = i[94];
  assign o[48475] = i[94];
  assign o[48476] = i[94];
  assign o[48477] = i[94];
  assign o[48478] = i[94];
  assign o[48479] = i[94];
  assign o[48480] = i[94];
  assign o[48481] = i[94];
  assign o[48482] = i[94];
  assign o[48483] = i[94];
  assign o[48484] = i[94];
  assign o[48485] = i[94];
  assign o[48486] = i[94];
  assign o[48487] = i[94];
  assign o[48488] = i[94];
  assign o[48489] = i[94];
  assign o[48490] = i[94];
  assign o[48491] = i[94];
  assign o[48492] = i[94];
  assign o[48493] = i[94];
  assign o[48494] = i[94];
  assign o[48495] = i[94];
  assign o[48496] = i[94];
  assign o[48497] = i[94];
  assign o[48498] = i[94];
  assign o[48499] = i[94];
  assign o[48500] = i[94];
  assign o[48501] = i[94];
  assign o[48502] = i[94];
  assign o[48503] = i[94];
  assign o[48504] = i[94];
  assign o[48505] = i[94];
  assign o[48506] = i[94];
  assign o[48507] = i[94];
  assign o[48508] = i[94];
  assign o[48509] = i[94];
  assign o[48510] = i[94];
  assign o[48511] = i[94];
  assign o[48512] = i[94];
  assign o[48513] = i[94];
  assign o[48514] = i[94];
  assign o[48515] = i[94];
  assign o[48516] = i[94];
  assign o[48517] = i[94];
  assign o[48518] = i[94];
  assign o[48519] = i[94];
  assign o[48520] = i[94];
  assign o[48521] = i[94];
  assign o[48522] = i[94];
  assign o[48523] = i[94];
  assign o[48524] = i[94];
  assign o[48525] = i[94];
  assign o[48526] = i[94];
  assign o[48527] = i[94];
  assign o[48528] = i[94];
  assign o[48529] = i[94];
  assign o[48530] = i[94];
  assign o[48531] = i[94];
  assign o[48532] = i[94];
  assign o[48533] = i[94];
  assign o[48534] = i[94];
  assign o[48535] = i[94];
  assign o[48536] = i[94];
  assign o[48537] = i[94];
  assign o[48538] = i[94];
  assign o[48539] = i[94];
  assign o[48540] = i[94];
  assign o[48541] = i[94];
  assign o[48542] = i[94];
  assign o[48543] = i[94];
  assign o[48544] = i[94];
  assign o[48545] = i[94];
  assign o[48546] = i[94];
  assign o[48547] = i[94];
  assign o[48548] = i[94];
  assign o[48549] = i[94];
  assign o[48550] = i[94];
  assign o[48551] = i[94];
  assign o[48552] = i[94];
  assign o[48553] = i[94];
  assign o[48554] = i[94];
  assign o[48555] = i[94];
  assign o[48556] = i[94];
  assign o[48557] = i[94];
  assign o[48558] = i[94];
  assign o[48559] = i[94];
  assign o[48560] = i[94];
  assign o[48561] = i[94];
  assign o[48562] = i[94];
  assign o[48563] = i[94];
  assign o[48564] = i[94];
  assign o[48565] = i[94];
  assign o[48566] = i[94];
  assign o[48567] = i[94];
  assign o[48568] = i[94];
  assign o[48569] = i[94];
  assign o[48570] = i[94];
  assign o[48571] = i[94];
  assign o[48572] = i[94];
  assign o[48573] = i[94];
  assign o[48574] = i[94];
  assign o[48575] = i[94];
  assign o[48576] = i[94];
  assign o[48577] = i[94];
  assign o[48578] = i[94];
  assign o[48579] = i[94];
  assign o[48580] = i[94];
  assign o[48581] = i[94];
  assign o[48582] = i[94];
  assign o[48583] = i[94];
  assign o[48584] = i[94];
  assign o[48585] = i[94];
  assign o[48586] = i[94];
  assign o[48587] = i[94];
  assign o[48588] = i[94];
  assign o[48589] = i[94];
  assign o[48590] = i[94];
  assign o[48591] = i[94];
  assign o[48592] = i[94];
  assign o[48593] = i[94];
  assign o[48594] = i[94];
  assign o[48595] = i[94];
  assign o[48596] = i[94];
  assign o[48597] = i[94];
  assign o[48598] = i[94];
  assign o[48599] = i[94];
  assign o[48600] = i[94];
  assign o[48601] = i[94];
  assign o[48602] = i[94];
  assign o[48603] = i[94];
  assign o[48604] = i[94];
  assign o[48605] = i[94];
  assign o[48606] = i[94];
  assign o[48607] = i[94];
  assign o[48608] = i[94];
  assign o[48609] = i[94];
  assign o[48610] = i[94];
  assign o[48611] = i[94];
  assign o[48612] = i[94];
  assign o[48613] = i[94];
  assign o[48614] = i[94];
  assign o[48615] = i[94];
  assign o[48616] = i[94];
  assign o[48617] = i[94];
  assign o[48618] = i[94];
  assign o[48619] = i[94];
  assign o[48620] = i[94];
  assign o[48621] = i[94];
  assign o[48622] = i[94];
  assign o[48623] = i[94];
  assign o[48624] = i[94];
  assign o[48625] = i[94];
  assign o[48626] = i[94];
  assign o[48627] = i[94];
  assign o[48628] = i[94];
  assign o[48629] = i[94];
  assign o[48630] = i[94];
  assign o[48631] = i[94];
  assign o[48632] = i[94];
  assign o[48633] = i[94];
  assign o[48634] = i[94];
  assign o[48635] = i[94];
  assign o[48636] = i[94];
  assign o[48637] = i[94];
  assign o[48638] = i[94];
  assign o[48639] = i[94];
  assign o[47616] = i[93];
  assign o[47617] = i[93];
  assign o[47618] = i[93];
  assign o[47619] = i[93];
  assign o[47620] = i[93];
  assign o[47621] = i[93];
  assign o[47622] = i[93];
  assign o[47623] = i[93];
  assign o[47624] = i[93];
  assign o[47625] = i[93];
  assign o[47626] = i[93];
  assign o[47627] = i[93];
  assign o[47628] = i[93];
  assign o[47629] = i[93];
  assign o[47630] = i[93];
  assign o[47631] = i[93];
  assign o[47632] = i[93];
  assign o[47633] = i[93];
  assign o[47634] = i[93];
  assign o[47635] = i[93];
  assign o[47636] = i[93];
  assign o[47637] = i[93];
  assign o[47638] = i[93];
  assign o[47639] = i[93];
  assign o[47640] = i[93];
  assign o[47641] = i[93];
  assign o[47642] = i[93];
  assign o[47643] = i[93];
  assign o[47644] = i[93];
  assign o[47645] = i[93];
  assign o[47646] = i[93];
  assign o[47647] = i[93];
  assign o[47648] = i[93];
  assign o[47649] = i[93];
  assign o[47650] = i[93];
  assign o[47651] = i[93];
  assign o[47652] = i[93];
  assign o[47653] = i[93];
  assign o[47654] = i[93];
  assign o[47655] = i[93];
  assign o[47656] = i[93];
  assign o[47657] = i[93];
  assign o[47658] = i[93];
  assign o[47659] = i[93];
  assign o[47660] = i[93];
  assign o[47661] = i[93];
  assign o[47662] = i[93];
  assign o[47663] = i[93];
  assign o[47664] = i[93];
  assign o[47665] = i[93];
  assign o[47666] = i[93];
  assign o[47667] = i[93];
  assign o[47668] = i[93];
  assign o[47669] = i[93];
  assign o[47670] = i[93];
  assign o[47671] = i[93];
  assign o[47672] = i[93];
  assign o[47673] = i[93];
  assign o[47674] = i[93];
  assign o[47675] = i[93];
  assign o[47676] = i[93];
  assign o[47677] = i[93];
  assign o[47678] = i[93];
  assign o[47679] = i[93];
  assign o[47680] = i[93];
  assign o[47681] = i[93];
  assign o[47682] = i[93];
  assign o[47683] = i[93];
  assign o[47684] = i[93];
  assign o[47685] = i[93];
  assign o[47686] = i[93];
  assign o[47687] = i[93];
  assign o[47688] = i[93];
  assign o[47689] = i[93];
  assign o[47690] = i[93];
  assign o[47691] = i[93];
  assign o[47692] = i[93];
  assign o[47693] = i[93];
  assign o[47694] = i[93];
  assign o[47695] = i[93];
  assign o[47696] = i[93];
  assign o[47697] = i[93];
  assign o[47698] = i[93];
  assign o[47699] = i[93];
  assign o[47700] = i[93];
  assign o[47701] = i[93];
  assign o[47702] = i[93];
  assign o[47703] = i[93];
  assign o[47704] = i[93];
  assign o[47705] = i[93];
  assign o[47706] = i[93];
  assign o[47707] = i[93];
  assign o[47708] = i[93];
  assign o[47709] = i[93];
  assign o[47710] = i[93];
  assign o[47711] = i[93];
  assign o[47712] = i[93];
  assign o[47713] = i[93];
  assign o[47714] = i[93];
  assign o[47715] = i[93];
  assign o[47716] = i[93];
  assign o[47717] = i[93];
  assign o[47718] = i[93];
  assign o[47719] = i[93];
  assign o[47720] = i[93];
  assign o[47721] = i[93];
  assign o[47722] = i[93];
  assign o[47723] = i[93];
  assign o[47724] = i[93];
  assign o[47725] = i[93];
  assign o[47726] = i[93];
  assign o[47727] = i[93];
  assign o[47728] = i[93];
  assign o[47729] = i[93];
  assign o[47730] = i[93];
  assign o[47731] = i[93];
  assign o[47732] = i[93];
  assign o[47733] = i[93];
  assign o[47734] = i[93];
  assign o[47735] = i[93];
  assign o[47736] = i[93];
  assign o[47737] = i[93];
  assign o[47738] = i[93];
  assign o[47739] = i[93];
  assign o[47740] = i[93];
  assign o[47741] = i[93];
  assign o[47742] = i[93];
  assign o[47743] = i[93];
  assign o[47744] = i[93];
  assign o[47745] = i[93];
  assign o[47746] = i[93];
  assign o[47747] = i[93];
  assign o[47748] = i[93];
  assign o[47749] = i[93];
  assign o[47750] = i[93];
  assign o[47751] = i[93];
  assign o[47752] = i[93];
  assign o[47753] = i[93];
  assign o[47754] = i[93];
  assign o[47755] = i[93];
  assign o[47756] = i[93];
  assign o[47757] = i[93];
  assign o[47758] = i[93];
  assign o[47759] = i[93];
  assign o[47760] = i[93];
  assign o[47761] = i[93];
  assign o[47762] = i[93];
  assign o[47763] = i[93];
  assign o[47764] = i[93];
  assign o[47765] = i[93];
  assign o[47766] = i[93];
  assign o[47767] = i[93];
  assign o[47768] = i[93];
  assign o[47769] = i[93];
  assign o[47770] = i[93];
  assign o[47771] = i[93];
  assign o[47772] = i[93];
  assign o[47773] = i[93];
  assign o[47774] = i[93];
  assign o[47775] = i[93];
  assign o[47776] = i[93];
  assign o[47777] = i[93];
  assign o[47778] = i[93];
  assign o[47779] = i[93];
  assign o[47780] = i[93];
  assign o[47781] = i[93];
  assign o[47782] = i[93];
  assign o[47783] = i[93];
  assign o[47784] = i[93];
  assign o[47785] = i[93];
  assign o[47786] = i[93];
  assign o[47787] = i[93];
  assign o[47788] = i[93];
  assign o[47789] = i[93];
  assign o[47790] = i[93];
  assign o[47791] = i[93];
  assign o[47792] = i[93];
  assign o[47793] = i[93];
  assign o[47794] = i[93];
  assign o[47795] = i[93];
  assign o[47796] = i[93];
  assign o[47797] = i[93];
  assign o[47798] = i[93];
  assign o[47799] = i[93];
  assign o[47800] = i[93];
  assign o[47801] = i[93];
  assign o[47802] = i[93];
  assign o[47803] = i[93];
  assign o[47804] = i[93];
  assign o[47805] = i[93];
  assign o[47806] = i[93];
  assign o[47807] = i[93];
  assign o[47808] = i[93];
  assign o[47809] = i[93];
  assign o[47810] = i[93];
  assign o[47811] = i[93];
  assign o[47812] = i[93];
  assign o[47813] = i[93];
  assign o[47814] = i[93];
  assign o[47815] = i[93];
  assign o[47816] = i[93];
  assign o[47817] = i[93];
  assign o[47818] = i[93];
  assign o[47819] = i[93];
  assign o[47820] = i[93];
  assign o[47821] = i[93];
  assign o[47822] = i[93];
  assign o[47823] = i[93];
  assign o[47824] = i[93];
  assign o[47825] = i[93];
  assign o[47826] = i[93];
  assign o[47827] = i[93];
  assign o[47828] = i[93];
  assign o[47829] = i[93];
  assign o[47830] = i[93];
  assign o[47831] = i[93];
  assign o[47832] = i[93];
  assign o[47833] = i[93];
  assign o[47834] = i[93];
  assign o[47835] = i[93];
  assign o[47836] = i[93];
  assign o[47837] = i[93];
  assign o[47838] = i[93];
  assign o[47839] = i[93];
  assign o[47840] = i[93];
  assign o[47841] = i[93];
  assign o[47842] = i[93];
  assign o[47843] = i[93];
  assign o[47844] = i[93];
  assign o[47845] = i[93];
  assign o[47846] = i[93];
  assign o[47847] = i[93];
  assign o[47848] = i[93];
  assign o[47849] = i[93];
  assign o[47850] = i[93];
  assign o[47851] = i[93];
  assign o[47852] = i[93];
  assign o[47853] = i[93];
  assign o[47854] = i[93];
  assign o[47855] = i[93];
  assign o[47856] = i[93];
  assign o[47857] = i[93];
  assign o[47858] = i[93];
  assign o[47859] = i[93];
  assign o[47860] = i[93];
  assign o[47861] = i[93];
  assign o[47862] = i[93];
  assign o[47863] = i[93];
  assign o[47864] = i[93];
  assign o[47865] = i[93];
  assign o[47866] = i[93];
  assign o[47867] = i[93];
  assign o[47868] = i[93];
  assign o[47869] = i[93];
  assign o[47870] = i[93];
  assign o[47871] = i[93];
  assign o[47872] = i[93];
  assign o[47873] = i[93];
  assign o[47874] = i[93];
  assign o[47875] = i[93];
  assign o[47876] = i[93];
  assign o[47877] = i[93];
  assign o[47878] = i[93];
  assign o[47879] = i[93];
  assign o[47880] = i[93];
  assign o[47881] = i[93];
  assign o[47882] = i[93];
  assign o[47883] = i[93];
  assign o[47884] = i[93];
  assign o[47885] = i[93];
  assign o[47886] = i[93];
  assign o[47887] = i[93];
  assign o[47888] = i[93];
  assign o[47889] = i[93];
  assign o[47890] = i[93];
  assign o[47891] = i[93];
  assign o[47892] = i[93];
  assign o[47893] = i[93];
  assign o[47894] = i[93];
  assign o[47895] = i[93];
  assign o[47896] = i[93];
  assign o[47897] = i[93];
  assign o[47898] = i[93];
  assign o[47899] = i[93];
  assign o[47900] = i[93];
  assign o[47901] = i[93];
  assign o[47902] = i[93];
  assign o[47903] = i[93];
  assign o[47904] = i[93];
  assign o[47905] = i[93];
  assign o[47906] = i[93];
  assign o[47907] = i[93];
  assign o[47908] = i[93];
  assign o[47909] = i[93];
  assign o[47910] = i[93];
  assign o[47911] = i[93];
  assign o[47912] = i[93];
  assign o[47913] = i[93];
  assign o[47914] = i[93];
  assign o[47915] = i[93];
  assign o[47916] = i[93];
  assign o[47917] = i[93];
  assign o[47918] = i[93];
  assign o[47919] = i[93];
  assign o[47920] = i[93];
  assign o[47921] = i[93];
  assign o[47922] = i[93];
  assign o[47923] = i[93];
  assign o[47924] = i[93];
  assign o[47925] = i[93];
  assign o[47926] = i[93];
  assign o[47927] = i[93];
  assign o[47928] = i[93];
  assign o[47929] = i[93];
  assign o[47930] = i[93];
  assign o[47931] = i[93];
  assign o[47932] = i[93];
  assign o[47933] = i[93];
  assign o[47934] = i[93];
  assign o[47935] = i[93];
  assign o[47936] = i[93];
  assign o[47937] = i[93];
  assign o[47938] = i[93];
  assign o[47939] = i[93];
  assign o[47940] = i[93];
  assign o[47941] = i[93];
  assign o[47942] = i[93];
  assign o[47943] = i[93];
  assign o[47944] = i[93];
  assign o[47945] = i[93];
  assign o[47946] = i[93];
  assign o[47947] = i[93];
  assign o[47948] = i[93];
  assign o[47949] = i[93];
  assign o[47950] = i[93];
  assign o[47951] = i[93];
  assign o[47952] = i[93];
  assign o[47953] = i[93];
  assign o[47954] = i[93];
  assign o[47955] = i[93];
  assign o[47956] = i[93];
  assign o[47957] = i[93];
  assign o[47958] = i[93];
  assign o[47959] = i[93];
  assign o[47960] = i[93];
  assign o[47961] = i[93];
  assign o[47962] = i[93];
  assign o[47963] = i[93];
  assign o[47964] = i[93];
  assign o[47965] = i[93];
  assign o[47966] = i[93];
  assign o[47967] = i[93];
  assign o[47968] = i[93];
  assign o[47969] = i[93];
  assign o[47970] = i[93];
  assign o[47971] = i[93];
  assign o[47972] = i[93];
  assign o[47973] = i[93];
  assign o[47974] = i[93];
  assign o[47975] = i[93];
  assign o[47976] = i[93];
  assign o[47977] = i[93];
  assign o[47978] = i[93];
  assign o[47979] = i[93];
  assign o[47980] = i[93];
  assign o[47981] = i[93];
  assign o[47982] = i[93];
  assign o[47983] = i[93];
  assign o[47984] = i[93];
  assign o[47985] = i[93];
  assign o[47986] = i[93];
  assign o[47987] = i[93];
  assign o[47988] = i[93];
  assign o[47989] = i[93];
  assign o[47990] = i[93];
  assign o[47991] = i[93];
  assign o[47992] = i[93];
  assign o[47993] = i[93];
  assign o[47994] = i[93];
  assign o[47995] = i[93];
  assign o[47996] = i[93];
  assign o[47997] = i[93];
  assign o[47998] = i[93];
  assign o[47999] = i[93];
  assign o[48000] = i[93];
  assign o[48001] = i[93];
  assign o[48002] = i[93];
  assign o[48003] = i[93];
  assign o[48004] = i[93];
  assign o[48005] = i[93];
  assign o[48006] = i[93];
  assign o[48007] = i[93];
  assign o[48008] = i[93];
  assign o[48009] = i[93];
  assign o[48010] = i[93];
  assign o[48011] = i[93];
  assign o[48012] = i[93];
  assign o[48013] = i[93];
  assign o[48014] = i[93];
  assign o[48015] = i[93];
  assign o[48016] = i[93];
  assign o[48017] = i[93];
  assign o[48018] = i[93];
  assign o[48019] = i[93];
  assign o[48020] = i[93];
  assign o[48021] = i[93];
  assign o[48022] = i[93];
  assign o[48023] = i[93];
  assign o[48024] = i[93];
  assign o[48025] = i[93];
  assign o[48026] = i[93];
  assign o[48027] = i[93];
  assign o[48028] = i[93];
  assign o[48029] = i[93];
  assign o[48030] = i[93];
  assign o[48031] = i[93];
  assign o[48032] = i[93];
  assign o[48033] = i[93];
  assign o[48034] = i[93];
  assign o[48035] = i[93];
  assign o[48036] = i[93];
  assign o[48037] = i[93];
  assign o[48038] = i[93];
  assign o[48039] = i[93];
  assign o[48040] = i[93];
  assign o[48041] = i[93];
  assign o[48042] = i[93];
  assign o[48043] = i[93];
  assign o[48044] = i[93];
  assign o[48045] = i[93];
  assign o[48046] = i[93];
  assign o[48047] = i[93];
  assign o[48048] = i[93];
  assign o[48049] = i[93];
  assign o[48050] = i[93];
  assign o[48051] = i[93];
  assign o[48052] = i[93];
  assign o[48053] = i[93];
  assign o[48054] = i[93];
  assign o[48055] = i[93];
  assign o[48056] = i[93];
  assign o[48057] = i[93];
  assign o[48058] = i[93];
  assign o[48059] = i[93];
  assign o[48060] = i[93];
  assign o[48061] = i[93];
  assign o[48062] = i[93];
  assign o[48063] = i[93];
  assign o[48064] = i[93];
  assign o[48065] = i[93];
  assign o[48066] = i[93];
  assign o[48067] = i[93];
  assign o[48068] = i[93];
  assign o[48069] = i[93];
  assign o[48070] = i[93];
  assign o[48071] = i[93];
  assign o[48072] = i[93];
  assign o[48073] = i[93];
  assign o[48074] = i[93];
  assign o[48075] = i[93];
  assign o[48076] = i[93];
  assign o[48077] = i[93];
  assign o[48078] = i[93];
  assign o[48079] = i[93];
  assign o[48080] = i[93];
  assign o[48081] = i[93];
  assign o[48082] = i[93];
  assign o[48083] = i[93];
  assign o[48084] = i[93];
  assign o[48085] = i[93];
  assign o[48086] = i[93];
  assign o[48087] = i[93];
  assign o[48088] = i[93];
  assign o[48089] = i[93];
  assign o[48090] = i[93];
  assign o[48091] = i[93];
  assign o[48092] = i[93];
  assign o[48093] = i[93];
  assign o[48094] = i[93];
  assign o[48095] = i[93];
  assign o[48096] = i[93];
  assign o[48097] = i[93];
  assign o[48098] = i[93];
  assign o[48099] = i[93];
  assign o[48100] = i[93];
  assign o[48101] = i[93];
  assign o[48102] = i[93];
  assign o[48103] = i[93];
  assign o[48104] = i[93];
  assign o[48105] = i[93];
  assign o[48106] = i[93];
  assign o[48107] = i[93];
  assign o[48108] = i[93];
  assign o[48109] = i[93];
  assign o[48110] = i[93];
  assign o[48111] = i[93];
  assign o[48112] = i[93];
  assign o[48113] = i[93];
  assign o[48114] = i[93];
  assign o[48115] = i[93];
  assign o[48116] = i[93];
  assign o[48117] = i[93];
  assign o[48118] = i[93];
  assign o[48119] = i[93];
  assign o[48120] = i[93];
  assign o[48121] = i[93];
  assign o[48122] = i[93];
  assign o[48123] = i[93];
  assign o[48124] = i[93];
  assign o[48125] = i[93];
  assign o[48126] = i[93];
  assign o[48127] = i[93];
  assign o[47104] = i[92];
  assign o[47105] = i[92];
  assign o[47106] = i[92];
  assign o[47107] = i[92];
  assign o[47108] = i[92];
  assign o[47109] = i[92];
  assign o[47110] = i[92];
  assign o[47111] = i[92];
  assign o[47112] = i[92];
  assign o[47113] = i[92];
  assign o[47114] = i[92];
  assign o[47115] = i[92];
  assign o[47116] = i[92];
  assign o[47117] = i[92];
  assign o[47118] = i[92];
  assign o[47119] = i[92];
  assign o[47120] = i[92];
  assign o[47121] = i[92];
  assign o[47122] = i[92];
  assign o[47123] = i[92];
  assign o[47124] = i[92];
  assign o[47125] = i[92];
  assign o[47126] = i[92];
  assign o[47127] = i[92];
  assign o[47128] = i[92];
  assign o[47129] = i[92];
  assign o[47130] = i[92];
  assign o[47131] = i[92];
  assign o[47132] = i[92];
  assign o[47133] = i[92];
  assign o[47134] = i[92];
  assign o[47135] = i[92];
  assign o[47136] = i[92];
  assign o[47137] = i[92];
  assign o[47138] = i[92];
  assign o[47139] = i[92];
  assign o[47140] = i[92];
  assign o[47141] = i[92];
  assign o[47142] = i[92];
  assign o[47143] = i[92];
  assign o[47144] = i[92];
  assign o[47145] = i[92];
  assign o[47146] = i[92];
  assign o[47147] = i[92];
  assign o[47148] = i[92];
  assign o[47149] = i[92];
  assign o[47150] = i[92];
  assign o[47151] = i[92];
  assign o[47152] = i[92];
  assign o[47153] = i[92];
  assign o[47154] = i[92];
  assign o[47155] = i[92];
  assign o[47156] = i[92];
  assign o[47157] = i[92];
  assign o[47158] = i[92];
  assign o[47159] = i[92];
  assign o[47160] = i[92];
  assign o[47161] = i[92];
  assign o[47162] = i[92];
  assign o[47163] = i[92];
  assign o[47164] = i[92];
  assign o[47165] = i[92];
  assign o[47166] = i[92];
  assign o[47167] = i[92];
  assign o[47168] = i[92];
  assign o[47169] = i[92];
  assign o[47170] = i[92];
  assign o[47171] = i[92];
  assign o[47172] = i[92];
  assign o[47173] = i[92];
  assign o[47174] = i[92];
  assign o[47175] = i[92];
  assign o[47176] = i[92];
  assign o[47177] = i[92];
  assign o[47178] = i[92];
  assign o[47179] = i[92];
  assign o[47180] = i[92];
  assign o[47181] = i[92];
  assign o[47182] = i[92];
  assign o[47183] = i[92];
  assign o[47184] = i[92];
  assign o[47185] = i[92];
  assign o[47186] = i[92];
  assign o[47187] = i[92];
  assign o[47188] = i[92];
  assign o[47189] = i[92];
  assign o[47190] = i[92];
  assign o[47191] = i[92];
  assign o[47192] = i[92];
  assign o[47193] = i[92];
  assign o[47194] = i[92];
  assign o[47195] = i[92];
  assign o[47196] = i[92];
  assign o[47197] = i[92];
  assign o[47198] = i[92];
  assign o[47199] = i[92];
  assign o[47200] = i[92];
  assign o[47201] = i[92];
  assign o[47202] = i[92];
  assign o[47203] = i[92];
  assign o[47204] = i[92];
  assign o[47205] = i[92];
  assign o[47206] = i[92];
  assign o[47207] = i[92];
  assign o[47208] = i[92];
  assign o[47209] = i[92];
  assign o[47210] = i[92];
  assign o[47211] = i[92];
  assign o[47212] = i[92];
  assign o[47213] = i[92];
  assign o[47214] = i[92];
  assign o[47215] = i[92];
  assign o[47216] = i[92];
  assign o[47217] = i[92];
  assign o[47218] = i[92];
  assign o[47219] = i[92];
  assign o[47220] = i[92];
  assign o[47221] = i[92];
  assign o[47222] = i[92];
  assign o[47223] = i[92];
  assign o[47224] = i[92];
  assign o[47225] = i[92];
  assign o[47226] = i[92];
  assign o[47227] = i[92];
  assign o[47228] = i[92];
  assign o[47229] = i[92];
  assign o[47230] = i[92];
  assign o[47231] = i[92];
  assign o[47232] = i[92];
  assign o[47233] = i[92];
  assign o[47234] = i[92];
  assign o[47235] = i[92];
  assign o[47236] = i[92];
  assign o[47237] = i[92];
  assign o[47238] = i[92];
  assign o[47239] = i[92];
  assign o[47240] = i[92];
  assign o[47241] = i[92];
  assign o[47242] = i[92];
  assign o[47243] = i[92];
  assign o[47244] = i[92];
  assign o[47245] = i[92];
  assign o[47246] = i[92];
  assign o[47247] = i[92];
  assign o[47248] = i[92];
  assign o[47249] = i[92];
  assign o[47250] = i[92];
  assign o[47251] = i[92];
  assign o[47252] = i[92];
  assign o[47253] = i[92];
  assign o[47254] = i[92];
  assign o[47255] = i[92];
  assign o[47256] = i[92];
  assign o[47257] = i[92];
  assign o[47258] = i[92];
  assign o[47259] = i[92];
  assign o[47260] = i[92];
  assign o[47261] = i[92];
  assign o[47262] = i[92];
  assign o[47263] = i[92];
  assign o[47264] = i[92];
  assign o[47265] = i[92];
  assign o[47266] = i[92];
  assign o[47267] = i[92];
  assign o[47268] = i[92];
  assign o[47269] = i[92];
  assign o[47270] = i[92];
  assign o[47271] = i[92];
  assign o[47272] = i[92];
  assign o[47273] = i[92];
  assign o[47274] = i[92];
  assign o[47275] = i[92];
  assign o[47276] = i[92];
  assign o[47277] = i[92];
  assign o[47278] = i[92];
  assign o[47279] = i[92];
  assign o[47280] = i[92];
  assign o[47281] = i[92];
  assign o[47282] = i[92];
  assign o[47283] = i[92];
  assign o[47284] = i[92];
  assign o[47285] = i[92];
  assign o[47286] = i[92];
  assign o[47287] = i[92];
  assign o[47288] = i[92];
  assign o[47289] = i[92];
  assign o[47290] = i[92];
  assign o[47291] = i[92];
  assign o[47292] = i[92];
  assign o[47293] = i[92];
  assign o[47294] = i[92];
  assign o[47295] = i[92];
  assign o[47296] = i[92];
  assign o[47297] = i[92];
  assign o[47298] = i[92];
  assign o[47299] = i[92];
  assign o[47300] = i[92];
  assign o[47301] = i[92];
  assign o[47302] = i[92];
  assign o[47303] = i[92];
  assign o[47304] = i[92];
  assign o[47305] = i[92];
  assign o[47306] = i[92];
  assign o[47307] = i[92];
  assign o[47308] = i[92];
  assign o[47309] = i[92];
  assign o[47310] = i[92];
  assign o[47311] = i[92];
  assign o[47312] = i[92];
  assign o[47313] = i[92];
  assign o[47314] = i[92];
  assign o[47315] = i[92];
  assign o[47316] = i[92];
  assign o[47317] = i[92];
  assign o[47318] = i[92];
  assign o[47319] = i[92];
  assign o[47320] = i[92];
  assign o[47321] = i[92];
  assign o[47322] = i[92];
  assign o[47323] = i[92];
  assign o[47324] = i[92];
  assign o[47325] = i[92];
  assign o[47326] = i[92];
  assign o[47327] = i[92];
  assign o[47328] = i[92];
  assign o[47329] = i[92];
  assign o[47330] = i[92];
  assign o[47331] = i[92];
  assign o[47332] = i[92];
  assign o[47333] = i[92];
  assign o[47334] = i[92];
  assign o[47335] = i[92];
  assign o[47336] = i[92];
  assign o[47337] = i[92];
  assign o[47338] = i[92];
  assign o[47339] = i[92];
  assign o[47340] = i[92];
  assign o[47341] = i[92];
  assign o[47342] = i[92];
  assign o[47343] = i[92];
  assign o[47344] = i[92];
  assign o[47345] = i[92];
  assign o[47346] = i[92];
  assign o[47347] = i[92];
  assign o[47348] = i[92];
  assign o[47349] = i[92];
  assign o[47350] = i[92];
  assign o[47351] = i[92];
  assign o[47352] = i[92];
  assign o[47353] = i[92];
  assign o[47354] = i[92];
  assign o[47355] = i[92];
  assign o[47356] = i[92];
  assign o[47357] = i[92];
  assign o[47358] = i[92];
  assign o[47359] = i[92];
  assign o[47360] = i[92];
  assign o[47361] = i[92];
  assign o[47362] = i[92];
  assign o[47363] = i[92];
  assign o[47364] = i[92];
  assign o[47365] = i[92];
  assign o[47366] = i[92];
  assign o[47367] = i[92];
  assign o[47368] = i[92];
  assign o[47369] = i[92];
  assign o[47370] = i[92];
  assign o[47371] = i[92];
  assign o[47372] = i[92];
  assign o[47373] = i[92];
  assign o[47374] = i[92];
  assign o[47375] = i[92];
  assign o[47376] = i[92];
  assign o[47377] = i[92];
  assign o[47378] = i[92];
  assign o[47379] = i[92];
  assign o[47380] = i[92];
  assign o[47381] = i[92];
  assign o[47382] = i[92];
  assign o[47383] = i[92];
  assign o[47384] = i[92];
  assign o[47385] = i[92];
  assign o[47386] = i[92];
  assign o[47387] = i[92];
  assign o[47388] = i[92];
  assign o[47389] = i[92];
  assign o[47390] = i[92];
  assign o[47391] = i[92];
  assign o[47392] = i[92];
  assign o[47393] = i[92];
  assign o[47394] = i[92];
  assign o[47395] = i[92];
  assign o[47396] = i[92];
  assign o[47397] = i[92];
  assign o[47398] = i[92];
  assign o[47399] = i[92];
  assign o[47400] = i[92];
  assign o[47401] = i[92];
  assign o[47402] = i[92];
  assign o[47403] = i[92];
  assign o[47404] = i[92];
  assign o[47405] = i[92];
  assign o[47406] = i[92];
  assign o[47407] = i[92];
  assign o[47408] = i[92];
  assign o[47409] = i[92];
  assign o[47410] = i[92];
  assign o[47411] = i[92];
  assign o[47412] = i[92];
  assign o[47413] = i[92];
  assign o[47414] = i[92];
  assign o[47415] = i[92];
  assign o[47416] = i[92];
  assign o[47417] = i[92];
  assign o[47418] = i[92];
  assign o[47419] = i[92];
  assign o[47420] = i[92];
  assign o[47421] = i[92];
  assign o[47422] = i[92];
  assign o[47423] = i[92];
  assign o[47424] = i[92];
  assign o[47425] = i[92];
  assign o[47426] = i[92];
  assign o[47427] = i[92];
  assign o[47428] = i[92];
  assign o[47429] = i[92];
  assign o[47430] = i[92];
  assign o[47431] = i[92];
  assign o[47432] = i[92];
  assign o[47433] = i[92];
  assign o[47434] = i[92];
  assign o[47435] = i[92];
  assign o[47436] = i[92];
  assign o[47437] = i[92];
  assign o[47438] = i[92];
  assign o[47439] = i[92];
  assign o[47440] = i[92];
  assign o[47441] = i[92];
  assign o[47442] = i[92];
  assign o[47443] = i[92];
  assign o[47444] = i[92];
  assign o[47445] = i[92];
  assign o[47446] = i[92];
  assign o[47447] = i[92];
  assign o[47448] = i[92];
  assign o[47449] = i[92];
  assign o[47450] = i[92];
  assign o[47451] = i[92];
  assign o[47452] = i[92];
  assign o[47453] = i[92];
  assign o[47454] = i[92];
  assign o[47455] = i[92];
  assign o[47456] = i[92];
  assign o[47457] = i[92];
  assign o[47458] = i[92];
  assign o[47459] = i[92];
  assign o[47460] = i[92];
  assign o[47461] = i[92];
  assign o[47462] = i[92];
  assign o[47463] = i[92];
  assign o[47464] = i[92];
  assign o[47465] = i[92];
  assign o[47466] = i[92];
  assign o[47467] = i[92];
  assign o[47468] = i[92];
  assign o[47469] = i[92];
  assign o[47470] = i[92];
  assign o[47471] = i[92];
  assign o[47472] = i[92];
  assign o[47473] = i[92];
  assign o[47474] = i[92];
  assign o[47475] = i[92];
  assign o[47476] = i[92];
  assign o[47477] = i[92];
  assign o[47478] = i[92];
  assign o[47479] = i[92];
  assign o[47480] = i[92];
  assign o[47481] = i[92];
  assign o[47482] = i[92];
  assign o[47483] = i[92];
  assign o[47484] = i[92];
  assign o[47485] = i[92];
  assign o[47486] = i[92];
  assign o[47487] = i[92];
  assign o[47488] = i[92];
  assign o[47489] = i[92];
  assign o[47490] = i[92];
  assign o[47491] = i[92];
  assign o[47492] = i[92];
  assign o[47493] = i[92];
  assign o[47494] = i[92];
  assign o[47495] = i[92];
  assign o[47496] = i[92];
  assign o[47497] = i[92];
  assign o[47498] = i[92];
  assign o[47499] = i[92];
  assign o[47500] = i[92];
  assign o[47501] = i[92];
  assign o[47502] = i[92];
  assign o[47503] = i[92];
  assign o[47504] = i[92];
  assign o[47505] = i[92];
  assign o[47506] = i[92];
  assign o[47507] = i[92];
  assign o[47508] = i[92];
  assign o[47509] = i[92];
  assign o[47510] = i[92];
  assign o[47511] = i[92];
  assign o[47512] = i[92];
  assign o[47513] = i[92];
  assign o[47514] = i[92];
  assign o[47515] = i[92];
  assign o[47516] = i[92];
  assign o[47517] = i[92];
  assign o[47518] = i[92];
  assign o[47519] = i[92];
  assign o[47520] = i[92];
  assign o[47521] = i[92];
  assign o[47522] = i[92];
  assign o[47523] = i[92];
  assign o[47524] = i[92];
  assign o[47525] = i[92];
  assign o[47526] = i[92];
  assign o[47527] = i[92];
  assign o[47528] = i[92];
  assign o[47529] = i[92];
  assign o[47530] = i[92];
  assign o[47531] = i[92];
  assign o[47532] = i[92];
  assign o[47533] = i[92];
  assign o[47534] = i[92];
  assign o[47535] = i[92];
  assign o[47536] = i[92];
  assign o[47537] = i[92];
  assign o[47538] = i[92];
  assign o[47539] = i[92];
  assign o[47540] = i[92];
  assign o[47541] = i[92];
  assign o[47542] = i[92];
  assign o[47543] = i[92];
  assign o[47544] = i[92];
  assign o[47545] = i[92];
  assign o[47546] = i[92];
  assign o[47547] = i[92];
  assign o[47548] = i[92];
  assign o[47549] = i[92];
  assign o[47550] = i[92];
  assign o[47551] = i[92];
  assign o[47552] = i[92];
  assign o[47553] = i[92];
  assign o[47554] = i[92];
  assign o[47555] = i[92];
  assign o[47556] = i[92];
  assign o[47557] = i[92];
  assign o[47558] = i[92];
  assign o[47559] = i[92];
  assign o[47560] = i[92];
  assign o[47561] = i[92];
  assign o[47562] = i[92];
  assign o[47563] = i[92];
  assign o[47564] = i[92];
  assign o[47565] = i[92];
  assign o[47566] = i[92];
  assign o[47567] = i[92];
  assign o[47568] = i[92];
  assign o[47569] = i[92];
  assign o[47570] = i[92];
  assign o[47571] = i[92];
  assign o[47572] = i[92];
  assign o[47573] = i[92];
  assign o[47574] = i[92];
  assign o[47575] = i[92];
  assign o[47576] = i[92];
  assign o[47577] = i[92];
  assign o[47578] = i[92];
  assign o[47579] = i[92];
  assign o[47580] = i[92];
  assign o[47581] = i[92];
  assign o[47582] = i[92];
  assign o[47583] = i[92];
  assign o[47584] = i[92];
  assign o[47585] = i[92];
  assign o[47586] = i[92];
  assign o[47587] = i[92];
  assign o[47588] = i[92];
  assign o[47589] = i[92];
  assign o[47590] = i[92];
  assign o[47591] = i[92];
  assign o[47592] = i[92];
  assign o[47593] = i[92];
  assign o[47594] = i[92];
  assign o[47595] = i[92];
  assign o[47596] = i[92];
  assign o[47597] = i[92];
  assign o[47598] = i[92];
  assign o[47599] = i[92];
  assign o[47600] = i[92];
  assign o[47601] = i[92];
  assign o[47602] = i[92];
  assign o[47603] = i[92];
  assign o[47604] = i[92];
  assign o[47605] = i[92];
  assign o[47606] = i[92];
  assign o[47607] = i[92];
  assign o[47608] = i[92];
  assign o[47609] = i[92];
  assign o[47610] = i[92];
  assign o[47611] = i[92];
  assign o[47612] = i[92];
  assign o[47613] = i[92];
  assign o[47614] = i[92];
  assign o[47615] = i[92];
  assign o[46592] = i[91];
  assign o[46593] = i[91];
  assign o[46594] = i[91];
  assign o[46595] = i[91];
  assign o[46596] = i[91];
  assign o[46597] = i[91];
  assign o[46598] = i[91];
  assign o[46599] = i[91];
  assign o[46600] = i[91];
  assign o[46601] = i[91];
  assign o[46602] = i[91];
  assign o[46603] = i[91];
  assign o[46604] = i[91];
  assign o[46605] = i[91];
  assign o[46606] = i[91];
  assign o[46607] = i[91];
  assign o[46608] = i[91];
  assign o[46609] = i[91];
  assign o[46610] = i[91];
  assign o[46611] = i[91];
  assign o[46612] = i[91];
  assign o[46613] = i[91];
  assign o[46614] = i[91];
  assign o[46615] = i[91];
  assign o[46616] = i[91];
  assign o[46617] = i[91];
  assign o[46618] = i[91];
  assign o[46619] = i[91];
  assign o[46620] = i[91];
  assign o[46621] = i[91];
  assign o[46622] = i[91];
  assign o[46623] = i[91];
  assign o[46624] = i[91];
  assign o[46625] = i[91];
  assign o[46626] = i[91];
  assign o[46627] = i[91];
  assign o[46628] = i[91];
  assign o[46629] = i[91];
  assign o[46630] = i[91];
  assign o[46631] = i[91];
  assign o[46632] = i[91];
  assign o[46633] = i[91];
  assign o[46634] = i[91];
  assign o[46635] = i[91];
  assign o[46636] = i[91];
  assign o[46637] = i[91];
  assign o[46638] = i[91];
  assign o[46639] = i[91];
  assign o[46640] = i[91];
  assign o[46641] = i[91];
  assign o[46642] = i[91];
  assign o[46643] = i[91];
  assign o[46644] = i[91];
  assign o[46645] = i[91];
  assign o[46646] = i[91];
  assign o[46647] = i[91];
  assign o[46648] = i[91];
  assign o[46649] = i[91];
  assign o[46650] = i[91];
  assign o[46651] = i[91];
  assign o[46652] = i[91];
  assign o[46653] = i[91];
  assign o[46654] = i[91];
  assign o[46655] = i[91];
  assign o[46656] = i[91];
  assign o[46657] = i[91];
  assign o[46658] = i[91];
  assign o[46659] = i[91];
  assign o[46660] = i[91];
  assign o[46661] = i[91];
  assign o[46662] = i[91];
  assign o[46663] = i[91];
  assign o[46664] = i[91];
  assign o[46665] = i[91];
  assign o[46666] = i[91];
  assign o[46667] = i[91];
  assign o[46668] = i[91];
  assign o[46669] = i[91];
  assign o[46670] = i[91];
  assign o[46671] = i[91];
  assign o[46672] = i[91];
  assign o[46673] = i[91];
  assign o[46674] = i[91];
  assign o[46675] = i[91];
  assign o[46676] = i[91];
  assign o[46677] = i[91];
  assign o[46678] = i[91];
  assign o[46679] = i[91];
  assign o[46680] = i[91];
  assign o[46681] = i[91];
  assign o[46682] = i[91];
  assign o[46683] = i[91];
  assign o[46684] = i[91];
  assign o[46685] = i[91];
  assign o[46686] = i[91];
  assign o[46687] = i[91];
  assign o[46688] = i[91];
  assign o[46689] = i[91];
  assign o[46690] = i[91];
  assign o[46691] = i[91];
  assign o[46692] = i[91];
  assign o[46693] = i[91];
  assign o[46694] = i[91];
  assign o[46695] = i[91];
  assign o[46696] = i[91];
  assign o[46697] = i[91];
  assign o[46698] = i[91];
  assign o[46699] = i[91];
  assign o[46700] = i[91];
  assign o[46701] = i[91];
  assign o[46702] = i[91];
  assign o[46703] = i[91];
  assign o[46704] = i[91];
  assign o[46705] = i[91];
  assign o[46706] = i[91];
  assign o[46707] = i[91];
  assign o[46708] = i[91];
  assign o[46709] = i[91];
  assign o[46710] = i[91];
  assign o[46711] = i[91];
  assign o[46712] = i[91];
  assign o[46713] = i[91];
  assign o[46714] = i[91];
  assign o[46715] = i[91];
  assign o[46716] = i[91];
  assign o[46717] = i[91];
  assign o[46718] = i[91];
  assign o[46719] = i[91];
  assign o[46720] = i[91];
  assign o[46721] = i[91];
  assign o[46722] = i[91];
  assign o[46723] = i[91];
  assign o[46724] = i[91];
  assign o[46725] = i[91];
  assign o[46726] = i[91];
  assign o[46727] = i[91];
  assign o[46728] = i[91];
  assign o[46729] = i[91];
  assign o[46730] = i[91];
  assign o[46731] = i[91];
  assign o[46732] = i[91];
  assign o[46733] = i[91];
  assign o[46734] = i[91];
  assign o[46735] = i[91];
  assign o[46736] = i[91];
  assign o[46737] = i[91];
  assign o[46738] = i[91];
  assign o[46739] = i[91];
  assign o[46740] = i[91];
  assign o[46741] = i[91];
  assign o[46742] = i[91];
  assign o[46743] = i[91];
  assign o[46744] = i[91];
  assign o[46745] = i[91];
  assign o[46746] = i[91];
  assign o[46747] = i[91];
  assign o[46748] = i[91];
  assign o[46749] = i[91];
  assign o[46750] = i[91];
  assign o[46751] = i[91];
  assign o[46752] = i[91];
  assign o[46753] = i[91];
  assign o[46754] = i[91];
  assign o[46755] = i[91];
  assign o[46756] = i[91];
  assign o[46757] = i[91];
  assign o[46758] = i[91];
  assign o[46759] = i[91];
  assign o[46760] = i[91];
  assign o[46761] = i[91];
  assign o[46762] = i[91];
  assign o[46763] = i[91];
  assign o[46764] = i[91];
  assign o[46765] = i[91];
  assign o[46766] = i[91];
  assign o[46767] = i[91];
  assign o[46768] = i[91];
  assign o[46769] = i[91];
  assign o[46770] = i[91];
  assign o[46771] = i[91];
  assign o[46772] = i[91];
  assign o[46773] = i[91];
  assign o[46774] = i[91];
  assign o[46775] = i[91];
  assign o[46776] = i[91];
  assign o[46777] = i[91];
  assign o[46778] = i[91];
  assign o[46779] = i[91];
  assign o[46780] = i[91];
  assign o[46781] = i[91];
  assign o[46782] = i[91];
  assign o[46783] = i[91];
  assign o[46784] = i[91];
  assign o[46785] = i[91];
  assign o[46786] = i[91];
  assign o[46787] = i[91];
  assign o[46788] = i[91];
  assign o[46789] = i[91];
  assign o[46790] = i[91];
  assign o[46791] = i[91];
  assign o[46792] = i[91];
  assign o[46793] = i[91];
  assign o[46794] = i[91];
  assign o[46795] = i[91];
  assign o[46796] = i[91];
  assign o[46797] = i[91];
  assign o[46798] = i[91];
  assign o[46799] = i[91];
  assign o[46800] = i[91];
  assign o[46801] = i[91];
  assign o[46802] = i[91];
  assign o[46803] = i[91];
  assign o[46804] = i[91];
  assign o[46805] = i[91];
  assign o[46806] = i[91];
  assign o[46807] = i[91];
  assign o[46808] = i[91];
  assign o[46809] = i[91];
  assign o[46810] = i[91];
  assign o[46811] = i[91];
  assign o[46812] = i[91];
  assign o[46813] = i[91];
  assign o[46814] = i[91];
  assign o[46815] = i[91];
  assign o[46816] = i[91];
  assign o[46817] = i[91];
  assign o[46818] = i[91];
  assign o[46819] = i[91];
  assign o[46820] = i[91];
  assign o[46821] = i[91];
  assign o[46822] = i[91];
  assign o[46823] = i[91];
  assign o[46824] = i[91];
  assign o[46825] = i[91];
  assign o[46826] = i[91];
  assign o[46827] = i[91];
  assign o[46828] = i[91];
  assign o[46829] = i[91];
  assign o[46830] = i[91];
  assign o[46831] = i[91];
  assign o[46832] = i[91];
  assign o[46833] = i[91];
  assign o[46834] = i[91];
  assign o[46835] = i[91];
  assign o[46836] = i[91];
  assign o[46837] = i[91];
  assign o[46838] = i[91];
  assign o[46839] = i[91];
  assign o[46840] = i[91];
  assign o[46841] = i[91];
  assign o[46842] = i[91];
  assign o[46843] = i[91];
  assign o[46844] = i[91];
  assign o[46845] = i[91];
  assign o[46846] = i[91];
  assign o[46847] = i[91];
  assign o[46848] = i[91];
  assign o[46849] = i[91];
  assign o[46850] = i[91];
  assign o[46851] = i[91];
  assign o[46852] = i[91];
  assign o[46853] = i[91];
  assign o[46854] = i[91];
  assign o[46855] = i[91];
  assign o[46856] = i[91];
  assign o[46857] = i[91];
  assign o[46858] = i[91];
  assign o[46859] = i[91];
  assign o[46860] = i[91];
  assign o[46861] = i[91];
  assign o[46862] = i[91];
  assign o[46863] = i[91];
  assign o[46864] = i[91];
  assign o[46865] = i[91];
  assign o[46866] = i[91];
  assign o[46867] = i[91];
  assign o[46868] = i[91];
  assign o[46869] = i[91];
  assign o[46870] = i[91];
  assign o[46871] = i[91];
  assign o[46872] = i[91];
  assign o[46873] = i[91];
  assign o[46874] = i[91];
  assign o[46875] = i[91];
  assign o[46876] = i[91];
  assign o[46877] = i[91];
  assign o[46878] = i[91];
  assign o[46879] = i[91];
  assign o[46880] = i[91];
  assign o[46881] = i[91];
  assign o[46882] = i[91];
  assign o[46883] = i[91];
  assign o[46884] = i[91];
  assign o[46885] = i[91];
  assign o[46886] = i[91];
  assign o[46887] = i[91];
  assign o[46888] = i[91];
  assign o[46889] = i[91];
  assign o[46890] = i[91];
  assign o[46891] = i[91];
  assign o[46892] = i[91];
  assign o[46893] = i[91];
  assign o[46894] = i[91];
  assign o[46895] = i[91];
  assign o[46896] = i[91];
  assign o[46897] = i[91];
  assign o[46898] = i[91];
  assign o[46899] = i[91];
  assign o[46900] = i[91];
  assign o[46901] = i[91];
  assign o[46902] = i[91];
  assign o[46903] = i[91];
  assign o[46904] = i[91];
  assign o[46905] = i[91];
  assign o[46906] = i[91];
  assign o[46907] = i[91];
  assign o[46908] = i[91];
  assign o[46909] = i[91];
  assign o[46910] = i[91];
  assign o[46911] = i[91];
  assign o[46912] = i[91];
  assign o[46913] = i[91];
  assign o[46914] = i[91];
  assign o[46915] = i[91];
  assign o[46916] = i[91];
  assign o[46917] = i[91];
  assign o[46918] = i[91];
  assign o[46919] = i[91];
  assign o[46920] = i[91];
  assign o[46921] = i[91];
  assign o[46922] = i[91];
  assign o[46923] = i[91];
  assign o[46924] = i[91];
  assign o[46925] = i[91];
  assign o[46926] = i[91];
  assign o[46927] = i[91];
  assign o[46928] = i[91];
  assign o[46929] = i[91];
  assign o[46930] = i[91];
  assign o[46931] = i[91];
  assign o[46932] = i[91];
  assign o[46933] = i[91];
  assign o[46934] = i[91];
  assign o[46935] = i[91];
  assign o[46936] = i[91];
  assign o[46937] = i[91];
  assign o[46938] = i[91];
  assign o[46939] = i[91];
  assign o[46940] = i[91];
  assign o[46941] = i[91];
  assign o[46942] = i[91];
  assign o[46943] = i[91];
  assign o[46944] = i[91];
  assign o[46945] = i[91];
  assign o[46946] = i[91];
  assign o[46947] = i[91];
  assign o[46948] = i[91];
  assign o[46949] = i[91];
  assign o[46950] = i[91];
  assign o[46951] = i[91];
  assign o[46952] = i[91];
  assign o[46953] = i[91];
  assign o[46954] = i[91];
  assign o[46955] = i[91];
  assign o[46956] = i[91];
  assign o[46957] = i[91];
  assign o[46958] = i[91];
  assign o[46959] = i[91];
  assign o[46960] = i[91];
  assign o[46961] = i[91];
  assign o[46962] = i[91];
  assign o[46963] = i[91];
  assign o[46964] = i[91];
  assign o[46965] = i[91];
  assign o[46966] = i[91];
  assign o[46967] = i[91];
  assign o[46968] = i[91];
  assign o[46969] = i[91];
  assign o[46970] = i[91];
  assign o[46971] = i[91];
  assign o[46972] = i[91];
  assign o[46973] = i[91];
  assign o[46974] = i[91];
  assign o[46975] = i[91];
  assign o[46976] = i[91];
  assign o[46977] = i[91];
  assign o[46978] = i[91];
  assign o[46979] = i[91];
  assign o[46980] = i[91];
  assign o[46981] = i[91];
  assign o[46982] = i[91];
  assign o[46983] = i[91];
  assign o[46984] = i[91];
  assign o[46985] = i[91];
  assign o[46986] = i[91];
  assign o[46987] = i[91];
  assign o[46988] = i[91];
  assign o[46989] = i[91];
  assign o[46990] = i[91];
  assign o[46991] = i[91];
  assign o[46992] = i[91];
  assign o[46993] = i[91];
  assign o[46994] = i[91];
  assign o[46995] = i[91];
  assign o[46996] = i[91];
  assign o[46997] = i[91];
  assign o[46998] = i[91];
  assign o[46999] = i[91];
  assign o[47000] = i[91];
  assign o[47001] = i[91];
  assign o[47002] = i[91];
  assign o[47003] = i[91];
  assign o[47004] = i[91];
  assign o[47005] = i[91];
  assign o[47006] = i[91];
  assign o[47007] = i[91];
  assign o[47008] = i[91];
  assign o[47009] = i[91];
  assign o[47010] = i[91];
  assign o[47011] = i[91];
  assign o[47012] = i[91];
  assign o[47013] = i[91];
  assign o[47014] = i[91];
  assign o[47015] = i[91];
  assign o[47016] = i[91];
  assign o[47017] = i[91];
  assign o[47018] = i[91];
  assign o[47019] = i[91];
  assign o[47020] = i[91];
  assign o[47021] = i[91];
  assign o[47022] = i[91];
  assign o[47023] = i[91];
  assign o[47024] = i[91];
  assign o[47025] = i[91];
  assign o[47026] = i[91];
  assign o[47027] = i[91];
  assign o[47028] = i[91];
  assign o[47029] = i[91];
  assign o[47030] = i[91];
  assign o[47031] = i[91];
  assign o[47032] = i[91];
  assign o[47033] = i[91];
  assign o[47034] = i[91];
  assign o[47035] = i[91];
  assign o[47036] = i[91];
  assign o[47037] = i[91];
  assign o[47038] = i[91];
  assign o[47039] = i[91];
  assign o[47040] = i[91];
  assign o[47041] = i[91];
  assign o[47042] = i[91];
  assign o[47043] = i[91];
  assign o[47044] = i[91];
  assign o[47045] = i[91];
  assign o[47046] = i[91];
  assign o[47047] = i[91];
  assign o[47048] = i[91];
  assign o[47049] = i[91];
  assign o[47050] = i[91];
  assign o[47051] = i[91];
  assign o[47052] = i[91];
  assign o[47053] = i[91];
  assign o[47054] = i[91];
  assign o[47055] = i[91];
  assign o[47056] = i[91];
  assign o[47057] = i[91];
  assign o[47058] = i[91];
  assign o[47059] = i[91];
  assign o[47060] = i[91];
  assign o[47061] = i[91];
  assign o[47062] = i[91];
  assign o[47063] = i[91];
  assign o[47064] = i[91];
  assign o[47065] = i[91];
  assign o[47066] = i[91];
  assign o[47067] = i[91];
  assign o[47068] = i[91];
  assign o[47069] = i[91];
  assign o[47070] = i[91];
  assign o[47071] = i[91];
  assign o[47072] = i[91];
  assign o[47073] = i[91];
  assign o[47074] = i[91];
  assign o[47075] = i[91];
  assign o[47076] = i[91];
  assign o[47077] = i[91];
  assign o[47078] = i[91];
  assign o[47079] = i[91];
  assign o[47080] = i[91];
  assign o[47081] = i[91];
  assign o[47082] = i[91];
  assign o[47083] = i[91];
  assign o[47084] = i[91];
  assign o[47085] = i[91];
  assign o[47086] = i[91];
  assign o[47087] = i[91];
  assign o[47088] = i[91];
  assign o[47089] = i[91];
  assign o[47090] = i[91];
  assign o[47091] = i[91];
  assign o[47092] = i[91];
  assign o[47093] = i[91];
  assign o[47094] = i[91];
  assign o[47095] = i[91];
  assign o[47096] = i[91];
  assign o[47097] = i[91];
  assign o[47098] = i[91];
  assign o[47099] = i[91];
  assign o[47100] = i[91];
  assign o[47101] = i[91];
  assign o[47102] = i[91];
  assign o[47103] = i[91];
  assign o[46080] = i[90];
  assign o[46081] = i[90];
  assign o[46082] = i[90];
  assign o[46083] = i[90];
  assign o[46084] = i[90];
  assign o[46085] = i[90];
  assign o[46086] = i[90];
  assign o[46087] = i[90];
  assign o[46088] = i[90];
  assign o[46089] = i[90];
  assign o[46090] = i[90];
  assign o[46091] = i[90];
  assign o[46092] = i[90];
  assign o[46093] = i[90];
  assign o[46094] = i[90];
  assign o[46095] = i[90];
  assign o[46096] = i[90];
  assign o[46097] = i[90];
  assign o[46098] = i[90];
  assign o[46099] = i[90];
  assign o[46100] = i[90];
  assign o[46101] = i[90];
  assign o[46102] = i[90];
  assign o[46103] = i[90];
  assign o[46104] = i[90];
  assign o[46105] = i[90];
  assign o[46106] = i[90];
  assign o[46107] = i[90];
  assign o[46108] = i[90];
  assign o[46109] = i[90];
  assign o[46110] = i[90];
  assign o[46111] = i[90];
  assign o[46112] = i[90];
  assign o[46113] = i[90];
  assign o[46114] = i[90];
  assign o[46115] = i[90];
  assign o[46116] = i[90];
  assign o[46117] = i[90];
  assign o[46118] = i[90];
  assign o[46119] = i[90];
  assign o[46120] = i[90];
  assign o[46121] = i[90];
  assign o[46122] = i[90];
  assign o[46123] = i[90];
  assign o[46124] = i[90];
  assign o[46125] = i[90];
  assign o[46126] = i[90];
  assign o[46127] = i[90];
  assign o[46128] = i[90];
  assign o[46129] = i[90];
  assign o[46130] = i[90];
  assign o[46131] = i[90];
  assign o[46132] = i[90];
  assign o[46133] = i[90];
  assign o[46134] = i[90];
  assign o[46135] = i[90];
  assign o[46136] = i[90];
  assign o[46137] = i[90];
  assign o[46138] = i[90];
  assign o[46139] = i[90];
  assign o[46140] = i[90];
  assign o[46141] = i[90];
  assign o[46142] = i[90];
  assign o[46143] = i[90];
  assign o[46144] = i[90];
  assign o[46145] = i[90];
  assign o[46146] = i[90];
  assign o[46147] = i[90];
  assign o[46148] = i[90];
  assign o[46149] = i[90];
  assign o[46150] = i[90];
  assign o[46151] = i[90];
  assign o[46152] = i[90];
  assign o[46153] = i[90];
  assign o[46154] = i[90];
  assign o[46155] = i[90];
  assign o[46156] = i[90];
  assign o[46157] = i[90];
  assign o[46158] = i[90];
  assign o[46159] = i[90];
  assign o[46160] = i[90];
  assign o[46161] = i[90];
  assign o[46162] = i[90];
  assign o[46163] = i[90];
  assign o[46164] = i[90];
  assign o[46165] = i[90];
  assign o[46166] = i[90];
  assign o[46167] = i[90];
  assign o[46168] = i[90];
  assign o[46169] = i[90];
  assign o[46170] = i[90];
  assign o[46171] = i[90];
  assign o[46172] = i[90];
  assign o[46173] = i[90];
  assign o[46174] = i[90];
  assign o[46175] = i[90];
  assign o[46176] = i[90];
  assign o[46177] = i[90];
  assign o[46178] = i[90];
  assign o[46179] = i[90];
  assign o[46180] = i[90];
  assign o[46181] = i[90];
  assign o[46182] = i[90];
  assign o[46183] = i[90];
  assign o[46184] = i[90];
  assign o[46185] = i[90];
  assign o[46186] = i[90];
  assign o[46187] = i[90];
  assign o[46188] = i[90];
  assign o[46189] = i[90];
  assign o[46190] = i[90];
  assign o[46191] = i[90];
  assign o[46192] = i[90];
  assign o[46193] = i[90];
  assign o[46194] = i[90];
  assign o[46195] = i[90];
  assign o[46196] = i[90];
  assign o[46197] = i[90];
  assign o[46198] = i[90];
  assign o[46199] = i[90];
  assign o[46200] = i[90];
  assign o[46201] = i[90];
  assign o[46202] = i[90];
  assign o[46203] = i[90];
  assign o[46204] = i[90];
  assign o[46205] = i[90];
  assign o[46206] = i[90];
  assign o[46207] = i[90];
  assign o[46208] = i[90];
  assign o[46209] = i[90];
  assign o[46210] = i[90];
  assign o[46211] = i[90];
  assign o[46212] = i[90];
  assign o[46213] = i[90];
  assign o[46214] = i[90];
  assign o[46215] = i[90];
  assign o[46216] = i[90];
  assign o[46217] = i[90];
  assign o[46218] = i[90];
  assign o[46219] = i[90];
  assign o[46220] = i[90];
  assign o[46221] = i[90];
  assign o[46222] = i[90];
  assign o[46223] = i[90];
  assign o[46224] = i[90];
  assign o[46225] = i[90];
  assign o[46226] = i[90];
  assign o[46227] = i[90];
  assign o[46228] = i[90];
  assign o[46229] = i[90];
  assign o[46230] = i[90];
  assign o[46231] = i[90];
  assign o[46232] = i[90];
  assign o[46233] = i[90];
  assign o[46234] = i[90];
  assign o[46235] = i[90];
  assign o[46236] = i[90];
  assign o[46237] = i[90];
  assign o[46238] = i[90];
  assign o[46239] = i[90];
  assign o[46240] = i[90];
  assign o[46241] = i[90];
  assign o[46242] = i[90];
  assign o[46243] = i[90];
  assign o[46244] = i[90];
  assign o[46245] = i[90];
  assign o[46246] = i[90];
  assign o[46247] = i[90];
  assign o[46248] = i[90];
  assign o[46249] = i[90];
  assign o[46250] = i[90];
  assign o[46251] = i[90];
  assign o[46252] = i[90];
  assign o[46253] = i[90];
  assign o[46254] = i[90];
  assign o[46255] = i[90];
  assign o[46256] = i[90];
  assign o[46257] = i[90];
  assign o[46258] = i[90];
  assign o[46259] = i[90];
  assign o[46260] = i[90];
  assign o[46261] = i[90];
  assign o[46262] = i[90];
  assign o[46263] = i[90];
  assign o[46264] = i[90];
  assign o[46265] = i[90];
  assign o[46266] = i[90];
  assign o[46267] = i[90];
  assign o[46268] = i[90];
  assign o[46269] = i[90];
  assign o[46270] = i[90];
  assign o[46271] = i[90];
  assign o[46272] = i[90];
  assign o[46273] = i[90];
  assign o[46274] = i[90];
  assign o[46275] = i[90];
  assign o[46276] = i[90];
  assign o[46277] = i[90];
  assign o[46278] = i[90];
  assign o[46279] = i[90];
  assign o[46280] = i[90];
  assign o[46281] = i[90];
  assign o[46282] = i[90];
  assign o[46283] = i[90];
  assign o[46284] = i[90];
  assign o[46285] = i[90];
  assign o[46286] = i[90];
  assign o[46287] = i[90];
  assign o[46288] = i[90];
  assign o[46289] = i[90];
  assign o[46290] = i[90];
  assign o[46291] = i[90];
  assign o[46292] = i[90];
  assign o[46293] = i[90];
  assign o[46294] = i[90];
  assign o[46295] = i[90];
  assign o[46296] = i[90];
  assign o[46297] = i[90];
  assign o[46298] = i[90];
  assign o[46299] = i[90];
  assign o[46300] = i[90];
  assign o[46301] = i[90];
  assign o[46302] = i[90];
  assign o[46303] = i[90];
  assign o[46304] = i[90];
  assign o[46305] = i[90];
  assign o[46306] = i[90];
  assign o[46307] = i[90];
  assign o[46308] = i[90];
  assign o[46309] = i[90];
  assign o[46310] = i[90];
  assign o[46311] = i[90];
  assign o[46312] = i[90];
  assign o[46313] = i[90];
  assign o[46314] = i[90];
  assign o[46315] = i[90];
  assign o[46316] = i[90];
  assign o[46317] = i[90];
  assign o[46318] = i[90];
  assign o[46319] = i[90];
  assign o[46320] = i[90];
  assign o[46321] = i[90];
  assign o[46322] = i[90];
  assign o[46323] = i[90];
  assign o[46324] = i[90];
  assign o[46325] = i[90];
  assign o[46326] = i[90];
  assign o[46327] = i[90];
  assign o[46328] = i[90];
  assign o[46329] = i[90];
  assign o[46330] = i[90];
  assign o[46331] = i[90];
  assign o[46332] = i[90];
  assign o[46333] = i[90];
  assign o[46334] = i[90];
  assign o[46335] = i[90];
  assign o[46336] = i[90];
  assign o[46337] = i[90];
  assign o[46338] = i[90];
  assign o[46339] = i[90];
  assign o[46340] = i[90];
  assign o[46341] = i[90];
  assign o[46342] = i[90];
  assign o[46343] = i[90];
  assign o[46344] = i[90];
  assign o[46345] = i[90];
  assign o[46346] = i[90];
  assign o[46347] = i[90];
  assign o[46348] = i[90];
  assign o[46349] = i[90];
  assign o[46350] = i[90];
  assign o[46351] = i[90];
  assign o[46352] = i[90];
  assign o[46353] = i[90];
  assign o[46354] = i[90];
  assign o[46355] = i[90];
  assign o[46356] = i[90];
  assign o[46357] = i[90];
  assign o[46358] = i[90];
  assign o[46359] = i[90];
  assign o[46360] = i[90];
  assign o[46361] = i[90];
  assign o[46362] = i[90];
  assign o[46363] = i[90];
  assign o[46364] = i[90];
  assign o[46365] = i[90];
  assign o[46366] = i[90];
  assign o[46367] = i[90];
  assign o[46368] = i[90];
  assign o[46369] = i[90];
  assign o[46370] = i[90];
  assign o[46371] = i[90];
  assign o[46372] = i[90];
  assign o[46373] = i[90];
  assign o[46374] = i[90];
  assign o[46375] = i[90];
  assign o[46376] = i[90];
  assign o[46377] = i[90];
  assign o[46378] = i[90];
  assign o[46379] = i[90];
  assign o[46380] = i[90];
  assign o[46381] = i[90];
  assign o[46382] = i[90];
  assign o[46383] = i[90];
  assign o[46384] = i[90];
  assign o[46385] = i[90];
  assign o[46386] = i[90];
  assign o[46387] = i[90];
  assign o[46388] = i[90];
  assign o[46389] = i[90];
  assign o[46390] = i[90];
  assign o[46391] = i[90];
  assign o[46392] = i[90];
  assign o[46393] = i[90];
  assign o[46394] = i[90];
  assign o[46395] = i[90];
  assign o[46396] = i[90];
  assign o[46397] = i[90];
  assign o[46398] = i[90];
  assign o[46399] = i[90];
  assign o[46400] = i[90];
  assign o[46401] = i[90];
  assign o[46402] = i[90];
  assign o[46403] = i[90];
  assign o[46404] = i[90];
  assign o[46405] = i[90];
  assign o[46406] = i[90];
  assign o[46407] = i[90];
  assign o[46408] = i[90];
  assign o[46409] = i[90];
  assign o[46410] = i[90];
  assign o[46411] = i[90];
  assign o[46412] = i[90];
  assign o[46413] = i[90];
  assign o[46414] = i[90];
  assign o[46415] = i[90];
  assign o[46416] = i[90];
  assign o[46417] = i[90];
  assign o[46418] = i[90];
  assign o[46419] = i[90];
  assign o[46420] = i[90];
  assign o[46421] = i[90];
  assign o[46422] = i[90];
  assign o[46423] = i[90];
  assign o[46424] = i[90];
  assign o[46425] = i[90];
  assign o[46426] = i[90];
  assign o[46427] = i[90];
  assign o[46428] = i[90];
  assign o[46429] = i[90];
  assign o[46430] = i[90];
  assign o[46431] = i[90];
  assign o[46432] = i[90];
  assign o[46433] = i[90];
  assign o[46434] = i[90];
  assign o[46435] = i[90];
  assign o[46436] = i[90];
  assign o[46437] = i[90];
  assign o[46438] = i[90];
  assign o[46439] = i[90];
  assign o[46440] = i[90];
  assign o[46441] = i[90];
  assign o[46442] = i[90];
  assign o[46443] = i[90];
  assign o[46444] = i[90];
  assign o[46445] = i[90];
  assign o[46446] = i[90];
  assign o[46447] = i[90];
  assign o[46448] = i[90];
  assign o[46449] = i[90];
  assign o[46450] = i[90];
  assign o[46451] = i[90];
  assign o[46452] = i[90];
  assign o[46453] = i[90];
  assign o[46454] = i[90];
  assign o[46455] = i[90];
  assign o[46456] = i[90];
  assign o[46457] = i[90];
  assign o[46458] = i[90];
  assign o[46459] = i[90];
  assign o[46460] = i[90];
  assign o[46461] = i[90];
  assign o[46462] = i[90];
  assign o[46463] = i[90];
  assign o[46464] = i[90];
  assign o[46465] = i[90];
  assign o[46466] = i[90];
  assign o[46467] = i[90];
  assign o[46468] = i[90];
  assign o[46469] = i[90];
  assign o[46470] = i[90];
  assign o[46471] = i[90];
  assign o[46472] = i[90];
  assign o[46473] = i[90];
  assign o[46474] = i[90];
  assign o[46475] = i[90];
  assign o[46476] = i[90];
  assign o[46477] = i[90];
  assign o[46478] = i[90];
  assign o[46479] = i[90];
  assign o[46480] = i[90];
  assign o[46481] = i[90];
  assign o[46482] = i[90];
  assign o[46483] = i[90];
  assign o[46484] = i[90];
  assign o[46485] = i[90];
  assign o[46486] = i[90];
  assign o[46487] = i[90];
  assign o[46488] = i[90];
  assign o[46489] = i[90];
  assign o[46490] = i[90];
  assign o[46491] = i[90];
  assign o[46492] = i[90];
  assign o[46493] = i[90];
  assign o[46494] = i[90];
  assign o[46495] = i[90];
  assign o[46496] = i[90];
  assign o[46497] = i[90];
  assign o[46498] = i[90];
  assign o[46499] = i[90];
  assign o[46500] = i[90];
  assign o[46501] = i[90];
  assign o[46502] = i[90];
  assign o[46503] = i[90];
  assign o[46504] = i[90];
  assign o[46505] = i[90];
  assign o[46506] = i[90];
  assign o[46507] = i[90];
  assign o[46508] = i[90];
  assign o[46509] = i[90];
  assign o[46510] = i[90];
  assign o[46511] = i[90];
  assign o[46512] = i[90];
  assign o[46513] = i[90];
  assign o[46514] = i[90];
  assign o[46515] = i[90];
  assign o[46516] = i[90];
  assign o[46517] = i[90];
  assign o[46518] = i[90];
  assign o[46519] = i[90];
  assign o[46520] = i[90];
  assign o[46521] = i[90];
  assign o[46522] = i[90];
  assign o[46523] = i[90];
  assign o[46524] = i[90];
  assign o[46525] = i[90];
  assign o[46526] = i[90];
  assign o[46527] = i[90];
  assign o[46528] = i[90];
  assign o[46529] = i[90];
  assign o[46530] = i[90];
  assign o[46531] = i[90];
  assign o[46532] = i[90];
  assign o[46533] = i[90];
  assign o[46534] = i[90];
  assign o[46535] = i[90];
  assign o[46536] = i[90];
  assign o[46537] = i[90];
  assign o[46538] = i[90];
  assign o[46539] = i[90];
  assign o[46540] = i[90];
  assign o[46541] = i[90];
  assign o[46542] = i[90];
  assign o[46543] = i[90];
  assign o[46544] = i[90];
  assign o[46545] = i[90];
  assign o[46546] = i[90];
  assign o[46547] = i[90];
  assign o[46548] = i[90];
  assign o[46549] = i[90];
  assign o[46550] = i[90];
  assign o[46551] = i[90];
  assign o[46552] = i[90];
  assign o[46553] = i[90];
  assign o[46554] = i[90];
  assign o[46555] = i[90];
  assign o[46556] = i[90];
  assign o[46557] = i[90];
  assign o[46558] = i[90];
  assign o[46559] = i[90];
  assign o[46560] = i[90];
  assign o[46561] = i[90];
  assign o[46562] = i[90];
  assign o[46563] = i[90];
  assign o[46564] = i[90];
  assign o[46565] = i[90];
  assign o[46566] = i[90];
  assign o[46567] = i[90];
  assign o[46568] = i[90];
  assign o[46569] = i[90];
  assign o[46570] = i[90];
  assign o[46571] = i[90];
  assign o[46572] = i[90];
  assign o[46573] = i[90];
  assign o[46574] = i[90];
  assign o[46575] = i[90];
  assign o[46576] = i[90];
  assign o[46577] = i[90];
  assign o[46578] = i[90];
  assign o[46579] = i[90];
  assign o[46580] = i[90];
  assign o[46581] = i[90];
  assign o[46582] = i[90];
  assign o[46583] = i[90];
  assign o[46584] = i[90];
  assign o[46585] = i[90];
  assign o[46586] = i[90];
  assign o[46587] = i[90];
  assign o[46588] = i[90];
  assign o[46589] = i[90];
  assign o[46590] = i[90];
  assign o[46591] = i[90];
  assign o[45568] = i[89];
  assign o[45569] = i[89];
  assign o[45570] = i[89];
  assign o[45571] = i[89];
  assign o[45572] = i[89];
  assign o[45573] = i[89];
  assign o[45574] = i[89];
  assign o[45575] = i[89];
  assign o[45576] = i[89];
  assign o[45577] = i[89];
  assign o[45578] = i[89];
  assign o[45579] = i[89];
  assign o[45580] = i[89];
  assign o[45581] = i[89];
  assign o[45582] = i[89];
  assign o[45583] = i[89];
  assign o[45584] = i[89];
  assign o[45585] = i[89];
  assign o[45586] = i[89];
  assign o[45587] = i[89];
  assign o[45588] = i[89];
  assign o[45589] = i[89];
  assign o[45590] = i[89];
  assign o[45591] = i[89];
  assign o[45592] = i[89];
  assign o[45593] = i[89];
  assign o[45594] = i[89];
  assign o[45595] = i[89];
  assign o[45596] = i[89];
  assign o[45597] = i[89];
  assign o[45598] = i[89];
  assign o[45599] = i[89];
  assign o[45600] = i[89];
  assign o[45601] = i[89];
  assign o[45602] = i[89];
  assign o[45603] = i[89];
  assign o[45604] = i[89];
  assign o[45605] = i[89];
  assign o[45606] = i[89];
  assign o[45607] = i[89];
  assign o[45608] = i[89];
  assign o[45609] = i[89];
  assign o[45610] = i[89];
  assign o[45611] = i[89];
  assign o[45612] = i[89];
  assign o[45613] = i[89];
  assign o[45614] = i[89];
  assign o[45615] = i[89];
  assign o[45616] = i[89];
  assign o[45617] = i[89];
  assign o[45618] = i[89];
  assign o[45619] = i[89];
  assign o[45620] = i[89];
  assign o[45621] = i[89];
  assign o[45622] = i[89];
  assign o[45623] = i[89];
  assign o[45624] = i[89];
  assign o[45625] = i[89];
  assign o[45626] = i[89];
  assign o[45627] = i[89];
  assign o[45628] = i[89];
  assign o[45629] = i[89];
  assign o[45630] = i[89];
  assign o[45631] = i[89];
  assign o[45632] = i[89];
  assign o[45633] = i[89];
  assign o[45634] = i[89];
  assign o[45635] = i[89];
  assign o[45636] = i[89];
  assign o[45637] = i[89];
  assign o[45638] = i[89];
  assign o[45639] = i[89];
  assign o[45640] = i[89];
  assign o[45641] = i[89];
  assign o[45642] = i[89];
  assign o[45643] = i[89];
  assign o[45644] = i[89];
  assign o[45645] = i[89];
  assign o[45646] = i[89];
  assign o[45647] = i[89];
  assign o[45648] = i[89];
  assign o[45649] = i[89];
  assign o[45650] = i[89];
  assign o[45651] = i[89];
  assign o[45652] = i[89];
  assign o[45653] = i[89];
  assign o[45654] = i[89];
  assign o[45655] = i[89];
  assign o[45656] = i[89];
  assign o[45657] = i[89];
  assign o[45658] = i[89];
  assign o[45659] = i[89];
  assign o[45660] = i[89];
  assign o[45661] = i[89];
  assign o[45662] = i[89];
  assign o[45663] = i[89];
  assign o[45664] = i[89];
  assign o[45665] = i[89];
  assign o[45666] = i[89];
  assign o[45667] = i[89];
  assign o[45668] = i[89];
  assign o[45669] = i[89];
  assign o[45670] = i[89];
  assign o[45671] = i[89];
  assign o[45672] = i[89];
  assign o[45673] = i[89];
  assign o[45674] = i[89];
  assign o[45675] = i[89];
  assign o[45676] = i[89];
  assign o[45677] = i[89];
  assign o[45678] = i[89];
  assign o[45679] = i[89];
  assign o[45680] = i[89];
  assign o[45681] = i[89];
  assign o[45682] = i[89];
  assign o[45683] = i[89];
  assign o[45684] = i[89];
  assign o[45685] = i[89];
  assign o[45686] = i[89];
  assign o[45687] = i[89];
  assign o[45688] = i[89];
  assign o[45689] = i[89];
  assign o[45690] = i[89];
  assign o[45691] = i[89];
  assign o[45692] = i[89];
  assign o[45693] = i[89];
  assign o[45694] = i[89];
  assign o[45695] = i[89];
  assign o[45696] = i[89];
  assign o[45697] = i[89];
  assign o[45698] = i[89];
  assign o[45699] = i[89];
  assign o[45700] = i[89];
  assign o[45701] = i[89];
  assign o[45702] = i[89];
  assign o[45703] = i[89];
  assign o[45704] = i[89];
  assign o[45705] = i[89];
  assign o[45706] = i[89];
  assign o[45707] = i[89];
  assign o[45708] = i[89];
  assign o[45709] = i[89];
  assign o[45710] = i[89];
  assign o[45711] = i[89];
  assign o[45712] = i[89];
  assign o[45713] = i[89];
  assign o[45714] = i[89];
  assign o[45715] = i[89];
  assign o[45716] = i[89];
  assign o[45717] = i[89];
  assign o[45718] = i[89];
  assign o[45719] = i[89];
  assign o[45720] = i[89];
  assign o[45721] = i[89];
  assign o[45722] = i[89];
  assign o[45723] = i[89];
  assign o[45724] = i[89];
  assign o[45725] = i[89];
  assign o[45726] = i[89];
  assign o[45727] = i[89];
  assign o[45728] = i[89];
  assign o[45729] = i[89];
  assign o[45730] = i[89];
  assign o[45731] = i[89];
  assign o[45732] = i[89];
  assign o[45733] = i[89];
  assign o[45734] = i[89];
  assign o[45735] = i[89];
  assign o[45736] = i[89];
  assign o[45737] = i[89];
  assign o[45738] = i[89];
  assign o[45739] = i[89];
  assign o[45740] = i[89];
  assign o[45741] = i[89];
  assign o[45742] = i[89];
  assign o[45743] = i[89];
  assign o[45744] = i[89];
  assign o[45745] = i[89];
  assign o[45746] = i[89];
  assign o[45747] = i[89];
  assign o[45748] = i[89];
  assign o[45749] = i[89];
  assign o[45750] = i[89];
  assign o[45751] = i[89];
  assign o[45752] = i[89];
  assign o[45753] = i[89];
  assign o[45754] = i[89];
  assign o[45755] = i[89];
  assign o[45756] = i[89];
  assign o[45757] = i[89];
  assign o[45758] = i[89];
  assign o[45759] = i[89];
  assign o[45760] = i[89];
  assign o[45761] = i[89];
  assign o[45762] = i[89];
  assign o[45763] = i[89];
  assign o[45764] = i[89];
  assign o[45765] = i[89];
  assign o[45766] = i[89];
  assign o[45767] = i[89];
  assign o[45768] = i[89];
  assign o[45769] = i[89];
  assign o[45770] = i[89];
  assign o[45771] = i[89];
  assign o[45772] = i[89];
  assign o[45773] = i[89];
  assign o[45774] = i[89];
  assign o[45775] = i[89];
  assign o[45776] = i[89];
  assign o[45777] = i[89];
  assign o[45778] = i[89];
  assign o[45779] = i[89];
  assign o[45780] = i[89];
  assign o[45781] = i[89];
  assign o[45782] = i[89];
  assign o[45783] = i[89];
  assign o[45784] = i[89];
  assign o[45785] = i[89];
  assign o[45786] = i[89];
  assign o[45787] = i[89];
  assign o[45788] = i[89];
  assign o[45789] = i[89];
  assign o[45790] = i[89];
  assign o[45791] = i[89];
  assign o[45792] = i[89];
  assign o[45793] = i[89];
  assign o[45794] = i[89];
  assign o[45795] = i[89];
  assign o[45796] = i[89];
  assign o[45797] = i[89];
  assign o[45798] = i[89];
  assign o[45799] = i[89];
  assign o[45800] = i[89];
  assign o[45801] = i[89];
  assign o[45802] = i[89];
  assign o[45803] = i[89];
  assign o[45804] = i[89];
  assign o[45805] = i[89];
  assign o[45806] = i[89];
  assign o[45807] = i[89];
  assign o[45808] = i[89];
  assign o[45809] = i[89];
  assign o[45810] = i[89];
  assign o[45811] = i[89];
  assign o[45812] = i[89];
  assign o[45813] = i[89];
  assign o[45814] = i[89];
  assign o[45815] = i[89];
  assign o[45816] = i[89];
  assign o[45817] = i[89];
  assign o[45818] = i[89];
  assign o[45819] = i[89];
  assign o[45820] = i[89];
  assign o[45821] = i[89];
  assign o[45822] = i[89];
  assign o[45823] = i[89];
  assign o[45824] = i[89];
  assign o[45825] = i[89];
  assign o[45826] = i[89];
  assign o[45827] = i[89];
  assign o[45828] = i[89];
  assign o[45829] = i[89];
  assign o[45830] = i[89];
  assign o[45831] = i[89];
  assign o[45832] = i[89];
  assign o[45833] = i[89];
  assign o[45834] = i[89];
  assign o[45835] = i[89];
  assign o[45836] = i[89];
  assign o[45837] = i[89];
  assign o[45838] = i[89];
  assign o[45839] = i[89];
  assign o[45840] = i[89];
  assign o[45841] = i[89];
  assign o[45842] = i[89];
  assign o[45843] = i[89];
  assign o[45844] = i[89];
  assign o[45845] = i[89];
  assign o[45846] = i[89];
  assign o[45847] = i[89];
  assign o[45848] = i[89];
  assign o[45849] = i[89];
  assign o[45850] = i[89];
  assign o[45851] = i[89];
  assign o[45852] = i[89];
  assign o[45853] = i[89];
  assign o[45854] = i[89];
  assign o[45855] = i[89];
  assign o[45856] = i[89];
  assign o[45857] = i[89];
  assign o[45858] = i[89];
  assign o[45859] = i[89];
  assign o[45860] = i[89];
  assign o[45861] = i[89];
  assign o[45862] = i[89];
  assign o[45863] = i[89];
  assign o[45864] = i[89];
  assign o[45865] = i[89];
  assign o[45866] = i[89];
  assign o[45867] = i[89];
  assign o[45868] = i[89];
  assign o[45869] = i[89];
  assign o[45870] = i[89];
  assign o[45871] = i[89];
  assign o[45872] = i[89];
  assign o[45873] = i[89];
  assign o[45874] = i[89];
  assign o[45875] = i[89];
  assign o[45876] = i[89];
  assign o[45877] = i[89];
  assign o[45878] = i[89];
  assign o[45879] = i[89];
  assign o[45880] = i[89];
  assign o[45881] = i[89];
  assign o[45882] = i[89];
  assign o[45883] = i[89];
  assign o[45884] = i[89];
  assign o[45885] = i[89];
  assign o[45886] = i[89];
  assign o[45887] = i[89];
  assign o[45888] = i[89];
  assign o[45889] = i[89];
  assign o[45890] = i[89];
  assign o[45891] = i[89];
  assign o[45892] = i[89];
  assign o[45893] = i[89];
  assign o[45894] = i[89];
  assign o[45895] = i[89];
  assign o[45896] = i[89];
  assign o[45897] = i[89];
  assign o[45898] = i[89];
  assign o[45899] = i[89];
  assign o[45900] = i[89];
  assign o[45901] = i[89];
  assign o[45902] = i[89];
  assign o[45903] = i[89];
  assign o[45904] = i[89];
  assign o[45905] = i[89];
  assign o[45906] = i[89];
  assign o[45907] = i[89];
  assign o[45908] = i[89];
  assign o[45909] = i[89];
  assign o[45910] = i[89];
  assign o[45911] = i[89];
  assign o[45912] = i[89];
  assign o[45913] = i[89];
  assign o[45914] = i[89];
  assign o[45915] = i[89];
  assign o[45916] = i[89];
  assign o[45917] = i[89];
  assign o[45918] = i[89];
  assign o[45919] = i[89];
  assign o[45920] = i[89];
  assign o[45921] = i[89];
  assign o[45922] = i[89];
  assign o[45923] = i[89];
  assign o[45924] = i[89];
  assign o[45925] = i[89];
  assign o[45926] = i[89];
  assign o[45927] = i[89];
  assign o[45928] = i[89];
  assign o[45929] = i[89];
  assign o[45930] = i[89];
  assign o[45931] = i[89];
  assign o[45932] = i[89];
  assign o[45933] = i[89];
  assign o[45934] = i[89];
  assign o[45935] = i[89];
  assign o[45936] = i[89];
  assign o[45937] = i[89];
  assign o[45938] = i[89];
  assign o[45939] = i[89];
  assign o[45940] = i[89];
  assign o[45941] = i[89];
  assign o[45942] = i[89];
  assign o[45943] = i[89];
  assign o[45944] = i[89];
  assign o[45945] = i[89];
  assign o[45946] = i[89];
  assign o[45947] = i[89];
  assign o[45948] = i[89];
  assign o[45949] = i[89];
  assign o[45950] = i[89];
  assign o[45951] = i[89];
  assign o[45952] = i[89];
  assign o[45953] = i[89];
  assign o[45954] = i[89];
  assign o[45955] = i[89];
  assign o[45956] = i[89];
  assign o[45957] = i[89];
  assign o[45958] = i[89];
  assign o[45959] = i[89];
  assign o[45960] = i[89];
  assign o[45961] = i[89];
  assign o[45962] = i[89];
  assign o[45963] = i[89];
  assign o[45964] = i[89];
  assign o[45965] = i[89];
  assign o[45966] = i[89];
  assign o[45967] = i[89];
  assign o[45968] = i[89];
  assign o[45969] = i[89];
  assign o[45970] = i[89];
  assign o[45971] = i[89];
  assign o[45972] = i[89];
  assign o[45973] = i[89];
  assign o[45974] = i[89];
  assign o[45975] = i[89];
  assign o[45976] = i[89];
  assign o[45977] = i[89];
  assign o[45978] = i[89];
  assign o[45979] = i[89];
  assign o[45980] = i[89];
  assign o[45981] = i[89];
  assign o[45982] = i[89];
  assign o[45983] = i[89];
  assign o[45984] = i[89];
  assign o[45985] = i[89];
  assign o[45986] = i[89];
  assign o[45987] = i[89];
  assign o[45988] = i[89];
  assign o[45989] = i[89];
  assign o[45990] = i[89];
  assign o[45991] = i[89];
  assign o[45992] = i[89];
  assign o[45993] = i[89];
  assign o[45994] = i[89];
  assign o[45995] = i[89];
  assign o[45996] = i[89];
  assign o[45997] = i[89];
  assign o[45998] = i[89];
  assign o[45999] = i[89];
  assign o[46000] = i[89];
  assign o[46001] = i[89];
  assign o[46002] = i[89];
  assign o[46003] = i[89];
  assign o[46004] = i[89];
  assign o[46005] = i[89];
  assign o[46006] = i[89];
  assign o[46007] = i[89];
  assign o[46008] = i[89];
  assign o[46009] = i[89];
  assign o[46010] = i[89];
  assign o[46011] = i[89];
  assign o[46012] = i[89];
  assign o[46013] = i[89];
  assign o[46014] = i[89];
  assign o[46015] = i[89];
  assign o[46016] = i[89];
  assign o[46017] = i[89];
  assign o[46018] = i[89];
  assign o[46019] = i[89];
  assign o[46020] = i[89];
  assign o[46021] = i[89];
  assign o[46022] = i[89];
  assign o[46023] = i[89];
  assign o[46024] = i[89];
  assign o[46025] = i[89];
  assign o[46026] = i[89];
  assign o[46027] = i[89];
  assign o[46028] = i[89];
  assign o[46029] = i[89];
  assign o[46030] = i[89];
  assign o[46031] = i[89];
  assign o[46032] = i[89];
  assign o[46033] = i[89];
  assign o[46034] = i[89];
  assign o[46035] = i[89];
  assign o[46036] = i[89];
  assign o[46037] = i[89];
  assign o[46038] = i[89];
  assign o[46039] = i[89];
  assign o[46040] = i[89];
  assign o[46041] = i[89];
  assign o[46042] = i[89];
  assign o[46043] = i[89];
  assign o[46044] = i[89];
  assign o[46045] = i[89];
  assign o[46046] = i[89];
  assign o[46047] = i[89];
  assign o[46048] = i[89];
  assign o[46049] = i[89];
  assign o[46050] = i[89];
  assign o[46051] = i[89];
  assign o[46052] = i[89];
  assign o[46053] = i[89];
  assign o[46054] = i[89];
  assign o[46055] = i[89];
  assign o[46056] = i[89];
  assign o[46057] = i[89];
  assign o[46058] = i[89];
  assign o[46059] = i[89];
  assign o[46060] = i[89];
  assign o[46061] = i[89];
  assign o[46062] = i[89];
  assign o[46063] = i[89];
  assign o[46064] = i[89];
  assign o[46065] = i[89];
  assign o[46066] = i[89];
  assign o[46067] = i[89];
  assign o[46068] = i[89];
  assign o[46069] = i[89];
  assign o[46070] = i[89];
  assign o[46071] = i[89];
  assign o[46072] = i[89];
  assign o[46073] = i[89];
  assign o[46074] = i[89];
  assign o[46075] = i[89];
  assign o[46076] = i[89];
  assign o[46077] = i[89];
  assign o[46078] = i[89];
  assign o[46079] = i[89];
  assign o[45056] = i[88];
  assign o[45057] = i[88];
  assign o[45058] = i[88];
  assign o[45059] = i[88];
  assign o[45060] = i[88];
  assign o[45061] = i[88];
  assign o[45062] = i[88];
  assign o[45063] = i[88];
  assign o[45064] = i[88];
  assign o[45065] = i[88];
  assign o[45066] = i[88];
  assign o[45067] = i[88];
  assign o[45068] = i[88];
  assign o[45069] = i[88];
  assign o[45070] = i[88];
  assign o[45071] = i[88];
  assign o[45072] = i[88];
  assign o[45073] = i[88];
  assign o[45074] = i[88];
  assign o[45075] = i[88];
  assign o[45076] = i[88];
  assign o[45077] = i[88];
  assign o[45078] = i[88];
  assign o[45079] = i[88];
  assign o[45080] = i[88];
  assign o[45081] = i[88];
  assign o[45082] = i[88];
  assign o[45083] = i[88];
  assign o[45084] = i[88];
  assign o[45085] = i[88];
  assign o[45086] = i[88];
  assign o[45087] = i[88];
  assign o[45088] = i[88];
  assign o[45089] = i[88];
  assign o[45090] = i[88];
  assign o[45091] = i[88];
  assign o[45092] = i[88];
  assign o[45093] = i[88];
  assign o[45094] = i[88];
  assign o[45095] = i[88];
  assign o[45096] = i[88];
  assign o[45097] = i[88];
  assign o[45098] = i[88];
  assign o[45099] = i[88];
  assign o[45100] = i[88];
  assign o[45101] = i[88];
  assign o[45102] = i[88];
  assign o[45103] = i[88];
  assign o[45104] = i[88];
  assign o[45105] = i[88];
  assign o[45106] = i[88];
  assign o[45107] = i[88];
  assign o[45108] = i[88];
  assign o[45109] = i[88];
  assign o[45110] = i[88];
  assign o[45111] = i[88];
  assign o[45112] = i[88];
  assign o[45113] = i[88];
  assign o[45114] = i[88];
  assign o[45115] = i[88];
  assign o[45116] = i[88];
  assign o[45117] = i[88];
  assign o[45118] = i[88];
  assign o[45119] = i[88];
  assign o[45120] = i[88];
  assign o[45121] = i[88];
  assign o[45122] = i[88];
  assign o[45123] = i[88];
  assign o[45124] = i[88];
  assign o[45125] = i[88];
  assign o[45126] = i[88];
  assign o[45127] = i[88];
  assign o[45128] = i[88];
  assign o[45129] = i[88];
  assign o[45130] = i[88];
  assign o[45131] = i[88];
  assign o[45132] = i[88];
  assign o[45133] = i[88];
  assign o[45134] = i[88];
  assign o[45135] = i[88];
  assign o[45136] = i[88];
  assign o[45137] = i[88];
  assign o[45138] = i[88];
  assign o[45139] = i[88];
  assign o[45140] = i[88];
  assign o[45141] = i[88];
  assign o[45142] = i[88];
  assign o[45143] = i[88];
  assign o[45144] = i[88];
  assign o[45145] = i[88];
  assign o[45146] = i[88];
  assign o[45147] = i[88];
  assign o[45148] = i[88];
  assign o[45149] = i[88];
  assign o[45150] = i[88];
  assign o[45151] = i[88];
  assign o[45152] = i[88];
  assign o[45153] = i[88];
  assign o[45154] = i[88];
  assign o[45155] = i[88];
  assign o[45156] = i[88];
  assign o[45157] = i[88];
  assign o[45158] = i[88];
  assign o[45159] = i[88];
  assign o[45160] = i[88];
  assign o[45161] = i[88];
  assign o[45162] = i[88];
  assign o[45163] = i[88];
  assign o[45164] = i[88];
  assign o[45165] = i[88];
  assign o[45166] = i[88];
  assign o[45167] = i[88];
  assign o[45168] = i[88];
  assign o[45169] = i[88];
  assign o[45170] = i[88];
  assign o[45171] = i[88];
  assign o[45172] = i[88];
  assign o[45173] = i[88];
  assign o[45174] = i[88];
  assign o[45175] = i[88];
  assign o[45176] = i[88];
  assign o[45177] = i[88];
  assign o[45178] = i[88];
  assign o[45179] = i[88];
  assign o[45180] = i[88];
  assign o[45181] = i[88];
  assign o[45182] = i[88];
  assign o[45183] = i[88];
  assign o[45184] = i[88];
  assign o[45185] = i[88];
  assign o[45186] = i[88];
  assign o[45187] = i[88];
  assign o[45188] = i[88];
  assign o[45189] = i[88];
  assign o[45190] = i[88];
  assign o[45191] = i[88];
  assign o[45192] = i[88];
  assign o[45193] = i[88];
  assign o[45194] = i[88];
  assign o[45195] = i[88];
  assign o[45196] = i[88];
  assign o[45197] = i[88];
  assign o[45198] = i[88];
  assign o[45199] = i[88];
  assign o[45200] = i[88];
  assign o[45201] = i[88];
  assign o[45202] = i[88];
  assign o[45203] = i[88];
  assign o[45204] = i[88];
  assign o[45205] = i[88];
  assign o[45206] = i[88];
  assign o[45207] = i[88];
  assign o[45208] = i[88];
  assign o[45209] = i[88];
  assign o[45210] = i[88];
  assign o[45211] = i[88];
  assign o[45212] = i[88];
  assign o[45213] = i[88];
  assign o[45214] = i[88];
  assign o[45215] = i[88];
  assign o[45216] = i[88];
  assign o[45217] = i[88];
  assign o[45218] = i[88];
  assign o[45219] = i[88];
  assign o[45220] = i[88];
  assign o[45221] = i[88];
  assign o[45222] = i[88];
  assign o[45223] = i[88];
  assign o[45224] = i[88];
  assign o[45225] = i[88];
  assign o[45226] = i[88];
  assign o[45227] = i[88];
  assign o[45228] = i[88];
  assign o[45229] = i[88];
  assign o[45230] = i[88];
  assign o[45231] = i[88];
  assign o[45232] = i[88];
  assign o[45233] = i[88];
  assign o[45234] = i[88];
  assign o[45235] = i[88];
  assign o[45236] = i[88];
  assign o[45237] = i[88];
  assign o[45238] = i[88];
  assign o[45239] = i[88];
  assign o[45240] = i[88];
  assign o[45241] = i[88];
  assign o[45242] = i[88];
  assign o[45243] = i[88];
  assign o[45244] = i[88];
  assign o[45245] = i[88];
  assign o[45246] = i[88];
  assign o[45247] = i[88];
  assign o[45248] = i[88];
  assign o[45249] = i[88];
  assign o[45250] = i[88];
  assign o[45251] = i[88];
  assign o[45252] = i[88];
  assign o[45253] = i[88];
  assign o[45254] = i[88];
  assign o[45255] = i[88];
  assign o[45256] = i[88];
  assign o[45257] = i[88];
  assign o[45258] = i[88];
  assign o[45259] = i[88];
  assign o[45260] = i[88];
  assign o[45261] = i[88];
  assign o[45262] = i[88];
  assign o[45263] = i[88];
  assign o[45264] = i[88];
  assign o[45265] = i[88];
  assign o[45266] = i[88];
  assign o[45267] = i[88];
  assign o[45268] = i[88];
  assign o[45269] = i[88];
  assign o[45270] = i[88];
  assign o[45271] = i[88];
  assign o[45272] = i[88];
  assign o[45273] = i[88];
  assign o[45274] = i[88];
  assign o[45275] = i[88];
  assign o[45276] = i[88];
  assign o[45277] = i[88];
  assign o[45278] = i[88];
  assign o[45279] = i[88];
  assign o[45280] = i[88];
  assign o[45281] = i[88];
  assign o[45282] = i[88];
  assign o[45283] = i[88];
  assign o[45284] = i[88];
  assign o[45285] = i[88];
  assign o[45286] = i[88];
  assign o[45287] = i[88];
  assign o[45288] = i[88];
  assign o[45289] = i[88];
  assign o[45290] = i[88];
  assign o[45291] = i[88];
  assign o[45292] = i[88];
  assign o[45293] = i[88];
  assign o[45294] = i[88];
  assign o[45295] = i[88];
  assign o[45296] = i[88];
  assign o[45297] = i[88];
  assign o[45298] = i[88];
  assign o[45299] = i[88];
  assign o[45300] = i[88];
  assign o[45301] = i[88];
  assign o[45302] = i[88];
  assign o[45303] = i[88];
  assign o[45304] = i[88];
  assign o[45305] = i[88];
  assign o[45306] = i[88];
  assign o[45307] = i[88];
  assign o[45308] = i[88];
  assign o[45309] = i[88];
  assign o[45310] = i[88];
  assign o[45311] = i[88];
  assign o[45312] = i[88];
  assign o[45313] = i[88];
  assign o[45314] = i[88];
  assign o[45315] = i[88];
  assign o[45316] = i[88];
  assign o[45317] = i[88];
  assign o[45318] = i[88];
  assign o[45319] = i[88];
  assign o[45320] = i[88];
  assign o[45321] = i[88];
  assign o[45322] = i[88];
  assign o[45323] = i[88];
  assign o[45324] = i[88];
  assign o[45325] = i[88];
  assign o[45326] = i[88];
  assign o[45327] = i[88];
  assign o[45328] = i[88];
  assign o[45329] = i[88];
  assign o[45330] = i[88];
  assign o[45331] = i[88];
  assign o[45332] = i[88];
  assign o[45333] = i[88];
  assign o[45334] = i[88];
  assign o[45335] = i[88];
  assign o[45336] = i[88];
  assign o[45337] = i[88];
  assign o[45338] = i[88];
  assign o[45339] = i[88];
  assign o[45340] = i[88];
  assign o[45341] = i[88];
  assign o[45342] = i[88];
  assign o[45343] = i[88];
  assign o[45344] = i[88];
  assign o[45345] = i[88];
  assign o[45346] = i[88];
  assign o[45347] = i[88];
  assign o[45348] = i[88];
  assign o[45349] = i[88];
  assign o[45350] = i[88];
  assign o[45351] = i[88];
  assign o[45352] = i[88];
  assign o[45353] = i[88];
  assign o[45354] = i[88];
  assign o[45355] = i[88];
  assign o[45356] = i[88];
  assign o[45357] = i[88];
  assign o[45358] = i[88];
  assign o[45359] = i[88];
  assign o[45360] = i[88];
  assign o[45361] = i[88];
  assign o[45362] = i[88];
  assign o[45363] = i[88];
  assign o[45364] = i[88];
  assign o[45365] = i[88];
  assign o[45366] = i[88];
  assign o[45367] = i[88];
  assign o[45368] = i[88];
  assign o[45369] = i[88];
  assign o[45370] = i[88];
  assign o[45371] = i[88];
  assign o[45372] = i[88];
  assign o[45373] = i[88];
  assign o[45374] = i[88];
  assign o[45375] = i[88];
  assign o[45376] = i[88];
  assign o[45377] = i[88];
  assign o[45378] = i[88];
  assign o[45379] = i[88];
  assign o[45380] = i[88];
  assign o[45381] = i[88];
  assign o[45382] = i[88];
  assign o[45383] = i[88];
  assign o[45384] = i[88];
  assign o[45385] = i[88];
  assign o[45386] = i[88];
  assign o[45387] = i[88];
  assign o[45388] = i[88];
  assign o[45389] = i[88];
  assign o[45390] = i[88];
  assign o[45391] = i[88];
  assign o[45392] = i[88];
  assign o[45393] = i[88];
  assign o[45394] = i[88];
  assign o[45395] = i[88];
  assign o[45396] = i[88];
  assign o[45397] = i[88];
  assign o[45398] = i[88];
  assign o[45399] = i[88];
  assign o[45400] = i[88];
  assign o[45401] = i[88];
  assign o[45402] = i[88];
  assign o[45403] = i[88];
  assign o[45404] = i[88];
  assign o[45405] = i[88];
  assign o[45406] = i[88];
  assign o[45407] = i[88];
  assign o[45408] = i[88];
  assign o[45409] = i[88];
  assign o[45410] = i[88];
  assign o[45411] = i[88];
  assign o[45412] = i[88];
  assign o[45413] = i[88];
  assign o[45414] = i[88];
  assign o[45415] = i[88];
  assign o[45416] = i[88];
  assign o[45417] = i[88];
  assign o[45418] = i[88];
  assign o[45419] = i[88];
  assign o[45420] = i[88];
  assign o[45421] = i[88];
  assign o[45422] = i[88];
  assign o[45423] = i[88];
  assign o[45424] = i[88];
  assign o[45425] = i[88];
  assign o[45426] = i[88];
  assign o[45427] = i[88];
  assign o[45428] = i[88];
  assign o[45429] = i[88];
  assign o[45430] = i[88];
  assign o[45431] = i[88];
  assign o[45432] = i[88];
  assign o[45433] = i[88];
  assign o[45434] = i[88];
  assign o[45435] = i[88];
  assign o[45436] = i[88];
  assign o[45437] = i[88];
  assign o[45438] = i[88];
  assign o[45439] = i[88];
  assign o[45440] = i[88];
  assign o[45441] = i[88];
  assign o[45442] = i[88];
  assign o[45443] = i[88];
  assign o[45444] = i[88];
  assign o[45445] = i[88];
  assign o[45446] = i[88];
  assign o[45447] = i[88];
  assign o[45448] = i[88];
  assign o[45449] = i[88];
  assign o[45450] = i[88];
  assign o[45451] = i[88];
  assign o[45452] = i[88];
  assign o[45453] = i[88];
  assign o[45454] = i[88];
  assign o[45455] = i[88];
  assign o[45456] = i[88];
  assign o[45457] = i[88];
  assign o[45458] = i[88];
  assign o[45459] = i[88];
  assign o[45460] = i[88];
  assign o[45461] = i[88];
  assign o[45462] = i[88];
  assign o[45463] = i[88];
  assign o[45464] = i[88];
  assign o[45465] = i[88];
  assign o[45466] = i[88];
  assign o[45467] = i[88];
  assign o[45468] = i[88];
  assign o[45469] = i[88];
  assign o[45470] = i[88];
  assign o[45471] = i[88];
  assign o[45472] = i[88];
  assign o[45473] = i[88];
  assign o[45474] = i[88];
  assign o[45475] = i[88];
  assign o[45476] = i[88];
  assign o[45477] = i[88];
  assign o[45478] = i[88];
  assign o[45479] = i[88];
  assign o[45480] = i[88];
  assign o[45481] = i[88];
  assign o[45482] = i[88];
  assign o[45483] = i[88];
  assign o[45484] = i[88];
  assign o[45485] = i[88];
  assign o[45486] = i[88];
  assign o[45487] = i[88];
  assign o[45488] = i[88];
  assign o[45489] = i[88];
  assign o[45490] = i[88];
  assign o[45491] = i[88];
  assign o[45492] = i[88];
  assign o[45493] = i[88];
  assign o[45494] = i[88];
  assign o[45495] = i[88];
  assign o[45496] = i[88];
  assign o[45497] = i[88];
  assign o[45498] = i[88];
  assign o[45499] = i[88];
  assign o[45500] = i[88];
  assign o[45501] = i[88];
  assign o[45502] = i[88];
  assign o[45503] = i[88];
  assign o[45504] = i[88];
  assign o[45505] = i[88];
  assign o[45506] = i[88];
  assign o[45507] = i[88];
  assign o[45508] = i[88];
  assign o[45509] = i[88];
  assign o[45510] = i[88];
  assign o[45511] = i[88];
  assign o[45512] = i[88];
  assign o[45513] = i[88];
  assign o[45514] = i[88];
  assign o[45515] = i[88];
  assign o[45516] = i[88];
  assign o[45517] = i[88];
  assign o[45518] = i[88];
  assign o[45519] = i[88];
  assign o[45520] = i[88];
  assign o[45521] = i[88];
  assign o[45522] = i[88];
  assign o[45523] = i[88];
  assign o[45524] = i[88];
  assign o[45525] = i[88];
  assign o[45526] = i[88];
  assign o[45527] = i[88];
  assign o[45528] = i[88];
  assign o[45529] = i[88];
  assign o[45530] = i[88];
  assign o[45531] = i[88];
  assign o[45532] = i[88];
  assign o[45533] = i[88];
  assign o[45534] = i[88];
  assign o[45535] = i[88];
  assign o[45536] = i[88];
  assign o[45537] = i[88];
  assign o[45538] = i[88];
  assign o[45539] = i[88];
  assign o[45540] = i[88];
  assign o[45541] = i[88];
  assign o[45542] = i[88];
  assign o[45543] = i[88];
  assign o[45544] = i[88];
  assign o[45545] = i[88];
  assign o[45546] = i[88];
  assign o[45547] = i[88];
  assign o[45548] = i[88];
  assign o[45549] = i[88];
  assign o[45550] = i[88];
  assign o[45551] = i[88];
  assign o[45552] = i[88];
  assign o[45553] = i[88];
  assign o[45554] = i[88];
  assign o[45555] = i[88];
  assign o[45556] = i[88];
  assign o[45557] = i[88];
  assign o[45558] = i[88];
  assign o[45559] = i[88];
  assign o[45560] = i[88];
  assign o[45561] = i[88];
  assign o[45562] = i[88];
  assign o[45563] = i[88];
  assign o[45564] = i[88];
  assign o[45565] = i[88];
  assign o[45566] = i[88];
  assign o[45567] = i[88];
  assign o[44544] = i[87];
  assign o[44545] = i[87];
  assign o[44546] = i[87];
  assign o[44547] = i[87];
  assign o[44548] = i[87];
  assign o[44549] = i[87];
  assign o[44550] = i[87];
  assign o[44551] = i[87];
  assign o[44552] = i[87];
  assign o[44553] = i[87];
  assign o[44554] = i[87];
  assign o[44555] = i[87];
  assign o[44556] = i[87];
  assign o[44557] = i[87];
  assign o[44558] = i[87];
  assign o[44559] = i[87];
  assign o[44560] = i[87];
  assign o[44561] = i[87];
  assign o[44562] = i[87];
  assign o[44563] = i[87];
  assign o[44564] = i[87];
  assign o[44565] = i[87];
  assign o[44566] = i[87];
  assign o[44567] = i[87];
  assign o[44568] = i[87];
  assign o[44569] = i[87];
  assign o[44570] = i[87];
  assign o[44571] = i[87];
  assign o[44572] = i[87];
  assign o[44573] = i[87];
  assign o[44574] = i[87];
  assign o[44575] = i[87];
  assign o[44576] = i[87];
  assign o[44577] = i[87];
  assign o[44578] = i[87];
  assign o[44579] = i[87];
  assign o[44580] = i[87];
  assign o[44581] = i[87];
  assign o[44582] = i[87];
  assign o[44583] = i[87];
  assign o[44584] = i[87];
  assign o[44585] = i[87];
  assign o[44586] = i[87];
  assign o[44587] = i[87];
  assign o[44588] = i[87];
  assign o[44589] = i[87];
  assign o[44590] = i[87];
  assign o[44591] = i[87];
  assign o[44592] = i[87];
  assign o[44593] = i[87];
  assign o[44594] = i[87];
  assign o[44595] = i[87];
  assign o[44596] = i[87];
  assign o[44597] = i[87];
  assign o[44598] = i[87];
  assign o[44599] = i[87];
  assign o[44600] = i[87];
  assign o[44601] = i[87];
  assign o[44602] = i[87];
  assign o[44603] = i[87];
  assign o[44604] = i[87];
  assign o[44605] = i[87];
  assign o[44606] = i[87];
  assign o[44607] = i[87];
  assign o[44608] = i[87];
  assign o[44609] = i[87];
  assign o[44610] = i[87];
  assign o[44611] = i[87];
  assign o[44612] = i[87];
  assign o[44613] = i[87];
  assign o[44614] = i[87];
  assign o[44615] = i[87];
  assign o[44616] = i[87];
  assign o[44617] = i[87];
  assign o[44618] = i[87];
  assign o[44619] = i[87];
  assign o[44620] = i[87];
  assign o[44621] = i[87];
  assign o[44622] = i[87];
  assign o[44623] = i[87];
  assign o[44624] = i[87];
  assign o[44625] = i[87];
  assign o[44626] = i[87];
  assign o[44627] = i[87];
  assign o[44628] = i[87];
  assign o[44629] = i[87];
  assign o[44630] = i[87];
  assign o[44631] = i[87];
  assign o[44632] = i[87];
  assign o[44633] = i[87];
  assign o[44634] = i[87];
  assign o[44635] = i[87];
  assign o[44636] = i[87];
  assign o[44637] = i[87];
  assign o[44638] = i[87];
  assign o[44639] = i[87];
  assign o[44640] = i[87];
  assign o[44641] = i[87];
  assign o[44642] = i[87];
  assign o[44643] = i[87];
  assign o[44644] = i[87];
  assign o[44645] = i[87];
  assign o[44646] = i[87];
  assign o[44647] = i[87];
  assign o[44648] = i[87];
  assign o[44649] = i[87];
  assign o[44650] = i[87];
  assign o[44651] = i[87];
  assign o[44652] = i[87];
  assign o[44653] = i[87];
  assign o[44654] = i[87];
  assign o[44655] = i[87];
  assign o[44656] = i[87];
  assign o[44657] = i[87];
  assign o[44658] = i[87];
  assign o[44659] = i[87];
  assign o[44660] = i[87];
  assign o[44661] = i[87];
  assign o[44662] = i[87];
  assign o[44663] = i[87];
  assign o[44664] = i[87];
  assign o[44665] = i[87];
  assign o[44666] = i[87];
  assign o[44667] = i[87];
  assign o[44668] = i[87];
  assign o[44669] = i[87];
  assign o[44670] = i[87];
  assign o[44671] = i[87];
  assign o[44672] = i[87];
  assign o[44673] = i[87];
  assign o[44674] = i[87];
  assign o[44675] = i[87];
  assign o[44676] = i[87];
  assign o[44677] = i[87];
  assign o[44678] = i[87];
  assign o[44679] = i[87];
  assign o[44680] = i[87];
  assign o[44681] = i[87];
  assign o[44682] = i[87];
  assign o[44683] = i[87];
  assign o[44684] = i[87];
  assign o[44685] = i[87];
  assign o[44686] = i[87];
  assign o[44687] = i[87];
  assign o[44688] = i[87];
  assign o[44689] = i[87];
  assign o[44690] = i[87];
  assign o[44691] = i[87];
  assign o[44692] = i[87];
  assign o[44693] = i[87];
  assign o[44694] = i[87];
  assign o[44695] = i[87];
  assign o[44696] = i[87];
  assign o[44697] = i[87];
  assign o[44698] = i[87];
  assign o[44699] = i[87];
  assign o[44700] = i[87];
  assign o[44701] = i[87];
  assign o[44702] = i[87];
  assign o[44703] = i[87];
  assign o[44704] = i[87];
  assign o[44705] = i[87];
  assign o[44706] = i[87];
  assign o[44707] = i[87];
  assign o[44708] = i[87];
  assign o[44709] = i[87];
  assign o[44710] = i[87];
  assign o[44711] = i[87];
  assign o[44712] = i[87];
  assign o[44713] = i[87];
  assign o[44714] = i[87];
  assign o[44715] = i[87];
  assign o[44716] = i[87];
  assign o[44717] = i[87];
  assign o[44718] = i[87];
  assign o[44719] = i[87];
  assign o[44720] = i[87];
  assign o[44721] = i[87];
  assign o[44722] = i[87];
  assign o[44723] = i[87];
  assign o[44724] = i[87];
  assign o[44725] = i[87];
  assign o[44726] = i[87];
  assign o[44727] = i[87];
  assign o[44728] = i[87];
  assign o[44729] = i[87];
  assign o[44730] = i[87];
  assign o[44731] = i[87];
  assign o[44732] = i[87];
  assign o[44733] = i[87];
  assign o[44734] = i[87];
  assign o[44735] = i[87];
  assign o[44736] = i[87];
  assign o[44737] = i[87];
  assign o[44738] = i[87];
  assign o[44739] = i[87];
  assign o[44740] = i[87];
  assign o[44741] = i[87];
  assign o[44742] = i[87];
  assign o[44743] = i[87];
  assign o[44744] = i[87];
  assign o[44745] = i[87];
  assign o[44746] = i[87];
  assign o[44747] = i[87];
  assign o[44748] = i[87];
  assign o[44749] = i[87];
  assign o[44750] = i[87];
  assign o[44751] = i[87];
  assign o[44752] = i[87];
  assign o[44753] = i[87];
  assign o[44754] = i[87];
  assign o[44755] = i[87];
  assign o[44756] = i[87];
  assign o[44757] = i[87];
  assign o[44758] = i[87];
  assign o[44759] = i[87];
  assign o[44760] = i[87];
  assign o[44761] = i[87];
  assign o[44762] = i[87];
  assign o[44763] = i[87];
  assign o[44764] = i[87];
  assign o[44765] = i[87];
  assign o[44766] = i[87];
  assign o[44767] = i[87];
  assign o[44768] = i[87];
  assign o[44769] = i[87];
  assign o[44770] = i[87];
  assign o[44771] = i[87];
  assign o[44772] = i[87];
  assign o[44773] = i[87];
  assign o[44774] = i[87];
  assign o[44775] = i[87];
  assign o[44776] = i[87];
  assign o[44777] = i[87];
  assign o[44778] = i[87];
  assign o[44779] = i[87];
  assign o[44780] = i[87];
  assign o[44781] = i[87];
  assign o[44782] = i[87];
  assign o[44783] = i[87];
  assign o[44784] = i[87];
  assign o[44785] = i[87];
  assign o[44786] = i[87];
  assign o[44787] = i[87];
  assign o[44788] = i[87];
  assign o[44789] = i[87];
  assign o[44790] = i[87];
  assign o[44791] = i[87];
  assign o[44792] = i[87];
  assign o[44793] = i[87];
  assign o[44794] = i[87];
  assign o[44795] = i[87];
  assign o[44796] = i[87];
  assign o[44797] = i[87];
  assign o[44798] = i[87];
  assign o[44799] = i[87];
  assign o[44800] = i[87];
  assign o[44801] = i[87];
  assign o[44802] = i[87];
  assign o[44803] = i[87];
  assign o[44804] = i[87];
  assign o[44805] = i[87];
  assign o[44806] = i[87];
  assign o[44807] = i[87];
  assign o[44808] = i[87];
  assign o[44809] = i[87];
  assign o[44810] = i[87];
  assign o[44811] = i[87];
  assign o[44812] = i[87];
  assign o[44813] = i[87];
  assign o[44814] = i[87];
  assign o[44815] = i[87];
  assign o[44816] = i[87];
  assign o[44817] = i[87];
  assign o[44818] = i[87];
  assign o[44819] = i[87];
  assign o[44820] = i[87];
  assign o[44821] = i[87];
  assign o[44822] = i[87];
  assign o[44823] = i[87];
  assign o[44824] = i[87];
  assign o[44825] = i[87];
  assign o[44826] = i[87];
  assign o[44827] = i[87];
  assign o[44828] = i[87];
  assign o[44829] = i[87];
  assign o[44830] = i[87];
  assign o[44831] = i[87];
  assign o[44832] = i[87];
  assign o[44833] = i[87];
  assign o[44834] = i[87];
  assign o[44835] = i[87];
  assign o[44836] = i[87];
  assign o[44837] = i[87];
  assign o[44838] = i[87];
  assign o[44839] = i[87];
  assign o[44840] = i[87];
  assign o[44841] = i[87];
  assign o[44842] = i[87];
  assign o[44843] = i[87];
  assign o[44844] = i[87];
  assign o[44845] = i[87];
  assign o[44846] = i[87];
  assign o[44847] = i[87];
  assign o[44848] = i[87];
  assign o[44849] = i[87];
  assign o[44850] = i[87];
  assign o[44851] = i[87];
  assign o[44852] = i[87];
  assign o[44853] = i[87];
  assign o[44854] = i[87];
  assign o[44855] = i[87];
  assign o[44856] = i[87];
  assign o[44857] = i[87];
  assign o[44858] = i[87];
  assign o[44859] = i[87];
  assign o[44860] = i[87];
  assign o[44861] = i[87];
  assign o[44862] = i[87];
  assign o[44863] = i[87];
  assign o[44864] = i[87];
  assign o[44865] = i[87];
  assign o[44866] = i[87];
  assign o[44867] = i[87];
  assign o[44868] = i[87];
  assign o[44869] = i[87];
  assign o[44870] = i[87];
  assign o[44871] = i[87];
  assign o[44872] = i[87];
  assign o[44873] = i[87];
  assign o[44874] = i[87];
  assign o[44875] = i[87];
  assign o[44876] = i[87];
  assign o[44877] = i[87];
  assign o[44878] = i[87];
  assign o[44879] = i[87];
  assign o[44880] = i[87];
  assign o[44881] = i[87];
  assign o[44882] = i[87];
  assign o[44883] = i[87];
  assign o[44884] = i[87];
  assign o[44885] = i[87];
  assign o[44886] = i[87];
  assign o[44887] = i[87];
  assign o[44888] = i[87];
  assign o[44889] = i[87];
  assign o[44890] = i[87];
  assign o[44891] = i[87];
  assign o[44892] = i[87];
  assign o[44893] = i[87];
  assign o[44894] = i[87];
  assign o[44895] = i[87];
  assign o[44896] = i[87];
  assign o[44897] = i[87];
  assign o[44898] = i[87];
  assign o[44899] = i[87];
  assign o[44900] = i[87];
  assign o[44901] = i[87];
  assign o[44902] = i[87];
  assign o[44903] = i[87];
  assign o[44904] = i[87];
  assign o[44905] = i[87];
  assign o[44906] = i[87];
  assign o[44907] = i[87];
  assign o[44908] = i[87];
  assign o[44909] = i[87];
  assign o[44910] = i[87];
  assign o[44911] = i[87];
  assign o[44912] = i[87];
  assign o[44913] = i[87];
  assign o[44914] = i[87];
  assign o[44915] = i[87];
  assign o[44916] = i[87];
  assign o[44917] = i[87];
  assign o[44918] = i[87];
  assign o[44919] = i[87];
  assign o[44920] = i[87];
  assign o[44921] = i[87];
  assign o[44922] = i[87];
  assign o[44923] = i[87];
  assign o[44924] = i[87];
  assign o[44925] = i[87];
  assign o[44926] = i[87];
  assign o[44927] = i[87];
  assign o[44928] = i[87];
  assign o[44929] = i[87];
  assign o[44930] = i[87];
  assign o[44931] = i[87];
  assign o[44932] = i[87];
  assign o[44933] = i[87];
  assign o[44934] = i[87];
  assign o[44935] = i[87];
  assign o[44936] = i[87];
  assign o[44937] = i[87];
  assign o[44938] = i[87];
  assign o[44939] = i[87];
  assign o[44940] = i[87];
  assign o[44941] = i[87];
  assign o[44942] = i[87];
  assign o[44943] = i[87];
  assign o[44944] = i[87];
  assign o[44945] = i[87];
  assign o[44946] = i[87];
  assign o[44947] = i[87];
  assign o[44948] = i[87];
  assign o[44949] = i[87];
  assign o[44950] = i[87];
  assign o[44951] = i[87];
  assign o[44952] = i[87];
  assign o[44953] = i[87];
  assign o[44954] = i[87];
  assign o[44955] = i[87];
  assign o[44956] = i[87];
  assign o[44957] = i[87];
  assign o[44958] = i[87];
  assign o[44959] = i[87];
  assign o[44960] = i[87];
  assign o[44961] = i[87];
  assign o[44962] = i[87];
  assign o[44963] = i[87];
  assign o[44964] = i[87];
  assign o[44965] = i[87];
  assign o[44966] = i[87];
  assign o[44967] = i[87];
  assign o[44968] = i[87];
  assign o[44969] = i[87];
  assign o[44970] = i[87];
  assign o[44971] = i[87];
  assign o[44972] = i[87];
  assign o[44973] = i[87];
  assign o[44974] = i[87];
  assign o[44975] = i[87];
  assign o[44976] = i[87];
  assign o[44977] = i[87];
  assign o[44978] = i[87];
  assign o[44979] = i[87];
  assign o[44980] = i[87];
  assign o[44981] = i[87];
  assign o[44982] = i[87];
  assign o[44983] = i[87];
  assign o[44984] = i[87];
  assign o[44985] = i[87];
  assign o[44986] = i[87];
  assign o[44987] = i[87];
  assign o[44988] = i[87];
  assign o[44989] = i[87];
  assign o[44990] = i[87];
  assign o[44991] = i[87];
  assign o[44992] = i[87];
  assign o[44993] = i[87];
  assign o[44994] = i[87];
  assign o[44995] = i[87];
  assign o[44996] = i[87];
  assign o[44997] = i[87];
  assign o[44998] = i[87];
  assign o[44999] = i[87];
  assign o[45000] = i[87];
  assign o[45001] = i[87];
  assign o[45002] = i[87];
  assign o[45003] = i[87];
  assign o[45004] = i[87];
  assign o[45005] = i[87];
  assign o[45006] = i[87];
  assign o[45007] = i[87];
  assign o[45008] = i[87];
  assign o[45009] = i[87];
  assign o[45010] = i[87];
  assign o[45011] = i[87];
  assign o[45012] = i[87];
  assign o[45013] = i[87];
  assign o[45014] = i[87];
  assign o[45015] = i[87];
  assign o[45016] = i[87];
  assign o[45017] = i[87];
  assign o[45018] = i[87];
  assign o[45019] = i[87];
  assign o[45020] = i[87];
  assign o[45021] = i[87];
  assign o[45022] = i[87];
  assign o[45023] = i[87];
  assign o[45024] = i[87];
  assign o[45025] = i[87];
  assign o[45026] = i[87];
  assign o[45027] = i[87];
  assign o[45028] = i[87];
  assign o[45029] = i[87];
  assign o[45030] = i[87];
  assign o[45031] = i[87];
  assign o[45032] = i[87];
  assign o[45033] = i[87];
  assign o[45034] = i[87];
  assign o[45035] = i[87];
  assign o[45036] = i[87];
  assign o[45037] = i[87];
  assign o[45038] = i[87];
  assign o[45039] = i[87];
  assign o[45040] = i[87];
  assign o[45041] = i[87];
  assign o[45042] = i[87];
  assign o[45043] = i[87];
  assign o[45044] = i[87];
  assign o[45045] = i[87];
  assign o[45046] = i[87];
  assign o[45047] = i[87];
  assign o[45048] = i[87];
  assign o[45049] = i[87];
  assign o[45050] = i[87];
  assign o[45051] = i[87];
  assign o[45052] = i[87];
  assign o[45053] = i[87];
  assign o[45054] = i[87];
  assign o[45055] = i[87];
  assign o[44032] = i[86];
  assign o[44033] = i[86];
  assign o[44034] = i[86];
  assign o[44035] = i[86];
  assign o[44036] = i[86];
  assign o[44037] = i[86];
  assign o[44038] = i[86];
  assign o[44039] = i[86];
  assign o[44040] = i[86];
  assign o[44041] = i[86];
  assign o[44042] = i[86];
  assign o[44043] = i[86];
  assign o[44044] = i[86];
  assign o[44045] = i[86];
  assign o[44046] = i[86];
  assign o[44047] = i[86];
  assign o[44048] = i[86];
  assign o[44049] = i[86];
  assign o[44050] = i[86];
  assign o[44051] = i[86];
  assign o[44052] = i[86];
  assign o[44053] = i[86];
  assign o[44054] = i[86];
  assign o[44055] = i[86];
  assign o[44056] = i[86];
  assign o[44057] = i[86];
  assign o[44058] = i[86];
  assign o[44059] = i[86];
  assign o[44060] = i[86];
  assign o[44061] = i[86];
  assign o[44062] = i[86];
  assign o[44063] = i[86];
  assign o[44064] = i[86];
  assign o[44065] = i[86];
  assign o[44066] = i[86];
  assign o[44067] = i[86];
  assign o[44068] = i[86];
  assign o[44069] = i[86];
  assign o[44070] = i[86];
  assign o[44071] = i[86];
  assign o[44072] = i[86];
  assign o[44073] = i[86];
  assign o[44074] = i[86];
  assign o[44075] = i[86];
  assign o[44076] = i[86];
  assign o[44077] = i[86];
  assign o[44078] = i[86];
  assign o[44079] = i[86];
  assign o[44080] = i[86];
  assign o[44081] = i[86];
  assign o[44082] = i[86];
  assign o[44083] = i[86];
  assign o[44084] = i[86];
  assign o[44085] = i[86];
  assign o[44086] = i[86];
  assign o[44087] = i[86];
  assign o[44088] = i[86];
  assign o[44089] = i[86];
  assign o[44090] = i[86];
  assign o[44091] = i[86];
  assign o[44092] = i[86];
  assign o[44093] = i[86];
  assign o[44094] = i[86];
  assign o[44095] = i[86];
  assign o[44096] = i[86];
  assign o[44097] = i[86];
  assign o[44098] = i[86];
  assign o[44099] = i[86];
  assign o[44100] = i[86];
  assign o[44101] = i[86];
  assign o[44102] = i[86];
  assign o[44103] = i[86];
  assign o[44104] = i[86];
  assign o[44105] = i[86];
  assign o[44106] = i[86];
  assign o[44107] = i[86];
  assign o[44108] = i[86];
  assign o[44109] = i[86];
  assign o[44110] = i[86];
  assign o[44111] = i[86];
  assign o[44112] = i[86];
  assign o[44113] = i[86];
  assign o[44114] = i[86];
  assign o[44115] = i[86];
  assign o[44116] = i[86];
  assign o[44117] = i[86];
  assign o[44118] = i[86];
  assign o[44119] = i[86];
  assign o[44120] = i[86];
  assign o[44121] = i[86];
  assign o[44122] = i[86];
  assign o[44123] = i[86];
  assign o[44124] = i[86];
  assign o[44125] = i[86];
  assign o[44126] = i[86];
  assign o[44127] = i[86];
  assign o[44128] = i[86];
  assign o[44129] = i[86];
  assign o[44130] = i[86];
  assign o[44131] = i[86];
  assign o[44132] = i[86];
  assign o[44133] = i[86];
  assign o[44134] = i[86];
  assign o[44135] = i[86];
  assign o[44136] = i[86];
  assign o[44137] = i[86];
  assign o[44138] = i[86];
  assign o[44139] = i[86];
  assign o[44140] = i[86];
  assign o[44141] = i[86];
  assign o[44142] = i[86];
  assign o[44143] = i[86];
  assign o[44144] = i[86];
  assign o[44145] = i[86];
  assign o[44146] = i[86];
  assign o[44147] = i[86];
  assign o[44148] = i[86];
  assign o[44149] = i[86];
  assign o[44150] = i[86];
  assign o[44151] = i[86];
  assign o[44152] = i[86];
  assign o[44153] = i[86];
  assign o[44154] = i[86];
  assign o[44155] = i[86];
  assign o[44156] = i[86];
  assign o[44157] = i[86];
  assign o[44158] = i[86];
  assign o[44159] = i[86];
  assign o[44160] = i[86];
  assign o[44161] = i[86];
  assign o[44162] = i[86];
  assign o[44163] = i[86];
  assign o[44164] = i[86];
  assign o[44165] = i[86];
  assign o[44166] = i[86];
  assign o[44167] = i[86];
  assign o[44168] = i[86];
  assign o[44169] = i[86];
  assign o[44170] = i[86];
  assign o[44171] = i[86];
  assign o[44172] = i[86];
  assign o[44173] = i[86];
  assign o[44174] = i[86];
  assign o[44175] = i[86];
  assign o[44176] = i[86];
  assign o[44177] = i[86];
  assign o[44178] = i[86];
  assign o[44179] = i[86];
  assign o[44180] = i[86];
  assign o[44181] = i[86];
  assign o[44182] = i[86];
  assign o[44183] = i[86];
  assign o[44184] = i[86];
  assign o[44185] = i[86];
  assign o[44186] = i[86];
  assign o[44187] = i[86];
  assign o[44188] = i[86];
  assign o[44189] = i[86];
  assign o[44190] = i[86];
  assign o[44191] = i[86];
  assign o[44192] = i[86];
  assign o[44193] = i[86];
  assign o[44194] = i[86];
  assign o[44195] = i[86];
  assign o[44196] = i[86];
  assign o[44197] = i[86];
  assign o[44198] = i[86];
  assign o[44199] = i[86];
  assign o[44200] = i[86];
  assign o[44201] = i[86];
  assign o[44202] = i[86];
  assign o[44203] = i[86];
  assign o[44204] = i[86];
  assign o[44205] = i[86];
  assign o[44206] = i[86];
  assign o[44207] = i[86];
  assign o[44208] = i[86];
  assign o[44209] = i[86];
  assign o[44210] = i[86];
  assign o[44211] = i[86];
  assign o[44212] = i[86];
  assign o[44213] = i[86];
  assign o[44214] = i[86];
  assign o[44215] = i[86];
  assign o[44216] = i[86];
  assign o[44217] = i[86];
  assign o[44218] = i[86];
  assign o[44219] = i[86];
  assign o[44220] = i[86];
  assign o[44221] = i[86];
  assign o[44222] = i[86];
  assign o[44223] = i[86];
  assign o[44224] = i[86];
  assign o[44225] = i[86];
  assign o[44226] = i[86];
  assign o[44227] = i[86];
  assign o[44228] = i[86];
  assign o[44229] = i[86];
  assign o[44230] = i[86];
  assign o[44231] = i[86];
  assign o[44232] = i[86];
  assign o[44233] = i[86];
  assign o[44234] = i[86];
  assign o[44235] = i[86];
  assign o[44236] = i[86];
  assign o[44237] = i[86];
  assign o[44238] = i[86];
  assign o[44239] = i[86];
  assign o[44240] = i[86];
  assign o[44241] = i[86];
  assign o[44242] = i[86];
  assign o[44243] = i[86];
  assign o[44244] = i[86];
  assign o[44245] = i[86];
  assign o[44246] = i[86];
  assign o[44247] = i[86];
  assign o[44248] = i[86];
  assign o[44249] = i[86];
  assign o[44250] = i[86];
  assign o[44251] = i[86];
  assign o[44252] = i[86];
  assign o[44253] = i[86];
  assign o[44254] = i[86];
  assign o[44255] = i[86];
  assign o[44256] = i[86];
  assign o[44257] = i[86];
  assign o[44258] = i[86];
  assign o[44259] = i[86];
  assign o[44260] = i[86];
  assign o[44261] = i[86];
  assign o[44262] = i[86];
  assign o[44263] = i[86];
  assign o[44264] = i[86];
  assign o[44265] = i[86];
  assign o[44266] = i[86];
  assign o[44267] = i[86];
  assign o[44268] = i[86];
  assign o[44269] = i[86];
  assign o[44270] = i[86];
  assign o[44271] = i[86];
  assign o[44272] = i[86];
  assign o[44273] = i[86];
  assign o[44274] = i[86];
  assign o[44275] = i[86];
  assign o[44276] = i[86];
  assign o[44277] = i[86];
  assign o[44278] = i[86];
  assign o[44279] = i[86];
  assign o[44280] = i[86];
  assign o[44281] = i[86];
  assign o[44282] = i[86];
  assign o[44283] = i[86];
  assign o[44284] = i[86];
  assign o[44285] = i[86];
  assign o[44286] = i[86];
  assign o[44287] = i[86];
  assign o[44288] = i[86];
  assign o[44289] = i[86];
  assign o[44290] = i[86];
  assign o[44291] = i[86];
  assign o[44292] = i[86];
  assign o[44293] = i[86];
  assign o[44294] = i[86];
  assign o[44295] = i[86];
  assign o[44296] = i[86];
  assign o[44297] = i[86];
  assign o[44298] = i[86];
  assign o[44299] = i[86];
  assign o[44300] = i[86];
  assign o[44301] = i[86];
  assign o[44302] = i[86];
  assign o[44303] = i[86];
  assign o[44304] = i[86];
  assign o[44305] = i[86];
  assign o[44306] = i[86];
  assign o[44307] = i[86];
  assign o[44308] = i[86];
  assign o[44309] = i[86];
  assign o[44310] = i[86];
  assign o[44311] = i[86];
  assign o[44312] = i[86];
  assign o[44313] = i[86];
  assign o[44314] = i[86];
  assign o[44315] = i[86];
  assign o[44316] = i[86];
  assign o[44317] = i[86];
  assign o[44318] = i[86];
  assign o[44319] = i[86];
  assign o[44320] = i[86];
  assign o[44321] = i[86];
  assign o[44322] = i[86];
  assign o[44323] = i[86];
  assign o[44324] = i[86];
  assign o[44325] = i[86];
  assign o[44326] = i[86];
  assign o[44327] = i[86];
  assign o[44328] = i[86];
  assign o[44329] = i[86];
  assign o[44330] = i[86];
  assign o[44331] = i[86];
  assign o[44332] = i[86];
  assign o[44333] = i[86];
  assign o[44334] = i[86];
  assign o[44335] = i[86];
  assign o[44336] = i[86];
  assign o[44337] = i[86];
  assign o[44338] = i[86];
  assign o[44339] = i[86];
  assign o[44340] = i[86];
  assign o[44341] = i[86];
  assign o[44342] = i[86];
  assign o[44343] = i[86];
  assign o[44344] = i[86];
  assign o[44345] = i[86];
  assign o[44346] = i[86];
  assign o[44347] = i[86];
  assign o[44348] = i[86];
  assign o[44349] = i[86];
  assign o[44350] = i[86];
  assign o[44351] = i[86];
  assign o[44352] = i[86];
  assign o[44353] = i[86];
  assign o[44354] = i[86];
  assign o[44355] = i[86];
  assign o[44356] = i[86];
  assign o[44357] = i[86];
  assign o[44358] = i[86];
  assign o[44359] = i[86];
  assign o[44360] = i[86];
  assign o[44361] = i[86];
  assign o[44362] = i[86];
  assign o[44363] = i[86];
  assign o[44364] = i[86];
  assign o[44365] = i[86];
  assign o[44366] = i[86];
  assign o[44367] = i[86];
  assign o[44368] = i[86];
  assign o[44369] = i[86];
  assign o[44370] = i[86];
  assign o[44371] = i[86];
  assign o[44372] = i[86];
  assign o[44373] = i[86];
  assign o[44374] = i[86];
  assign o[44375] = i[86];
  assign o[44376] = i[86];
  assign o[44377] = i[86];
  assign o[44378] = i[86];
  assign o[44379] = i[86];
  assign o[44380] = i[86];
  assign o[44381] = i[86];
  assign o[44382] = i[86];
  assign o[44383] = i[86];
  assign o[44384] = i[86];
  assign o[44385] = i[86];
  assign o[44386] = i[86];
  assign o[44387] = i[86];
  assign o[44388] = i[86];
  assign o[44389] = i[86];
  assign o[44390] = i[86];
  assign o[44391] = i[86];
  assign o[44392] = i[86];
  assign o[44393] = i[86];
  assign o[44394] = i[86];
  assign o[44395] = i[86];
  assign o[44396] = i[86];
  assign o[44397] = i[86];
  assign o[44398] = i[86];
  assign o[44399] = i[86];
  assign o[44400] = i[86];
  assign o[44401] = i[86];
  assign o[44402] = i[86];
  assign o[44403] = i[86];
  assign o[44404] = i[86];
  assign o[44405] = i[86];
  assign o[44406] = i[86];
  assign o[44407] = i[86];
  assign o[44408] = i[86];
  assign o[44409] = i[86];
  assign o[44410] = i[86];
  assign o[44411] = i[86];
  assign o[44412] = i[86];
  assign o[44413] = i[86];
  assign o[44414] = i[86];
  assign o[44415] = i[86];
  assign o[44416] = i[86];
  assign o[44417] = i[86];
  assign o[44418] = i[86];
  assign o[44419] = i[86];
  assign o[44420] = i[86];
  assign o[44421] = i[86];
  assign o[44422] = i[86];
  assign o[44423] = i[86];
  assign o[44424] = i[86];
  assign o[44425] = i[86];
  assign o[44426] = i[86];
  assign o[44427] = i[86];
  assign o[44428] = i[86];
  assign o[44429] = i[86];
  assign o[44430] = i[86];
  assign o[44431] = i[86];
  assign o[44432] = i[86];
  assign o[44433] = i[86];
  assign o[44434] = i[86];
  assign o[44435] = i[86];
  assign o[44436] = i[86];
  assign o[44437] = i[86];
  assign o[44438] = i[86];
  assign o[44439] = i[86];
  assign o[44440] = i[86];
  assign o[44441] = i[86];
  assign o[44442] = i[86];
  assign o[44443] = i[86];
  assign o[44444] = i[86];
  assign o[44445] = i[86];
  assign o[44446] = i[86];
  assign o[44447] = i[86];
  assign o[44448] = i[86];
  assign o[44449] = i[86];
  assign o[44450] = i[86];
  assign o[44451] = i[86];
  assign o[44452] = i[86];
  assign o[44453] = i[86];
  assign o[44454] = i[86];
  assign o[44455] = i[86];
  assign o[44456] = i[86];
  assign o[44457] = i[86];
  assign o[44458] = i[86];
  assign o[44459] = i[86];
  assign o[44460] = i[86];
  assign o[44461] = i[86];
  assign o[44462] = i[86];
  assign o[44463] = i[86];
  assign o[44464] = i[86];
  assign o[44465] = i[86];
  assign o[44466] = i[86];
  assign o[44467] = i[86];
  assign o[44468] = i[86];
  assign o[44469] = i[86];
  assign o[44470] = i[86];
  assign o[44471] = i[86];
  assign o[44472] = i[86];
  assign o[44473] = i[86];
  assign o[44474] = i[86];
  assign o[44475] = i[86];
  assign o[44476] = i[86];
  assign o[44477] = i[86];
  assign o[44478] = i[86];
  assign o[44479] = i[86];
  assign o[44480] = i[86];
  assign o[44481] = i[86];
  assign o[44482] = i[86];
  assign o[44483] = i[86];
  assign o[44484] = i[86];
  assign o[44485] = i[86];
  assign o[44486] = i[86];
  assign o[44487] = i[86];
  assign o[44488] = i[86];
  assign o[44489] = i[86];
  assign o[44490] = i[86];
  assign o[44491] = i[86];
  assign o[44492] = i[86];
  assign o[44493] = i[86];
  assign o[44494] = i[86];
  assign o[44495] = i[86];
  assign o[44496] = i[86];
  assign o[44497] = i[86];
  assign o[44498] = i[86];
  assign o[44499] = i[86];
  assign o[44500] = i[86];
  assign o[44501] = i[86];
  assign o[44502] = i[86];
  assign o[44503] = i[86];
  assign o[44504] = i[86];
  assign o[44505] = i[86];
  assign o[44506] = i[86];
  assign o[44507] = i[86];
  assign o[44508] = i[86];
  assign o[44509] = i[86];
  assign o[44510] = i[86];
  assign o[44511] = i[86];
  assign o[44512] = i[86];
  assign o[44513] = i[86];
  assign o[44514] = i[86];
  assign o[44515] = i[86];
  assign o[44516] = i[86];
  assign o[44517] = i[86];
  assign o[44518] = i[86];
  assign o[44519] = i[86];
  assign o[44520] = i[86];
  assign o[44521] = i[86];
  assign o[44522] = i[86];
  assign o[44523] = i[86];
  assign o[44524] = i[86];
  assign o[44525] = i[86];
  assign o[44526] = i[86];
  assign o[44527] = i[86];
  assign o[44528] = i[86];
  assign o[44529] = i[86];
  assign o[44530] = i[86];
  assign o[44531] = i[86];
  assign o[44532] = i[86];
  assign o[44533] = i[86];
  assign o[44534] = i[86];
  assign o[44535] = i[86];
  assign o[44536] = i[86];
  assign o[44537] = i[86];
  assign o[44538] = i[86];
  assign o[44539] = i[86];
  assign o[44540] = i[86];
  assign o[44541] = i[86];
  assign o[44542] = i[86];
  assign o[44543] = i[86];
  assign o[43520] = i[85];
  assign o[43521] = i[85];
  assign o[43522] = i[85];
  assign o[43523] = i[85];
  assign o[43524] = i[85];
  assign o[43525] = i[85];
  assign o[43526] = i[85];
  assign o[43527] = i[85];
  assign o[43528] = i[85];
  assign o[43529] = i[85];
  assign o[43530] = i[85];
  assign o[43531] = i[85];
  assign o[43532] = i[85];
  assign o[43533] = i[85];
  assign o[43534] = i[85];
  assign o[43535] = i[85];
  assign o[43536] = i[85];
  assign o[43537] = i[85];
  assign o[43538] = i[85];
  assign o[43539] = i[85];
  assign o[43540] = i[85];
  assign o[43541] = i[85];
  assign o[43542] = i[85];
  assign o[43543] = i[85];
  assign o[43544] = i[85];
  assign o[43545] = i[85];
  assign o[43546] = i[85];
  assign o[43547] = i[85];
  assign o[43548] = i[85];
  assign o[43549] = i[85];
  assign o[43550] = i[85];
  assign o[43551] = i[85];
  assign o[43552] = i[85];
  assign o[43553] = i[85];
  assign o[43554] = i[85];
  assign o[43555] = i[85];
  assign o[43556] = i[85];
  assign o[43557] = i[85];
  assign o[43558] = i[85];
  assign o[43559] = i[85];
  assign o[43560] = i[85];
  assign o[43561] = i[85];
  assign o[43562] = i[85];
  assign o[43563] = i[85];
  assign o[43564] = i[85];
  assign o[43565] = i[85];
  assign o[43566] = i[85];
  assign o[43567] = i[85];
  assign o[43568] = i[85];
  assign o[43569] = i[85];
  assign o[43570] = i[85];
  assign o[43571] = i[85];
  assign o[43572] = i[85];
  assign o[43573] = i[85];
  assign o[43574] = i[85];
  assign o[43575] = i[85];
  assign o[43576] = i[85];
  assign o[43577] = i[85];
  assign o[43578] = i[85];
  assign o[43579] = i[85];
  assign o[43580] = i[85];
  assign o[43581] = i[85];
  assign o[43582] = i[85];
  assign o[43583] = i[85];
  assign o[43584] = i[85];
  assign o[43585] = i[85];
  assign o[43586] = i[85];
  assign o[43587] = i[85];
  assign o[43588] = i[85];
  assign o[43589] = i[85];
  assign o[43590] = i[85];
  assign o[43591] = i[85];
  assign o[43592] = i[85];
  assign o[43593] = i[85];
  assign o[43594] = i[85];
  assign o[43595] = i[85];
  assign o[43596] = i[85];
  assign o[43597] = i[85];
  assign o[43598] = i[85];
  assign o[43599] = i[85];
  assign o[43600] = i[85];
  assign o[43601] = i[85];
  assign o[43602] = i[85];
  assign o[43603] = i[85];
  assign o[43604] = i[85];
  assign o[43605] = i[85];
  assign o[43606] = i[85];
  assign o[43607] = i[85];
  assign o[43608] = i[85];
  assign o[43609] = i[85];
  assign o[43610] = i[85];
  assign o[43611] = i[85];
  assign o[43612] = i[85];
  assign o[43613] = i[85];
  assign o[43614] = i[85];
  assign o[43615] = i[85];
  assign o[43616] = i[85];
  assign o[43617] = i[85];
  assign o[43618] = i[85];
  assign o[43619] = i[85];
  assign o[43620] = i[85];
  assign o[43621] = i[85];
  assign o[43622] = i[85];
  assign o[43623] = i[85];
  assign o[43624] = i[85];
  assign o[43625] = i[85];
  assign o[43626] = i[85];
  assign o[43627] = i[85];
  assign o[43628] = i[85];
  assign o[43629] = i[85];
  assign o[43630] = i[85];
  assign o[43631] = i[85];
  assign o[43632] = i[85];
  assign o[43633] = i[85];
  assign o[43634] = i[85];
  assign o[43635] = i[85];
  assign o[43636] = i[85];
  assign o[43637] = i[85];
  assign o[43638] = i[85];
  assign o[43639] = i[85];
  assign o[43640] = i[85];
  assign o[43641] = i[85];
  assign o[43642] = i[85];
  assign o[43643] = i[85];
  assign o[43644] = i[85];
  assign o[43645] = i[85];
  assign o[43646] = i[85];
  assign o[43647] = i[85];
  assign o[43648] = i[85];
  assign o[43649] = i[85];
  assign o[43650] = i[85];
  assign o[43651] = i[85];
  assign o[43652] = i[85];
  assign o[43653] = i[85];
  assign o[43654] = i[85];
  assign o[43655] = i[85];
  assign o[43656] = i[85];
  assign o[43657] = i[85];
  assign o[43658] = i[85];
  assign o[43659] = i[85];
  assign o[43660] = i[85];
  assign o[43661] = i[85];
  assign o[43662] = i[85];
  assign o[43663] = i[85];
  assign o[43664] = i[85];
  assign o[43665] = i[85];
  assign o[43666] = i[85];
  assign o[43667] = i[85];
  assign o[43668] = i[85];
  assign o[43669] = i[85];
  assign o[43670] = i[85];
  assign o[43671] = i[85];
  assign o[43672] = i[85];
  assign o[43673] = i[85];
  assign o[43674] = i[85];
  assign o[43675] = i[85];
  assign o[43676] = i[85];
  assign o[43677] = i[85];
  assign o[43678] = i[85];
  assign o[43679] = i[85];
  assign o[43680] = i[85];
  assign o[43681] = i[85];
  assign o[43682] = i[85];
  assign o[43683] = i[85];
  assign o[43684] = i[85];
  assign o[43685] = i[85];
  assign o[43686] = i[85];
  assign o[43687] = i[85];
  assign o[43688] = i[85];
  assign o[43689] = i[85];
  assign o[43690] = i[85];
  assign o[43691] = i[85];
  assign o[43692] = i[85];
  assign o[43693] = i[85];
  assign o[43694] = i[85];
  assign o[43695] = i[85];
  assign o[43696] = i[85];
  assign o[43697] = i[85];
  assign o[43698] = i[85];
  assign o[43699] = i[85];
  assign o[43700] = i[85];
  assign o[43701] = i[85];
  assign o[43702] = i[85];
  assign o[43703] = i[85];
  assign o[43704] = i[85];
  assign o[43705] = i[85];
  assign o[43706] = i[85];
  assign o[43707] = i[85];
  assign o[43708] = i[85];
  assign o[43709] = i[85];
  assign o[43710] = i[85];
  assign o[43711] = i[85];
  assign o[43712] = i[85];
  assign o[43713] = i[85];
  assign o[43714] = i[85];
  assign o[43715] = i[85];
  assign o[43716] = i[85];
  assign o[43717] = i[85];
  assign o[43718] = i[85];
  assign o[43719] = i[85];
  assign o[43720] = i[85];
  assign o[43721] = i[85];
  assign o[43722] = i[85];
  assign o[43723] = i[85];
  assign o[43724] = i[85];
  assign o[43725] = i[85];
  assign o[43726] = i[85];
  assign o[43727] = i[85];
  assign o[43728] = i[85];
  assign o[43729] = i[85];
  assign o[43730] = i[85];
  assign o[43731] = i[85];
  assign o[43732] = i[85];
  assign o[43733] = i[85];
  assign o[43734] = i[85];
  assign o[43735] = i[85];
  assign o[43736] = i[85];
  assign o[43737] = i[85];
  assign o[43738] = i[85];
  assign o[43739] = i[85];
  assign o[43740] = i[85];
  assign o[43741] = i[85];
  assign o[43742] = i[85];
  assign o[43743] = i[85];
  assign o[43744] = i[85];
  assign o[43745] = i[85];
  assign o[43746] = i[85];
  assign o[43747] = i[85];
  assign o[43748] = i[85];
  assign o[43749] = i[85];
  assign o[43750] = i[85];
  assign o[43751] = i[85];
  assign o[43752] = i[85];
  assign o[43753] = i[85];
  assign o[43754] = i[85];
  assign o[43755] = i[85];
  assign o[43756] = i[85];
  assign o[43757] = i[85];
  assign o[43758] = i[85];
  assign o[43759] = i[85];
  assign o[43760] = i[85];
  assign o[43761] = i[85];
  assign o[43762] = i[85];
  assign o[43763] = i[85];
  assign o[43764] = i[85];
  assign o[43765] = i[85];
  assign o[43766] = i[85];
  assign o[43767] = i[85];
  assign o[43768] = i[85];
  assign o[43769] = i[85];
  assign o[43770] = i[85];
  assign o[43771] = i[85];
  assign o[43772] = i[85];
  assign o[43773] = i[85];
  assign o[43774] = i[85];
  assign o[43775] = i[85];
  assign o[43776] = i[85];
  assign o[43777] = i[85];
  assign o[43778] = i[85];
  assign o[43779] = i[85];
  assign o[43780] = i[85];
  assign o[43781] = i[85];
  assign o[43782] = i[85];
  assign o[43783] = i[85];
  assign o[43784] = i[85];
  assign o[43785] = i[85];
  assign o[43786] = i[85];
  assign o[43787] = i[85];
  assign o[43788] = i[85];
  assign o[43789] = i[85];
  assign o[43790] = i[85];
  assign o[43791] = i[85];
  assign o[43792] = i[85];
  assign o[43793] = i[85];
  assign o[43794] = i[85];
  assign o[43795] = i[85];
  assign o[43796] = i[85];
  assign o[43797] = i[85];
  assign o[43798] = i[85];
  assign o[43799] = i[85];
  assign o[43800] = i[85];
  assign o[43801] = i[85];
  assign o[43802] = i[85];
  assign o[43803] = i[85];
  assign o[43804] = i[85];
  assign o[43805] = i[85];
  assign o[43806] = i[85];
  assign o[43807] = i[85];
  assign o[43808] = i[85];
  assign o[43809] = i[85];
  assign o[43810] = i[85];
  assign o[43811] = i[85];
  assign o[43812] = i[85];
  assign o[43813] = i[85];
  assign o[43814] = i[85];
  assign o[43815] = i[85];
  assign o[43816] = i[85];
  assign o[43817] = i[85];
  assign o[43818] = i[85];
  assign o[43819] = i[85];
  assign o[43820] = i[85];
  assign o[43821] = i[85];
  assign o[43822] = i[85];
  assign o[43823] = i[85];
  assign o[43824] = i[85];
  assign o[43825] = i[85];
  assign o[43826] = i[85];
  assign o[43827] = i[85];
  assign o[43828] = i[85];
  assign o[43829] = i[85];
  assign o[43830] = i[85];
  assign o[43831] = i[85];
  assign o[43832] = i[85];
  assign o[43833] = i[85];
  assign o[43834] = i[85];
  assign o[43835] = i[85];
  assign o[43836] = i[85];
  assign o[43837] = i[85];
  assign o[43838] = i[85];
  assign o[43839] = i[85];
  assign o[43840] = i[85];
  assign o[43841] = i[85];
  assign o[43842] = i[85];
  assign o[43843] = i[85];
  assign o[43844] = i[85];
  assign o[43845] = i[85];
  assign o[43846] = i[85];
  assign o[43847] = i[85];
  assign o[43848] = i[85];
  assign o[43849] = i[85];
  assign o[43850] = i[85];
  assign o[43851] = i[85];
  assign o[43852] = i[85];
  assign o[43853] = i[85];
  assign o[43854] = i[85];
  assign o[43855] = i[85];
  assign o[43856] = i[85];
  assign o[43857] = i[85];
  assign o[43858] = i[85];
  assign o[43859] = i[85];
  assign o[43860] = i[85];
  assign o[43861] = i[85];
  assign o[43862] = i[85];
  assign o[43863] = i[85];
  assign o[43864] = i[85];
  assign o[43865] = i[85];
  assign o[43866] = i[85];
  assign o[43867] = i[85];
  assign o[43868] = i[85];
  assign o[43869] = i[85];
  assign o[43870] = i[85];
  assign o[43871] = i[85];
  assign o[43872] = i[85];
  assign o[43873] = i[85];
  assign o[43874] = i[85];
  assign o[43875] = i[85];
  assign o[43876] = i[85];
  assign o[43877] = i[85];
  assign o[43878] = i[85];
  assign o[43879] = i[85];
  assign o[43880] = i[85];
  assign o[43881] = i[85];
  assign o[43882] = i[85];
  assign o[43883] = i[85];
  assign o[43884] = i[85];
  assign o[43885] = i[85];
  assign o[43886] = i[85];
  assign o[43887] = i[85];
  assign o[43888] = i[85];
  assign o[43889] = i[85];
  assign o[43890] = i[85];
  assign o[43891] = i[85];
  assign o[43892] = i[85];
  assign o[43893] = i[85];
  assign o[43894] = i[85];
  assign o[43895] = i[85];
  assign o[43896] = i[85];
  assign o[43897] = i[85];
  assign o[43898] = i[85];
  assign o[43899] = i[85];
  assign o[43900] = i[85];
  assign o[43901] = i[85];
  assign o[43902] = i[85];
  assign o[43903] = i[85];
  assign o[43904] = i[85];
  assign o[43905] = i[85];
  assign o[43906] = i[85];
  assign o[43907] = i[85];
  assign o[43908] = i[85];
  assign o[43909] = i[85];
  assign o[43910] = i[85];
  assign o[43911] = i[85];
  assign o[43912] = i[85];
  assign o[43913] = i[85];
  assign o[43914] = i[85];
  assign o[43915] = i[85];
  assign o[43916] = i[85];
  assign o[43917] = i[85];
  assign o[43918] = i[85];
  assign o[43919] = i[85];
  assign o[43920] = i[85];
  assign o[43921] = i[85];
  assign o[43922] = i[85];
  assign o[43923] = i[85];
  assign o[43924] = i[85];
  assign o[43925] = i[85];
  assign o[43926] = i[85];
  assign o[43927] = i[85];
  assign o[43928] = i[85];
  assign o[43929] = i[85];
  assign o[43930] = i[85];
  assign o[43931] = i[85];
  assign o[43932] = i[85];
  assign o[43933] = i[85];
  assign o[43934] = i[85];
  assign o[43935] = i[85];
  assign o[43936] = i[85];
  assign o[43937] = i[85];
  assign o[43938] = i[85];
  assign o[43939] = i[85];
  assign o[43940] = i[85];
  assign o[43941] = i[85];
  assign o[43942] = i[85];
  assign o[43943] = i[85];
  assign o[43944] = i[85];
  assign o[43945] = i[85];
  assign o[43946] = i[85];
  assign o[43947] = i[85];
  assign o[43948] = i[85];
  assign o[43949] = i[85];
  assign o[43950] = i[85];
  assign o[43951] = i[85];
  assign o[43952] = i[85];
  assign o[43953] = i[85];
  assign o[43954] = i[85];
  assign o[43955] = i[85];
  assign o[43956] = i[85];
  assign o[43957] = i[85];
  assign o[43958] = i[85];
  assign o[43959] = i[85];
  assign o[43960] = i[85];
  assign o[43961] = i[85];
  assign o[43962] = i[85];
  assign o[43963] = i[85];
  assign o[43964] = i[85];
  assign o[43965] = i[85];
  assign o[43966] = i[85];
  assign o[43967] = i[85];
  assign o[43968] = i[85];
  assign o[43969] = i[85];
  assign o[43970] = i[85];
  assign o[43971] = i[85];
  assign o[43972] = i[85];
  assign o[43973] = i[85];
  assign o[43974] = i[85];
  assign o[43975] = i[85];
  assign o[43976] = i[85];
  assign o[43977] = i[85];
  assign o[43978] = i[85];
  assign o[43979] = i[85];
  assign o[43980] = i[85];
  assign o[43981] = i[85];
  assign o[43982] = i[85];
  assign o[43983] = i[85];
  assign o[43984] = i[85];
  assign o[43985] = i[85];
  assign o[43986] = i[85];
  assign o[43987] = i[85];
  assign o[43988] = i[85];
  assign o[43989] = i[85];
  assign o[43990] = i[85];
  assign o[43991] = i[85];
  assign o[43992] = i[85];
  assign o[43993] = i[85];
  assign o[43994] = i[85];
  assign o[43995] = i[85];
  assign o[43996] = i[85];
  assign o[43997] = i[85];
  assign o[43998] = i[85];
  assign o[43999] = i[85];
  assign o[44000] = i[85];
  assign o[44001] = i[85];
  assign o[44002] = i[85];
  assign o[44003] = i[85];
  assign o[44004] = i[85];
  assign o[44005] = i[85];
  assign o[44006] = i[85];
  assign o[44007] = i[85];
  assign o[44008] = i[85];
  assign o[44009] = i[85];
  assign o[44010] = i[85];
  assign o[44011] = i[85];
  assign o[44012] = i[85];
  assign o[44013] = i[85];
  assign o[44014] = i[85];
  assign o[44015] = i[85];
  assign o[44016] = i[85];
  assign o[44017] = i[85];
  assign o[44018] = i[85];
  assign o[44019] = i[85];
  assign o[44020] = i[85];
  assign o[44021] = i[85];
  assign o[44022] = i[85];
  assign o[44023] = i[85];
  assign o[44024] = i[85];
  assign o[44025] = i[85];
  assign o[44026] = i[85];
  assign o[44027] = i[85];
  assign o[44028] = i[85];
  assign o[44029] = i[85];
  assign o[44030] = i[85];
  assign o[44031] = i[85];
  assign o[43008] = i[84];
  assign o[43009] = i[84];
  assign o[43010] = i[84];
  assign o[43011] = i[84];
  assign o[43012] = i[84];
  assign o[43013] = i[84];
  assign o[43014] = i[84];
  assign o[43015] = i[84];
  assign o[43016] = i[84];
  assign o[43017] = i[84];
  assign o[43018] = i[84];
  assign o[43019] = i[84];
  assign o[43020] = i[84];
  assign o[43021] = i[84];
  assign o[43022] = i[84];
  assign o[43023] = i[84];
  assign o[43024] = i[84];
  assign o[43025] = i[84];
  assign o[43026] = i[84];
  assign o[43027] = i[84];
  assign o[43028] = i[84];
  assign o[43029] = i[84];
  assign o[43030] = i[84];
  assign o[43031] = i[84];
  assign o[43032] = i[84];
  assign o[43033] = i[84];
  assign o[43034] = i[84];
  assign o[43035] = i[84];
  assign o[43036] = i[84];
  assign o[43037] = i[84];
  assign o[43038] = i[84];
  assign o[43039] = i[84];
  assign o[43040] = i[84];
  assign o[43041] = i[84];
  assign o[43042] = i[84];
  assign o[43043] = i[84];
  assign o[43044] = i[84];
  assign o[43045] = i[84];
  assign o[43046] = i[84];
  assign o[43047] = i[84];
  assign o[43048] = i[84];
  assign o[43049] = i[84];
  assign o[43050] = i[84];
  assign o[43051] = i[84];
  assign o[43052] = i[84];
  assign o[43053] = i[84];
  assign o[43054] = i[84];
  assign o[43055] = i[84];
  assign o[43056] = i[84];
  assign o[43057] = i[84];
  assign o[43058] = i[84];
  assign o[43059] = i[84];
  assign o[43060] = i[84];
  assign o[43061] = i[84];
  assign o[43062] = i[84];
  assign o[43063] = i[84];
  assign o[43064] = i[84];
  assign o[43065] = i[84];
  assign o[43066] = i[84];
  assign o[43067] = i[84];
  assign o[43068] = i[84];
  assign o[43069] = i[84];
  assign o[43070] = i[84];
  assign o[43071] = i[84];
  assign o[43072] = i[84];
  assign o[43073] = i[84];
  assign o[43074] = i[84];
  assign o[43075] = i[84];
  assign o[43076] = i[84];
  assign o[43077] = i[84];
  assign o[43078] = i[84];
  assign o[43079] = i[84];
  assign o[43080] = i[84];
  assign o[43081] = i[84];
  assign o[43082] = i[84];
  assign o[43083] = i[84];
  assign o[43084] = i[84];
  assign o[43085] = i[84];
  assign o[43086] = i[84];
  assign o[43087] = i[84];
  assign o[43088] = i[84];
  assign o[43089] = i[84];
  assign o[43090] = i[84];
  assign o[43091] = i[84];
  assign o[43092] = i[84];
  assign o[43093] = i[84];
  assign o[43094] = i[84];
  assign o[43095] = i[84];
  assign o[43096] = i[84];
  assign o[43097] = i[84];
  assign o[43098] = i[84];
  assign o[43099] = i[84];
  assign o[43100] = i[84];
  assign o[43101] = i[84];
  assign o[43102] = i[84];
  assign o[43103] = i[84];
  assign o[43104] = i[84];
  assign o[43105] = i[84];
  assign o[43106] = i[84];
  assign o[43107] = i[84];
  assign o[43108] = i[84];
  assign o[43109] = i[84];
  assign o[43110] = i[84];
  assign o[43111] = i[84];
  assign o[43112] = i[84];
  assign o[43113] = i[84];
  assign o[43114] = i[84];
  assign o[43115] = i[84];
  assign o[43116] = i[84];
  assign o[43117] = i[84];
  assign o[43118] = i[84];
  assign o[43119] = i[84];
  assign o[43120] = i[84];
  assign o[43121] = i[84];
  assign o[43122] = i[84];
  assign o[43123] = i[84];
  assign o[43124] = i[84];
  assign o[43125] = i[84];
  assign o[43126] = i[84];
  assign o[43127] = i[84];
  assign o[43128] = i[84];
  assign o[43129] = i[84];
  assign o[43130] = i[84];
  assign o[43131] = i[84];
  assign o[43132] = i[84];
  assign o[43133] = i[84];
  assign o[43134] = i[84];
  assign o[43135] = i[84];
  assign o[43136] = i[84];
  assign o[43137] = i[84];
  assign o[43138] = i[84];
  assign o[43139] = i[84];
  assign o[43140] = i[84];
  assign o[43141] = i[84];
  assign o[43142] = i[84];
  assign o[43143] = i[84];
  assign o[43144] = i[84];
  assign o[43145] = i[84];
  assign o[43146] = i[84];
  assign o[43147] = i[84];
  assign o[43148] = i[84];
  assign o[43149] = i[84];
  assign o[43150] = i[84];
  assign o[43151] = i[84];
  assign o[43152] = i[84];
  assign o[43153] = i[84];
  assign o[43154] = i[84];
  assign o[43155] = i[84];
  assign o[43156] = i[84];
  assign o[43157] = i[84];
  assign o[43158] = i[84];
  assign o[43159] = i[84];
  assign o[43160] = i[84];
  assign o[43161] = i[84];
  assign o[43162] = i[84];
  assign o[43163] = i[84];
  assign o[43164] = i[84];
  assign o[43165] = i[84];
  assign o[43166] = i[84];
  assign o[43167] = i[84];
  assign o[43168] = i[84];
  assign o[43169] = i[84];
  assign o[43170] = i[84];
  assign o[43171] = i[84];
  assign o[43172] = i[84];
  assign o[43173] = i[84];
  assign o[43174] = i[84];
  assign o[43175] = i[84];
  assign o[43176] = i[84];
  assign o[43177] = i[84];
  assign o[43178] = i[84];
  assign o[43179] = i[84];
  assign o[43180] = i[84];
  assign o[43181] = i[84];
  assign o[43182] = i[84];
  assign o[43183] = i[84];
  assign o[43184] = i[84];
  assign o[43185] = i[84];
  assign o[43186] = i[84];
  assign o[43187] = i[84];
  assign o[43188] = i[84];
  assign o[43189] = i[84];
  assign o[43190] = i[84];
  assign o[43191] = i[84];
  assign o[43192] = i[84];
  assign o[43193] = i[84];
  assign o[43194] = i[84];
  assign o[43195] = i[84];
  assign o[43196] = i[84];
  assign o[43197] = i[84];
  assign o[43198] = i[84];
  assign o[43199] = i[84];
  assign o[43200] = i[84];
  assign o[43201] = i[84];
  assign o[43202] = i[84];
  assign o[43203] = i[84];
  assign o[43204] = i[84];
  assign o[43205] = i[84];
  assign o[43206] = i[84];
  assign o[43207] = i[84];
  assign o[43208] = i[84];
  assign o[43209] = i[84];
  assign o[43210] = i[84];
  assign o[43211] = i[84];
  assign o[43212] = i[84];
  assign o[43213] = i[84];
  assign o[43214] = i[84];
  assign o[43215] = i[84];
  assign o[43216] = i[84];
  assign o[43217] = i[84];
  assign o[43218] = i[84];
  assign o[43219] = i[84];
  assign o[43220] = i[84];
  assign o[43221] = i[84];
  assign o[43222] = i[84];
  assign o[43223] = i[84];
  assign o[43224] = i[84];
  assign o[43225] = i[84];
  assign o[43226] = i[84];
  assign o[43227] = i[84];
  assign o[43228] = i[84];
  assign o[43229] = i[84];
  assign o[43230] = i[84];
  assign o[43231] = i[84];
  assign o[43232] = i[84];
  assign o[43233] = i[84];
  assign o[43234] = i[84];
  assign o[43235] = i[84];
  assign o[43236] = i[84];
  assign o[43237] = i[84];
  assign o[43238] = i[84];
  assign o[43239] = i[84];
  assign o[43240] = i[84];
  assign o[43241] = i[84];
  assign o[43242] = i[84];
  assign o[43243] = i[84];
  assign o[43244] = i[84];
  assign o[43245] = i[84];
  assign o[43246] = i[84];
  assign o[43247] = i[84];
  assign o[43248] = i[84];
  assign o[43249] = i[84];
  assign o[43250] = i[84];
  assign o[43251] = i[84];
  assign o[43252] = i[84];
  assign o[43253] = i[84];
  assign o[43254] = i[84];
  assign o[43255] = i[84];
  assign o[43256] = i[84];
  assign o[43257] = i[84];
  assign o[43258] = i[84];
  assign o[43259] = i[84];
  assign o[43260] = i[84];
  assign o[43261] = i[84];
  assign o[43262] = i[84];
  assign o[43263] = i[84];
  assign o[43264] = i[84];
  assign o[43265] = i[84];
  assign o[43266] = i[84];
  assign o[43267] = i[84];
  assign o[43268] = i[84];
  assign o[43269] = i[84];
  assign o[43270] = i[84];
  assign o[43271] = i[84];
  assign o[43272] = i[84];
  assign o[43273] = i[84];
  assign o[43274] = i[84];
  assign o[43275] = i[84];
  assign o[43276] = i[84];
  assign o[43277] = i[84];
  assign o[43278] = i[84];
  assign o[43279] = i[84];
  assign o[43280] = i[84];
  assign o[43281] = i[84];
  assign o[43282] = i[84];
  assign o[43283] = i[84];
  assign o[43284] = i[84];
  assign o[43285] = i[84];
  assign o[43286] = i[84];
  assign o[43287] = i[84];
  assign o[43288] = i[84];
  assign o[43289] = i[84];
  assign o[43290] = i[84];
  assign o[43291] = i[84];
  assign o[43292] = i[84];
  assign o[43293] = i[84];
  assign o[43294] = i[84];
  assign o[43295] = i[84];
  assign o[43296] = i[84];
  assign o[43297] = i[84];
  assign o[43298] = i[84];
  assign o[43299] = i[84];
  assign o[43300] = i[84];
  assign o[43301] = i[84];
  assign o[43302] = i[84];
  assign o[43303] = i[84];
  assign o[43304] = i[84];
  assign o[43305] = i[84];
  assign o[43306] = i[84];
  assign o[43307] = i[84];
  assign o[43308] = i[84];
  assign o[43309] = i[84];
  assign o[43310] = i[84];
  assign o[43311] = i[84];
  assign o[43312] = i[84];
  assign o[43313] = i[84];
  assign o[43314] = i[84];
  assign o[43315] = i[84];
  assign o[43316] = i[84];
  assign o[43317] = i[84];
  assign o[43318] = i[84];
  assign o[43319] = i[84];
  assign o[43320] = i[84];
  assign o[43321] = i[84];
  assign o[43322] = i[84];
  assign o[43323] = i[84];
  assign o[43324] = i[84];
  assign o[43325] = i[84];
  assign o[43326] = i[84];
  assign o[43327] = i[84];
  assign o[43328] = i[84];
  assign o[43329] = i[84];
  assign o[43330] = i[84];
  assign o[43331] = i[84];
  assign o[43332] = i[84];
  assign o[43333] = i[84];
  assign o[43334] = i[84];
  assign o[43335] = i[84];
  assign o[43336] = i[84];
  assign o[43337] = i[84];
  assign o[43338] = i[84];
  assign o[43339] = i[84];
  assign o[43340] = i[84];
  assign o[43341] = i[84];
  assign o[43342] = i[84];
  assign o[43343] = i[84];
  assign o[43344] = i[84];
  assign o[43345] = i[84];
  assign o[43346] = i[84];
  assign o[43347] = i[84];
  assign o[43348] = i[84];
  assign o[43349] = i[84];
  assign o[43350] = i[84];
  assign o[43351] = i[84];
  assign o[43352] = i[84];
  assign o[43353] = i[84];
  assign o[43354] = i[84];
  assign o[43355] = i[84];
  assign o[43356] = i[84];
  assign o[43357] = i[84];
  assign o[43358] = i[84];
  assign o[43359] = i[84];
  assign o[43360] = i[84];
  assign o[43361] = i[84];
  assign o[43362] = i[84];
  assign o[43363] = i[84];
  assign o[43364] = i[84];
  assign o[43365] = i[84];
  assign o[43366] = i[84];
  assign o[43367] = i[84];
  assign o[43368] = i[84];
  assign o[43369] = i[84];
  assign o[43370] = i[84];
  assign o[43371] = i[84];
  assign o[43372] = i[84];
  assign o[43373] = i[84];
  assign o[43374] = i[84];
  assign o[43375] = i[84];
  assign o[43376] = i[84];
  assign o[43377] = i[84];
  assign o[43378] = i[84];
  assign o[43379] = i[84];
  assign o[43380] = i[84];
  assign o[43381] = i[84];
  assign o[43382] = i[84];
  assign o[43383] = i[84];
  assign o[43384] = i[84];
  assign o[43385] = i[84];
  assign o[43386] = i[84];
  assign o[43387] = i[84];
  assign o[43388] = i[84];
  assign o[43389] = i[84];
  assign o[43390] = i[84];
  assign o[43391] = i[84];
  assign o[43392] = i[84];
  assign o[43393] = i[84];
  assign o[43394] = i[84];
  assign o[43395] = i[84];
  assign o[43396] = i[84];
  assign o[43397] = i[84];
  assign o[43398] = i[84];
  assign o[43399] = i[84];
  assign o[43400] = i[84];
  assign o[43401] = i[84];
  assign o[43402] = i[84];
  assign o[43403] = i[84];
  assign o[43404] = i[84];
  assign o[43405] = i[84];
  assign o[43406] = i[84];
  assign o[43407] = i[84];
  assign o[43408] = i[84];
  assign o[43409] = i[84];
  assign o[43410] = i[84];
  assign o[43411] = i[84];
  assign o[43412] = i[84];
  assign o[43413] = i[84];
  assign o[43414] = i[84];
  assign o[43415] = i[84];
  assign o[43416] = i[84];
  assign o[43417] = i[84];
  assign o[43418] = i[84];
  assign o[43419] = i[84];
  assign o[43420] = i[84];
  assign o[43421] = i[84];
  assign o[43422] = i[84];
  assign o[43423] = i[84];
  assign o[43424] = i[84];
  assign o[43425] = i[84];
  assign o[43426] = i[84];
  assign o[43427] = i[84];
  assign o[43428] = i[84];
  assign o[43429] = i[84];
  assign o[43430] = i[84];
  assign o[43431] = i[84];
  assign o[43432] = i[84];
  assign o[43433] = i[84];
  assign o[43434] = i[84];
  assign o[43435] = i[84];
  assign o[43436] = i[84];
  assign o[43437] = i[84];
  assign o[43438] = i[84];
  assign o[43439] = i[84];
  assign o[43440] = i[84];
  assign o[43441] = i[84];
  assign o[43442] = i[84];
  assign o[43443] = i[84];
  assign o[43444] = i[84];
  assign o[43445] = i[84];
  assign o[43446] = i[84];
  assign o[43447] = i[84];
  assign o[43448] = i[84];
  assign o[43449] = i[84];
  assign o[43450] = i[84];
  assign o[43451] = i[84];
  assign o[43452] = i[84];
  assign o[43453] = i[84];
  assign o[43454] = i[84];
  assign o[43455] = i[84];
  assign o[43456] = i[84];
  assign o[43457] = i[84];
  assign o[43458] = i[84];
  assign o[43459] = i[84];
  assign o[43460] = i[84];
  assign o[43461] = i[84];
  assign o[43462] = i[84];
  assign o[43463] = i[84];
  assign o[43464] = i[84];
  assign o[43465] = i[84];
  assign o[43466] = i[84];
  assign o[43467] = i[84];
  assign o[43468] = i[84];
  assign o[43469] = i[84];
  assign o[43470] = i[84];
  assign o[43471] = i[84];
  assign o[43472] = i[84];
  assign o[43473] = i[84];
  assign o[43474] = i[84];
  assign o[43475] = i[84];
  assign o[43476] = i[84];
  assign o[43477] = i[84];
  assign o[43478] = i[84];
  assign o[43479] = i[84];
  assign o[43480] = i[84];
  assign o[43481] = i[84];
  assign o[43482] = i[84];
  assign o[43483] = i[84];
  assign o[43484] = i[84];
  assign o[43485] = i[84];
  assign o[43486] = i[84];
  assign o[43487] = i[84];
  assign o[43488] = i[84];
  assign o[43489] = i[84];
  assign o[43490] = i[84];
  assign o[43491] = i[84];
  assign o[43492] = i[84];
  assign o[43493] = i[84];
  assign o[43494] = i[84];
  assign o[43495] = i[84];
  assign o[43496] = i[84];
  assign o[43497] = i[84];
  assign o[43498] = i[84];
  assign o[43499] = i[84];
  assign o[43500] = i[84];
  assign o[43501] = i[84];
  assign o[43502] = i[84];
  assign o[43503] = i[84];
  assign o[43504] = i[84];
  assign o[43505] = i[84];
  assign o[43506] = i[84];
  assign o[43507] = i[84];
  assign o[43508] = i[84];
  assign o[43509] = i[84];
  assign o[43510] = i[84];
  assign o[43511] = i[84];
  assign o[43512] = i[84];
  assign o[43513] = i[84];
  assign o[43514] = i[84];
  assign o[43515] = i[84];
  assign o[43516] = i[84];
  assign o[43517] = i[84];
  assign o[43518] = i[84];
  assign o[43519] = i[84];
  assign o[42496] = i[83];
  assign o[42497] = i[83];
  assign o[42498] = i[83];
  assign o[42499] = i[83];
  assign o[42500] = i[83];
  assign o[42501] = i[83];
  assign o[42502] = i[83];
  assign o[42503] = i[83];
  assign o[42504] = i[83];
  assign o[42505] = i[83];
  assign o[42506] = i[83];
  assign o[42507] = i[83];
  assign o[42508] = i[83];
  assign o[42509] = i[83];
  assign o[42510] = i[83];
  assign o[42511] = i[83];
  assign o[42512] = i[83];
  assign o[42513] = i[83];
  assign o[42514] = i[83];
  assign o[42515] = i[83];
  assign o[42516] = i[83];
  assign o[42517] = i[83];
  assign o[42518] = i[83];
  assign o[42519] = i[83];
  assign o[42520] = i[83];
  assign o[42521] = i[83];
  assign o[42522] = i[83];
  assign o[42523] = i[83];
  assign o[42524] = i[83];
  assign o[42525] = i[83];
  assign o[42526] = i[83];
  assign o[42527] = i[83];
  assign o[42528] = i[83];
  assign o[42529] = i[83];
  assign o[42530] = i[83];
  assign o[42531] = i[83];
  assign o[42532] = i[83];
  assign o[42533] = i[83];
  assign o[42534] = i[83];
  assign o[42535] = i[83];
  assign o[42536] = i[83];
  assign o[42537] = i[83];
  assign o[42538] = i[83];
  assign o[42539] = i[83];
  assign o[42540] = i[83];
  assign o[42541] = i[83];
  assign o[42542] = i[83];
  assign o[42543] = i[83];
  assign o[42544] = i[83];
  assign o[42545] = i[83];
  assign o[42546] = i[83];
  assign o[42547] = i[83];
  assign o[42548] = i[83];
  assign o[42549] = i[83];
  assign o[42550] = i[83];
  assign o[42551] = i[83];
  assign o[42552] = i[83];
  assign o[42553] = i[83];
  assign o[42554] = i[83];
  assign o[42555] = i[83];
  assign o[42556] = i[83];
  assign o[42557] = i[83];
  assign o[42558] = i[83];
  assign o[42559] = i[83];
  assign o[42560] = i[83];
  assign o[42561] = i[83];
  assign o[42562] = i[83];
  assign o[42563] = i[83];
  assign o[42564] = i[83];
  assign o[42565] = i[83];
  assign o[42566] = i[83];
  assign o[42567] = i[83];
  assign o[42568] = i[83];
  assign o[42569] = i[83];
  assign o[42570] = i[83];
  assign o[42571] = i[83];
  assign o[42572] = i[83];
  assign o[42573] = i[83];
  assign o[42574] = i[83];
  assign o[42575] = i[83];
  assign o[42576] = i[83];
  assign o[42577] = i[83];
  assign o[42578] = i[83];
  assign o[42579] = i[83];
  assign o[42580] = i[83];
  assign o[42581] = i[83];
  assign o[42582] = i[83];
  assign o[42583] = i[83];
  assign o[42584] = i[83];
  assign o[42585] = i[83];
  assign o[42586] = i[83];
  assign o[42587] = i[83];
  assign o[42588] = i[83];
  assign o[42589] = i[83];
  assign o[42590] = i[83];
  assign o[42591] = i[83];
  assign o[42592] = i[83];
  assign o[42593] = i[83];
  assign o[42594] = i[83];
  assign o[42595] = i[83];
  assign o[42596] = i[83];
  assign o[42597] = i[83];
  assign o[42598] = i[83];
  assign o[42599] = i[83];
  assign o[42600] = i[83];
  assign o[42601] = i[83];
  assign o[42602] = i[83];
  assign o[42603] = i[83];
  assign o[42604] = i[83];
  assign o[42605] = i[83];
  assign o[42606] = i[83];
  assign o[42607] = i[83];
  assign o[42608] = i[83];
  assign o[42609] = i[83];
  assign o[42610] = i[83];
  assign o[42611] = i[83];
  assign o[42612] = i[83];
  assign o[42613] = i[83];
  assign o[42614] = i[83];
  assign o[42615] = i[83];
  assign o[42616] = i[83];
  assign o[42617] = i[83];
  assign o[42618] = i[83];
  assign o[42619] = i[83];
  assign o[42620] = i[83];
  assign o[42621] = i[83];
  assign o[42622] = i[83];
  assign o[42623] = i[83];
  assign o[42624] = i[83];
  assign o[42625] = i[83];
  assign o[42626] = i[83];
  assign o[42627] = i[83];
  assign o[42628] = i[83];
  assign o[42629] = i[83];
  assign o[42630] = i[83];
  assign o[42631] = i[83];
  assign o[42632] = i[83];
  assign o[42633] = i[83];
  assign o[42634] = i[83];
  assign o[42635] = i[83];
  assign o[42636] = i[83];
  assign o[42637] = i[83];
  assign o[42638] = i[83];
  assign o[42639] = i[83];
  assign o[42640] = i[83];
  assign o[42641] = i[83];
  assign o[42642] = i[83];
  assign o[42643] = i[83];
  assign o[42644] = i[83];
  assign o[42645] = i[83];
  assign o[42646] = i[83];
  assign o[42647] = i[83];
  assign o[42648] = i[83];
  assign o[42649] = i[83];
  assign o[42650] = i[83];
  assign o[42651] = i[83];
  assign o[42652] = i[83];
  assign o[42653] = i[83];
  assign o[42654] = i[83];
  assign o[42655] = i[83];
  assign o[42656] = i[83];
  assign o[42657] = i[83];
  assign o[42658] = i[83];
  assign o[42659] = i[83];
  assign o[42660] = i[83];
  assign o[42661] = i[83];
  assign o[42662] = i[83];
  assign o[42663] = i[83];
  assign o[42664] = i[83];
  assign o[42665] = i[83];
  assign o[42666] = i[83];
  assign o[42667] = i[83];
  assign o[42668] = i[83];
  assign o[42669] = i[83];
  assign o[42670] = i[83];
  assign o[42671] = i[83];
  assign o[42672] = i[83];
  assign o[42673] = i[83];
  assign o[42674] = i[83];
  assign o[42675] = i[83];
  assign o[42676] = i[83];
  assign o[42677] = i[83];
  assign o[42678] = i[83];
  assign o[42679] = i[83];
  assign o[42680] = i[83];
  assign o[42681] = i[83];
  assign o[42682] = i[83];
  assign o[42683] = i[83];
  assign o[42684] = i[83];
  assign o[42685] = i[83];
  assign o[42686] = i[83];
  assign o[42687] = i[83];
  assign o[42688] = i[83];
  assign o[42689] = i[83];
  assign o[42690] = i[83];
  assign o[42691] = i[83];
  assign o[42692] = i[83];
  assign o[42693] = i[83];
  assign o[42694] = i[83];
  assign o[42695] = i[83];
  assign o[42696] = i[83];
  assign o[42697] = i[83];
  assign o[42698] = i[83];
  assign o[42699] = i[83];
  assign o[42700] = i[83];
  assign o[42701] = i[83];
  assign o[42702] = i[83];
  assign o[42703] = i[83];
  assign o[42704] = i[83];
  assign o[42705] = i[83];
  assign o[42706] = i[83];
  assign o[42707] = i[83];
  assign o[42708] = i[83];
  assign o[42709] = i[83];
  assign o[42710] = i[83];
  assign o[42711] = i[83];
  assign o[42712] = i[83];
  assign o[42713] = i[83];
  assign o[42714] = i[83];
  assign o[42715] = i[83];
  assign o[42716] = i[83];
  assign o[42717] = i[83];
  assign o[42718] = i[83];
  assign o[42719] = i[83];
  assign o[42720] = i[83];
  assign o[42721] = i[83];
  assign o[42722] = i[83];
  assign o[42723] = i[83];
  assign o[42724] = i[83];
  assign o[42725] = i[83];
  assign o[42726] = i[83];
  assign o[42727] = i[83];
  assign o[42728] = i[83];
  assign o[42729] = i[83];
  assign o[42730] = i[83];
  assign o[42731] = i[83];
  assign o[42732] = i[83];
  assign o[42733] = i[83];
  assign o[42734] = i[83];
  assign o[42735] = i[83];
  assign o[42736] = i[83];
  assign o[42737] = i[83];
  assign o[42738] = i[83];
  assign o[42739] = i[83];
  assign o[42740] = i[83];
  assign o[42741] = i[83];
  assign o[42742] = i[83];
  assign o[42743] = i[83];
  assign o[42744] = i[83];
  assign o[42745] = i[83];
  assign o[42746] = i[83];
  assign o[42747] = i[83];
  assign o[42748] = i[83];
  assign o[42749] = i[83];
  assign o[42750] = i[83];
  assign o[42751] = i[83];
  assign o[42752] = i[83];
  assign o[42753] = i[83];
  assign o[42754] = i[83];
  assign o[42755] = i[83];
  assign o[42756] = i[83];
  assign o[42757] = i[83];
  assign o[42758] = i[83];
  assign o[42759] = i[83];
  assign o[42760] = i[83];
  assign o[42761] = i[83];
  assign o[42762] = i[83];
  assign o[42763] = i[83];
  assign o[42764] = i[83];
  assign o[42765] = i[83];
  assign o[42766] = i[83];
  assign o[42767] = i[83];
  assign o[42768] = i[83];
  assign o[42769] = i[83];
  assign o[42770] = i[83];
  assign o[42771] = i[83];
  assign o[42772] = i[83];
  assign o[42773] = i[83];
  assign o[42774] = i[83];
  assign o[42775] = i[83];
  assign o[42776] = i[83];
  assign o[42777] = i[83];
  assign o[42778] = i[83];
  assign o[42779] = i[83];
  assign o[42780] = i[83];
  assign o[42781] = i[83];
  assign o[42782] = i[83];
  assign o[42783] = i[83];
  assign o[42784] = i[83];
  assign o[42785] = i[83];
  assign o[42786] = i[83];
  assign o[42787] = i[83];
  assign o[42788] = i[83];
  assign o[42789] = i[83];
  assign o[42790] = i[83];
  assign o[42791] = i[83];
  assign o[42792] = i[83];
  assign o[42793] = i[83];
  assign o[42794] = i[83];
  assign o[42795] = i[83];
  assign o[42796] = i[83];
  assign o[42797] = i[83];
  assign o[42798] = i[83];
  assign o[42799] = i[83];
  assign o[42800] = i[83];
  assign o[42801] = i[83];
  assign o[42802] = i[83];
  assign o[42803] = i[83];
  assign o[42804] = i[83];
  assign o[42805] = i[83];
  assign o[42806] = i[83];
  assign o[42807] = i[83];
  assign o[42808] = i[83];
  assign o[42809] = i[83];
  assign o[42810] = i[83];
  assign o[42811] = i[83];
  assign o[42812] = i[83];
  assign o[42813] = i[83];
  assign o[42814] = i[83];
  assign o[42815] = i[83];
  assign o[42816] = i[83];
  assign o[42817] = i[83];
  assign o[42818] = i[83];
  assign o[42819] = i[83];
  assign o[42820] = i[83];
  assign o[42821] = i[83];
  assign o[42822] = i[83];
  assign o[42823] = i[83];
  assign o[42824] = i[83];
  assign o[42825] = i[83];
  assign o[42826] = i[83];
  assign o[42827] = i[83];
  assign o[42828] = i[83];
  assign o[42829] = i[83];
  assign o[42830] = i[83];
  assign o[42831] = i[83];
  assign o[42832] = i[83];
  assign o[42833] = i[83];
  assign o[42834] = i[83];
  assign o[42835] = i[83];
  assign o[42836] = i[83];
  assign o[42837] = i[83];
  assign o[42838] = i[83];
  assign o[42839] = i[83];
  assign o[42840] = i[83];
  assign o[42841] = i[83];
  assign o[42842] = i[83];
  assign o[42843] = i[83];
  assign o[42844] = i[83];
  assign o[42845] = i[83];
  assign o[42846] = i[83];
  assign o[42847] = i[83];
  assign o[42848] = i[83];
  assign o[42849] = i[83];
  assign o[42850] = i[83];
  assign o[42851] = i[83];
  assign o[42852] = i[83];
  assign o[42853] = i[83];
  assign o[42854] = i[83];
  assign o[42855] = i[83];
  assign o[42856] = i[83];
  assign o[42857] = i[83];
  assign o[42858] = i[83];
  assign o[42859] = i[83];
  assign o[42860] = i[83];
  assign o[42861] = i[83];
  assign o[42862] = i[83];
  assign o[42863] = i[83];
  assign o[42864] = i[83];
  assign o[42865] = i[83];
  assign o[42866] = i[83];
  assign o[42867] = i[83];
  assign o[42868] = i[83];
  assign o[42869] = i[83];
  assign o[42870] = i[83];
  assign o[42871] = i[83];
  assign o[42872] = i[83];
  assign o[42873] = i[83];
  assign o[42874] = i[83];
  assign o[42875] = i[83];
  assign o[42876] = i[83];
  assign o[42877] = i[83];
  assign o[42878] = i[83];
  assign o[42879] = i[83];
  assign o[42880] = i[83];
  assign o[42881] = i[83];
  assign o[42882] = i[83];
  assign o[42883] = i[83];
  assign o[42884] = i[83];
  assign o[42885] = i[83];
  assign o[42886] = i[83];
  assign o[42887] = i[83];
  assign o[42888] = i[83];
  assign o[42889] = i[83];
  assign o[42890] = i[83];
  assign o[42891] = i[83];
  assign o[42892] = i[83];
  assign o[42893] = i[83];
  assign o[42894] = i[83];
  assign o[42895] = i[83];
  assign o[42896] = i[83];
  assign o[42897] = i[83];
  assign o[42898] = i[83];
  assign o[42899] = i[83];
  assign o[42900] = i[83];
  assign o[42901] = i[83];
  assign o[42902] = i[83];
  assign o[42903] = i[83];
  assign o[42904] = i[83];
  assign o[42905] = i[83];
  assign o[42906] = i[83];
  assign o[42907] = i[83];
  assign o[42908] = i[83];
  assign o[42909] = i[83];
  assign o[42910] = i[83];
  assign o[42911] = i[83];
  assign o[42912] = i[83];
  assign o[42913] = i[83];
  assign o[42914] = i[83];
  assign o[42915] = i[83];
  assign o[42916] = i[83];
  assign o[42917] = i[83];
  assign o[42918] = i[83];
  assign o[42919] = i[83];
  assign o[42920] = i[83];
  assign o[42921] = i[83];
  assign o[42922] = i[83];
  assign o[42923] = i[83];
  assign o[42924] = i[83];
  assign o[42925] = i[83];
  assign o[42926] = i[83];
  assign o[42927] = i[83];
  assign o[42928] = i[83];
  assign o[42929] = i[83];
  assign o[42930] = i[83];
  assign o[42931] = i[83];
  assign o[42932] = i[83];
  assign o[42933] = i[83];
  assign o[42934] = i[83];
  assign o[42935] = i[83];
  assign o[42936] = i[83];
  assign o[42937] = i[83];
  assign o[42938] = i[83];
  assign o[42939] = i[83];
  assign o[42940] = i[83];
  assign o[42941] = i[83];
  assign o[42942] = i[83];
  assign o[42943] = i[83];
  assign o[42944] = i[83];
  assign o[42945] = i[83];
  assign o[42946] = i[83];
  assign o[42947] = i[83];
  assign o[42948] = i[83];
  assign o[42949] = i[83];
  assign o[42950] = i[83];
  assign o[42951] = i[83];
  assign o[42952] = i[83];
  assign o[42953] = i[83];
  assign o[42954] = i[83];
  assign o[42955] = i[83];
  assign o[42956] = i[83];
  assign o[42957] = i[83];
  assign o[42958] = i[83];
  assign o[42959] = i[83];
  assign o[42960] = i[83];
  assign o[42961] = i[83];
  assign o[42962] = i[83];
  assign o[42963] = i[83];
  assign o[42964] = i[83];
  assign o[42965] = i[83];
  assign o[42966] = i[83];
  assign o[42967] = i[83];
  assign o[42968] = i[83];
  assign o[42969] = i[83];
  assign o[42970] = i[83];
  assign o[42971] = i[83];
  assign o[42972] = i[83];
  assign o[42973] = i[83];
  assign o[42974] = i[83];
  assign o[42975] = i[83];
  assign o[42976] = i[83];
  assign o[42977] = i[83];
  assign o[42978] = i[83];
  assign o[42979] = i[83];
  assign o[42980] = i[83];
  assign o[42981] = i[83];
  assign o[42982] = i[83];
  assign o[42983] = i[83];
  assign o[42984] = i[83];
  assign o[42985] = i[83];
  assign o[42986] = i[83];
  assign o[42987] = i[83];
  assign o[42988] = i[83];
  assign o[42989] = i[83];
  assign o[42990] = i[83];
  assign o[42991] = i[83];
  assign o[42992] = i[83];
  assign o[42993] = i[83];
  assign o[42994] = i[83];
  assign o[42995] = i[83];
  assign o[42996] = i[83];
  assign o[42997] = i[83];
  assign o[42998] = i[83];
  assign o[42999] = i[83];
  assign o[43000] = i[83];
  assign o[43001] = i[83];
  assign o[43002] = i[83];
  assign o[43003] = i[83];
  assign o[43004] = i[83];
  assign o[43005] = i[83];
  assign o[43006] = i[83];
  assign o[43007] = i[83];
  assign o[41984] = i[82];
  assign o[41985] = i[82];
  assign o[41986] = i[82];
  assign o[41987] = i[82];
  assign o[41988] = i[82];
  assign o[41989] = i[82];
  assign o[41990] = i[82];
  assign o[41991] = i[82];
  assign o[41992] = i[82];
  assign o[41993] = i[82];
  assign o[41994] = i[82];
  assign o[41995] = i[82];
  assign o[41996] = i[82];
  assign o[41997] = i[82];
  assign o[41998] = i[82];
  assign o[41999] = i[82];
  assign o[42000] = i[82];
  assign o[42001] = i[82];
  assign o[42002] = i[82];
  assign o[42003] = i[82];
  assign o[42004] = i[82];
  assign o[42005] = i[82];
  assign o[42006] = i[82];
  assign o[42007] = i[82];
  assign o[42008] = i[82];
  assign o[42009] = i[82];
  assign o[42010] = i[82];
  assign o[42011] = i[82];
  assign o[42012] = i[82];
  assign o[42013] = i[82];
  assign o[42014] = i[82];
  assign o[42015] = i[82];
  assign o[42016] = i[82];
  assign o[42017] = i[82];
  assign o[42018] = i[82];
  assign o[42019] = i[82];
  assign o[42020] = i[82];
  assign o[42021] = i[82];
  assign o[42022] = i[82];
  assign o[42023] = i[82];
  assign o[42024] = i[82];
  assign o[42025] = i[82];
  assign o[42026] = i[82];
  assign o[42027] = i[82];
  assign o[42028] = i[82];
  assign o[42029] = i[82];
  assign o[42030] = i[82];
  assign o[42031] = i[82];
  assign o[42032] = i[82];
  assign o[42033] = i[82];
  assign o[42034] = i[82];
  assign o[42035] = i[82];
  assign o[42036] = i[82];
  assign o[42037] = i[82];
  assign o[42038] = i[82];
  assign o[42039] = i[82];
  assign o[42040] = i[82];
  assign o[42041] = i[82];
  assign o[42042] = i[82];
  assign o[42043] = i[82];
  assign o[42044] = i[82];
  assign o[42045] = i[82];
  assign o[42046] = i[82];
  assign o[42047] = i[82];
  assign o[42048] = i[82];
  assign o[42049] = i[82];
  assign o[42050] = i[82];
  assign o[42051] = i[82];
  assign o[42052] = i[82];
  assign o[42053] = i[82];
  assign o[42054] = i[82];
  assign o[42055] = i[82];
  assign o[42056] = i[82];
  assign o[42057] = i[82];
  assign o[42058] = i[82];
  assign o[42059] = i[82];
  assign o[42060] = i[82];
  assign o[42061] = i[82];
  assign o[42062] = i[82];
  assign o[42063] = i[82];
  assign o[42064] = i[82];
  assign o[42065] = i[82];
  assign o[42066] = i[82];
  assign o[42067] = i[82];
  assign o[42068] = i[82];
  assign o[42069] = i[82];
  assign o[42070] = i[82];
  assign o[42071] = i[82];
  assign o[42072] = i[82];
  assign o[42073] = i[82];
  assign o[42074] = i[82];
  assign o[42075] = i[82];
  assign o[42076] = i[82];
  assign o[42077] = i[82];
  assign o[42078] = i[82];
  assign o[42079] = i[82];
  assign o[42080] = i[82];
  assign o[42081] = i[82];
  assign o[42082] = i[82];
  assign o[42083] = i[82];
  assign o[42084] = i[82];
  assign o[42085] = i[82];
  assign o[42086] = i[82];
  assign o[42087] = i[82];
  assign o[42088] = i[82];
  assign o[42089] = i[82];
  assign o[42090] = i[82];
  assign o[42091] = i[82];
  assign o[42092] = i[82];
  assign o[42093] = i[82];
  assign o[42094] = i[82];
  assign o[42095] = i[82];
  assign o[42096] = i[82];
  assign o[42097] = i[82];
  assign o[42098] = i[82];
  assign o[42099] = i[82];
  assign o[42100] = i[82];
  assign o[42101] = i[82];
  assign o[42102] = i[82];
  assign o[42103] = i[82];
  assign o[42104] = i[82];
  assign o[42105] = i[82];
  assign o[42106] = i[82];
  assign o[42107] = i[82];
  assign o[42108] = i[82];
  assign o[42109] = i[82];
  assign o[42110] = i[82];
  assign o[42111] = i[82];
  assign o[42112] = i[82];
  assign o[42113] = i[82];
  assign o[42114] = i[82];
  assign o[42115] = i[82];
  assign o[42116] = i[82];
  assign o[42117] = i[82];
  assign o[42118] = i[82];
  assign o[42119] = i[82];
  assign o[42120] = i[82];
  assign o[42121] = i[82];
  assign o[42122] = i[82];
  assign o[42123] = i[82];
  assign o[42124] = i[82];
  assign o[42125] = i[82];
  assign o[42126] = i[82];
  assign o[42127] = i[82];
  assign o[42128] = i[82];
  assign o[42129] = i[82];
  assign o[42130] = i[82];
  assign o[42131] = i[82];
  assign o[42132] = i[82];
  assign o[42133] = i[82];
  assign o[42134] = i[82];
  assign o[42135] = i[82];
  assign o[42136] = i[82];
  assign o[42137] = i[82];
  assign o[42138] = i[82];
  assign o[42139] = i[82];
  assign o[42140] = i[82];
  assign o[42141] = i[82];
  assign o[42142] = i[82];
  assign o[42143] = i[82];
  assign o[42144] = i[82];
  assign o[42145] = i[82];
  assign o[42146] = i[82];
  assign o[42147] = i[82];
  assign o[42148] = i[82];
  assign o[42149] = i[82];
  assign o[42150] = i[82];
  assign o[42151] = i[82];
  assign o[42152] = i[82];
  assign o[42153] = i[82];
  assign o[42154] = i[82];
  assign o[42155] = i[82];
  assign o[42156] = i[82];
  assign o[42157] = i[82];
  assign o[42158] = i[82];
  assign o[42159] = i[82];
  assign o[42160] = i[82];
  assign o[42161] = i[82];
  assign o[42162] = i[82];
  assign o[42163] = i[82];
  assign o[42164] = i[82];
  assign o[42165] = i[82];
  assign o[42166] = i[82];
  assign o[42167] = i[82];
  assign o[42168] = i[82];
  assign o[42169] = i[82];
  assign o[42170] = i[82];
  assign o[42171] = i[82];
  assign o[42172] = i[82];
  assign o[42173] = i[82];
  assign o[42174] = i[82];
  assign o[42175] = i[82];
  assign o[42176] = i[82];
  assign o[42177] = i[82];
  assign o[42178] = i[82];
  assign o[42179] = i[82];
  assign o[42180] = i[82];
  assign o[42181] = i[82];
  assign o[42182] = i[82];
  assign o[42183] = i[82];
  assign o[42184] = i[82];
  assign o[42185] = i[82];
  assign o[42186] = i[82];
  assign o[42187] = i[82];
  assign o[42188] = i[82];
  assign o[42189] = i[82];
  assign o[42190] = i[82];
  assign o[42191] = i[82];
  assign o[42192] = i[82];
  assign o[42193] = i[82];
  assign o[42194] = i[82];
  assign o[42195] = i[82];
  assign o[42196] = i[82];
  assign o[42197] = i[82];
  assign o[42198] = i[82];
  assign o[42199] = i[82];
  assign o[42200] = i[82];
  assign o[42201] = i[82];
  assign o[42202] = i[82];
  assign o[42203] = i[82];
  assign o[42204] = i[82];
  assign o[42205] = i[82];
  assign o[42206] = i[82];
  assign o[42207] = i[82];
  assign o[42208] = i[82];
  assign o[42209] = i[82];
  assign o[42210] = i[82];
  assign o[42211] = i[82];
  assign o[42212] = i[82];
  assign o[42213] = i[82];
  assign o[42214] = i[82];
  assign o[42215] = i[82];
  assign o[42216] = i[82];
  assign o[42217] = i[82];
  assign o[42218] = i[82];
  assign o[42219] = i[82];
  assign o[42220] = i[82];
  assign o[42221] = i[82];
  assign o[42222] = i[82];
  assign o[42223] = i[82];
  assign o[42224] = i[82];
  assign o[42225] = i[82];
  assign o[42226] = i[82];
  assign o[42227] = i[82];
  assign o[42228] = i[82];
  assign o[42229] = i[82];
  assign o[42230] = i[82];
  assign o[42231] = i[82];
  assign o[42232] = i[82];
  assign o[42233] = i[82];
  assign o[42234] = i[82];
  assign o[42235] = i[82];
  assign o[42236] = i[82];
  assign o[42237] = i[82];
  assign o[42238] = i[82];
  assign o[42239] = i[82];
  assign o[42240] = i[82];
  assign o[42241] = i[82];
  assign o[42242] = i[82];
  assign o[42243] = i[82];
  assign o[42244] = i[82];
  assign o[42245] = i[82];
  assign o[42246] = i[82];
  assign o[42247] = i[82];
  assign o[42248] = i[82];
  assign o[42249] = i[82];
  assign o[42250] = i[82];
  assign o[42251] = i[82];
  assign o[42252] = i[82];
  assign o[42253] = i[82];
  assign o[42254] = i[82];
  assign o[42255] = i[82];
  assign o[42256] = i[82];
  assign o[42257] = i[82];
  assign o[42258] = i[82];
  assign o[42259] = i[82];
  assign o[42260] = i[82];
  assign o[42261] = i[82];
  assign o[42262] = i[82];
  assign o[42263] = i[82];
  assign o[42264] = i[82];
  assign o[42265] = i[82];
  assign o[42266] = i[82];
  assign o[42267] = i[82];
  assign o[42268] = i[82];
  assign o[42269] = i[82];
  assign o[42270] = i[82];
  assign o[42271] = i[82];
  assign o[42272] = i[82];
  assign o[42273] = i[82];
  assign o[42274] = i[82];
  assign o[42275] = i[82];
  assign o[42276] = i[82];
  assign o[42277] = i[82];
  assign o[42278] = i[82];
  assign o[42279] = i[82];
  assign o[42280] = i[82];
  assign o[42281] = i[82];
  assign o[42282] = i[82];
  assign o[42283] = i[82];
  assign o[42284] = i[82];
  assign o[42285] = i[82];
  assign o[42286] = i[82];
  assign o[42287] = i[82];
  assign o[42288] = i[82];
  assign o[42289] = i[82];
  assign o[42290] = i[82];
  assign o[42291] = i[82];
  assign o[42292] = i[82];
  assign o[42293] = i[82];
  assign o[42294] = i[82];
  assign o[42295] = i[82];
  assign o[42296] = i[82];
  assign o[42297] = i[82];
  assign o[42298] = i[82];
  assign o[42299] = i[82];
  assign o[42300] = i[82];
  assign o[42301] = i[82];
  assign o[42302] = i[82];
  assign o[42303] = i[82];
  assign o[42304] = i[82];
  assign o[42305] = i[82];
  assign o[42306] = i[82];
  assign o[42307] = i[82];
  assign o[42308] = i[82];
  assign o[42309] = i[82];
  assign o[42310] = i[82];
  assign o[42311] = i[82];
  assign o[42312] = i[82];
  assign o[42313] = i[82];
  assign o[42314] = i[82];
  assign o[42315] = i[82];
  assign o[42316] = i[82];
  assign o[42317] = i[82];
  assign o[42318] = i[82];
  assign o[42319] = i[82];
  assign o[42320] = i[82];
  assign o[42321] = i[82];
  assign o[42322] = i[82];
  assign o[42323] = i[82];
  assign o[42324] = i[82];
  assign o[42325] = i[82];
  assign o[42326] = i[82];
  assign o[42327] = i[82];
  assign o[42328] = i[82];
  assign o[42329] = i[82];
  assign o[42330] = i[82];
  assign o[42331] = i[82];
  assign o[42332] = i[82];
  assign o[42333] = i[82];
  assign o[42334] = i[82];
  assign o[42335] = i[82];
  assign o[42336] = i[82];
  assign o[42337] = i[82];
  assign o[42338] = i[82];
  assign o[42339] = i[82];
  assign o[42340] = i[82];
  assign o[42341] = i[82];
  assign o[42342] = i[82];
  assign o[42343] = i[82];
  assign o[42344] = i[82];
  assign o[42345] = i[82];
  assign o[42346] = i[82];
  assign o[42347] = i[82];
  assign o[42348] = i[82];
  assign o[42349] = i[82];
  assign o[42350] = i[82];
  assign o[42351] = i[82];
  assign o[42352] = i[82];
  assign o[42353] = i[82];
  assign o[42354] = i[82];
  assign o[42355] = i[82];
  assign o[42356] = i[82];
  assign o[42357] = i[82];
  assign o[42358] = i[82];
  assign o[42359] = i[82];
  assign o[42360] = i[82];
  assign o[42361] = i[82];
  assign o[42362] = i[82];
  assign o[42363] = i[82];
  assign o[42364] = i[82];
  assign o[42365] = i[82];
  assign o[42366] = i[82];
  assign o[42367] = i[82];
  assign o[42368] = i[82];
  assign o[42369] = i[82];
  assign o[42370] = i[82];
  assign o[42371] = i[82];
  assign o[42372] = i[82];
  assign o[42373] = i[82];
  assign o[42374] = i[82];
  assign o[42375] = i[82];
  assign o[42376] = i[82];
  assign o[42377] = i[82];
  assign o[42378] = i[82];
  assign o[42379] = i[82];
  assign o[42380] = i[82];
  assign o[42381] = i[82];
  assign o[42382] = i[82];
  assign o[42383] = i[82];
  assign o[42384] = i[82];
  assign o[42385] = i[82];
  assign o[42386] = i[82];
  assign o[42387] = i[82];
  assign o[42388] = i[82];
  assign o[42389] = i[82];
  assign o[42390] = i[82];
  assign o[42391] = i[82];
  assign o[42392] = i[82];
  assign o[42393] = i[82];
  assign o[42394] = i[82];
  assign o[42395] = i[82];
  assign o[42396] = i[82];
  assign o[42397] = i[82];
  assign o[42398] = i[82];
  assign o[42399] = i[82];
  assign o[42400] = i[82];
  assign o[42401] = i[82];
  assign o[42402] = i[82];
  assign o[42403] = i[82];
  assign o[42404] = i[82];
  assign o[42405] = i[82];
  assign o[42406] = i[82];
  assign o[42407] = i[82];
  assign o[42408] = i[82];
  assign o[42409] = i[82];
  assign o[42410] = i[82];
  assign o[42411] = i[82];
  assign o[42412] = i[82];
  assign o[42413] = i[82];
  assign o[42414] = i[82];
  assign o[42415] = i[82];
  assign o[42416] = i[82];
  assign o[42417] = i[82];
  assign o[42418] = i[82];
  assign o[42419] = i[82];
  assign o[42420] = i[82];
  assign o[42421] = i[82];
  assign o[42422] = i[82];
  assign o[42423] = i[82];
  assign o[42424] = i[82];
  assign o[42425] = i[82];
  assign o[42426] = i[82];
  assign o[42427] = i[82];
  assign o[42428] = i[82];
  assign o[42429] = i[82];
  assign o[42430] = i[82];
  assign o[42431] = i[82];
  assign o[42432] = i[82];
  assign o[42433] = i[82];
  assign o[42434] = i[82];
  assign o[42435] = i[82];
  assign o[42436] = i[82];
  assign o[42437] = i[82];
  assign o[42438] = i[82];
  assign o[42439] = i[82];
  assign o[42440] = i[82];
  assign o[42441] = i[82];
  assign o[42442] = i[82];
  assign o[42443] = i[82];
  assign o[42444] = i[82];
  assign o[42445] = i[82];
  assign o[42446] = i[82];
  assign o[42447] = i[82];
  assign o[42448] = i[82];
  assign o[42449] = i[82];
  assign o[42450] = i[82];
  assign o[42451] = i[82];
  assign o[42452] = i[82];
  assign o[42453] = i[82];
  assign o[42454] = i[82];
  assign o[42455] = i[82];
  assign o[42456] = i[82];
  assign o[42457] = i[82];
  assign o[42458] = i[82];
  assign o[42459] = i[82];
  assign o[42460] = i[82];
  assign o[42461] = i[82];
  assign o[42462] = i[82];
  assign o[42463] = i[82];
  assign o[42464] = i[82];
  assign o[42465] = i[82];
  assign o[42466] = i[82];
  assign o[42467] = i[82];
  assign o[42468] = i[82];
  assign o[42469] = i[82];
  assign o[42470] = i[82];
  assign o[42471] = i[82];
  assign o[42472] = i[82];
  assign o[42473] = i[82];
  assign o[42474] = i[82];
  assign o[42475] = i[82];
  assign o[42476] = i[82];
  assign o[42477] = i[82];
  assign o[42478] = i[82];
  assign o[42479] = i[82];
  assign o[42480] = i[82];
  assign o[42481] = i[82];
  assign o[42482] = i[82];
  assign o[42483] = i[82];
  assign o[42484] = i[82];
  assign o[42485] = i[82];
  assign o[42486] = i[82];
  assign o[42487] = i[82];
  assign o[42488] = i[82];
  assign o[42489] = i[82];
  assign o[42490] = i[82];
  assign o[42491] = i[82];
  assign o[42492] = i[82];
  assign o[42493] = i[82];
  assign o[42494] = i[82];
  assign o[42495] = i[82];
  assign o[41472] = i[81];
  assign o[41473] = i[81];
  assign o[41474] = i[81];
  assign o[41475] = i[81];
  assign o[41476] = i[81];
  assign o[41477] = i[81];
  assign o[41478] = i[81];
  assign o[41479] = i[81];
  assign o[41480] = i[81];
  assign o[41481] = i[81];
  assign o[41482] = i[81];
  assign o[41483] = i[81];
  assign o[41484] = i[81];
  assign o[41485] = i[81];
  assign o[41486] = i[81];
  assign o[41487] = i[81];
  assign o[41488] = i[81];
  assign o[41489] = i[81];
  assign o[41490] = i[81];
  assign o[41491] = i[81];
  assign o[41492] = i[81];
  assign o[41493] = i[81];
  assign o[41494] = i[81];
  assign o[41495] = i[81];
  assign o[41496] = i[81];
  assign o[41497] = i[81];
  assign o[41498] = i[81];
  assign o[41499] = i[81];
  assign o[41500] = i[81];
  assign o[41501] = i[81];
  assign o[41502] = i[81];
  assign o[41503] = i[81];
  assign o[41504] = i[81];
  assign o[41505] = i[81];
  assign o[41506] = i[81];
  assign o[41507] = i[81];
  assign o[41508] = i[81];
  assign o[41509] = i[81];
  assign o[41510] = i[81];
  assign o[41511] = i[81];
  assign o[41512] = i[81];
  assign o[41513] = i[81];
  assign o[41514] = i[81];
  assign o[41515] = i[81];
  assign o[41516] = i[81];
  assign o[41517] = i[81];
  assign o[41518] = i[81];
  assign o[41519] = i[81];
  assign o[41520] = i[81];
  assign o[41521] = i[81];
  assign o[41522] = i[81];
  assign o[41523] = i[81];
  assign o[41524] = i[81];
  assign o[41525] = i[81];
  assign o[41526] = i[81];
  assign o[41527] = i[81];
  assign o[41528] = i[81];
  assign o[41529] = i[81];
  assign o[41530] = i[81];
  assign o[41531] = i[81];
  assign o[41532] = i[81];
  assign o[41533] = i[81];
  assign o[41534] = i[81];
  assign o[41535] = i[81];
  assign o[41536] = i[81];
  assign o[41537] = i[81];
  assign o[41538] = i[81];
  assign o[41539] = i[81];
  assign o[41540] = i[81];
  assign o[41541] = i[81];
  assign o[41542] = i[81];
  assign o[41543] = i[81];
  assign o[41544] = i[81];
  assign o[41545] = i[81];
  assign o[41546] = i[81];
  assign o[41547] = i[81];
  assign o[41548] = i[81];
  assign o[41549] = i[81];
  assign o[41550] = i[81];
  assign o[41551] = i[81];
  assign o[41552] = i[81];
  assign o[41553] = i[81];
  assign o[41554] = i[81];
  assign o[41555] = i[81];
  assign o[41556] = i[81];
  assign o[41557] = i[81];
  assign o[41558] = i[81];
  assign o[41559] = i[81];
  assign o[41560] = i[81];
  assign o[41561] = i[81];
  assign o[41562] = i[81];
  assign o[41563] = i[81];
  assign o[41564] = i[81];
  assign o[41565] = i[81];
  assign o[41566] = i[81];
  assign o[41567] = i[81];
  assign o[41568] = i[81];
  assign o[41569] = i[81];
  assign o[41570] = i[81];
  assign o[41571] = i[81];
  assign o[41572] = i[81];
  assign o[41573] = i[81];
  assign o[41574] = i[81];
  assign o[41575] = i[81];
  assign o[41576] = i[81];
  assign o[41577] = i[81];
  assign o[41578] = i[81];
  assign o[41579] = i[81];
  assign o[41580] = i[81];
  assign o[41581] = i[81];
  assign o[41582] = i[81];
  assign o[41583] = i[81];
  assign o[41584] = i[81];
  assign o[41585] = i[81];
  assign o[41586] = i[81];
  assign o[41587] = i[81];
  assign o[41588] = i[81];
  assign o[41589] = i[81];
  assign o[41590] = i[81];
  assign o[41591] = i[81];
  assign o[41592] = i[81];
  assign o[41593] = i[81];
  assign o[41594] = i[81];
  assign o[41595] = i[81];
  assign o[41596] = i[81];
  assign o[41597] = i[81];
  assign o[41598] = i[81];
  assign o[41599] = i[81];
  assign o[41600] = i[81];
  assign o[41601] = i[81];
  assign o[41602] = i[81];
  assign o[41603] = i[81];
  assign o[41604] = i[81];
  assign o[41605] = i[81];
  assign o[41606] = i[81];
  assign o[41607] = i[81];
  assign o[41608] = i[81];
  assign o[41609] = i[81];
  assign o[41610] = i[81];
  assign o[41611] = i[81];
  assign o[41612] = i[81];
  assign o[41613] = i[81];
  assign o[41614] = i[81];
  assign o[41615] = i[81];
  assign o[41616] = i[81];
  assign o[41617] = i[81];
  assign o[41618] = i[81];
  assign o[41619] = i[81];
  assign o[41620] = i[81];
  assign o[41621] = i[81];
  assign o[41622] = i[81];
  assign o[41623] = i[81];
  assign o[41624] = i[81];
  assign o[41625] = i[81];
  assign o[41626] = i[81];
  assign o[41627] = i[81];
  assign o[41628] = i[81];
  assign o[41629] = i[81];
  assign o[41630] = i[81];
  assign o[41631] = i[81];
  assign o[41632] = i[81];
  assign o[41633] = i[81];
  assign o[41634] = i[81];
  assign o[41635] = i[81];
  assign o[41636] = i[81];
  assign o[41637] = i[81];
  assign o[41638] = i[81];
  assign o[41639] = i[81];
  assign o[41640] = i[81];
  assign o[41641] = i[81];
  assign o[41642] = i[81];
  assign o[41643] = i[81];
  assign o[41644] = i[81];
  assign o[41645] = i[81];
  assign o[41646] = i[81];
  assign o[41647] = i[81];
  assign o[41648] = i[81];
  assign o[41649] = i[81];
  assign o[41650] = i[81];
  assign o[41651] = i[81];
  assign o[41652] = i[81];
  assign o[41653] = i[81];
  assign o[41654] = i[81];
  assign o[41655] = i[81];
  assign o[41656] = i[81];
  assign o[41657] = i[81];
  assign o[41658] = i[81];
  assign o[41659] = i[81];
  assign o[41660] = i[81];
  assign o[41661] = i[81];
  assign o[41662] = i[81];
  assign o[41663] = i[81];
  assign o[41664] = i[81];
  assign o[41665] = i[81];
  assign o[41666] = i[81];
  assign o[41667] = i[81];
  assign o[41668] = i[81];
  assign o[41669] = i[81];
  assign o[41670] = i[81];
  assign o[41671] = i[81];
  assign o[41672] = i[81];
  assign o[41673] = i[81];
  assign o[41674] = i[81];
  assign o[41675] = i[81];
  assign o[41676] = i[81];
  assign o[41677] = i[81];
  assign o[41678] = i[81];
  assign o[41679] = i[81];
  assign o[41680] = i[81];
  assign o[41681] = i[81];
  assign o[41682] = i[81];
  assign o[41683] = i[81];
  assign o[41684] = i[81];
  assign o[41685] = i[81];
  assign o[41686] = i[81];
  assign o[41687] = i[81];
  assign o[41688] = i[81];
  assign o[41689] = i[81];
  assign o[41690] = i[81];
  assign o[41691] = i[81];
  assign o[41692] = i[81];
  assign o[41693] = i[81];
  assign o[41694] = i[81];
  assign o[41695] = i[81];
  assign o[41696] = i[81];
  assign o[41697] = i[81];
  assign o[41698] = i[81];
  assign o[41699] = i[81];
  assign o[41700] = i[81];
  assign o[41701] = i[81];
  assign o[41702] = i[81];
  assign o[41703] = i[81];
  assign o[41704] = i[81];
  assign o[41705] = i[81];
  assign o[41706] = i[81];
  assign o[41707] = i[81];
  assign o[41708] = i[81];
  assign o[41709] = i[81];
  assign o[41710] = i[81];
  assign o[41711] = i[81];
  assign o[41712] = i[81];
  assign o[41713] = i[81];
  assign o[41714] = i[81];
  assign o[41715] = i[81];
  assign o[41716] = i[81];
  assign o[41717] = i[81];
  assign o[41718] = i[81];
  assign o[41719] = i[81];
  assign o[41720] = i[81];
  assign o[41721] = i[81];
  assign o[41722] = i[81];
  assign o[41723] = i[81];
  assign o[41724] = i[81];
  assign o[41725] = i[81];
  assign o[41726] = i[81];
  assign o[41727] = i[81];
  assign o[41728] = i[81];
  assign o[41729] = i[81];
  assign o[41730] = i[81];
  assign o[41731] = i[81];
  assign o[41732] = i[81];
  assign o[41733] = i[81];
  assign o[41734] = i[81];
  assign o[41735] = i[81];
  assign o[41736] = i[81];
  assign o[41737] = i[81];
  assign o[41738] = i[81];
  assign o[41739] = i[81];
  assign o[41740] = i[81];
  assign o[41741] = i[81];
  assign o[41742] = i[81];
  assign o[41743] = i[81];
  assign o[41744] = i[81];
  assign o[41745] = i[81];
  assign o[41746] = i[81];
  assign o[41747] = i[81];
  assign o[41748] = i[81];
  assign o[41749] = i[81];
  assign o[41750] = i[81];
  assign o[41751] = i[81];
  assign o[41752] = i[81];
  assign o[41753] = i[81];
  assign o[41754] = i[81];
  assign o[41755] = i[81];
  assign o[41756] = i[81];
  assign o[41757] = i[81];
  assign o[41758] = i[81];
  assign o[41759] = i[81];
  assign o[41760] = i[81];
  assign o[41761] = i[81];
  assign o[41762] = i[81];
  assign o[41763] = i[81];
  assign o[41764] = i[81];
  assign o[41765] = i[81];
  assign o[41766] = i[81];
  assign o[41767] = i[81];
  assign o[41768] = i[81];
  assign o[41769] = i[81];
  assign o[41770] = i[81];
  assign o[41771] = i[81];
  assign o[41772] = i[81];
  assign o[41773] = i[81];
  assign o[41774] = i[81];
  assign o[41775] = i[81];
  assign o[41776] = i[81];
  assign o[41777] = i[81];
  assign o[41778] = i[81];
  assign o[41779] = i[81];
  assign o[41780] = i[81];
  assign o[41781] = i[81];
  assign o[41782] = i[81];
  assign o[41783] = i[81];
  assign o[41784] = i[81];
  assign o[41785] = i[81];
  assign o[41786] = i[81];
  assign o[41787] = i[81];
  assign o[41788] = i[81];
  assign o[41789] = i[81];
  assign o[41790] = i[81];
  assign o[41791] = i[81];
  assign o[41792] = i[81];
  assign o[41793] = i[81];
  assign o[41794] = i[81];
  assign o[41795] = i[81];
  assign o[41796] = i[81];
  assign o[41797] = i[81];
  assign o[41798] = i[81];
  assign o[41799] = i[81];
  assign o[41800] = i[81];
  assign o[41801] = i[81];
  assign o[41802] = i[81];
  assign o[41803] = i[81];
  assign o[41804] = i[81];
  assign o[41805] = i[81];
  assign o[41806] = i[81];
  assign o[41807] = i[81];
  assign o[41808] = i[81];
  assign o[41809] = i[81];
  assign o[41810] = i[81];
  assign o[41811] = i[81];
  assign o[41812] = i[81];
  assign o[41813] = i[81];
  assign o[41814] = i[81];
  assign o[41815] = i[81];
  assign o[41816] = i[81];
  assign o[41817] = i[81];
  assign o[41818] = i[81];
  assign o[41819] = i[81];
  assign o[41820] = i[81];
  assign o[41821] = i[81];
  assign o[41822] = i[81];
  assign o[41823] = i[81];
  assign o[41824] = i[81];
  assign o[41825] = i[81];
  assign o[41826] = i[81];
  assign o[41827] = i[81];
  assign o[41828] = i[81];
  assign o[41829] = i[81];
  assign o[41830] = i[81];
  assign o[41831] = i[81];
  assign o[41832] = i[81];
  assign o[41833] = i[81];
  assign o[41834] = i[81];
  assign o[41835] = i[81];
  assign o[41836] = i[81];
  assign o[41837] = i[81];
  assign o[41838] = i[81];
  assign o[41839] = i[81];
  assign o[41840] = i[81];
  assign o[41841] = i[81];
  assign o[41842] = i[81];
  assign o[41843] = i[81];
  assign o[41844] = i[81];
  assign o[41845] = i[81];
  assign o[41846] = i[81];
  assign o[41847] = i[81];
  assign o[41848] = i[81];
  assign o[41849] = i[81];
  assign o[41850] = i[81];
  assign o[41851] = i[81];
  assign o[41852] = i[81];
  assign o[41853] = i[81];
  assign o[41854] = i[81];
  assign o[41855] = i[81];
  assign o[41856] = i[81];
  assign o[41857] = i[81];
  assign o[41858] = i[81];
  assign o[41859] = i[81];
  assign o[41860] = i[81];
  assign o[41861] = i[81];
  assign o[41862] = i[81];
  assign o[41863] = i[81];
  assign o[41864] = i[81];
  assign o[41865] = i[81];
  assign o[41866] = i[81];
  assign o[41867] = i[81];
  assign o[41868] = i[81];
  assign o[41869] = i[81];
  assign o[41870] = i[81];
  assign o[41871] = i[81];
  assign o[41872] = i[81];
  assign o[41873] = i[81];
  assign o[41874] = i[81];
  assign o[41875] = i[81];
  assign o[41876] = i[81];
  assign o[41877] = i[81];
  assign o[41878] = i[81];
  assign o[41879] = i[81];
  assign o[41880] = i[81];
  assign o[41881] = i[81];
  assign o[41882] = i[81];
  assign o[41883] = i[81];
  assign o[41884] = i[81];
  assign o[41885] = i[81];
  assign o[41886] = i[81];
  assign o[41887] = i[81];
  assign o[41888] = i[81];
  assign o[41889] = i[81];
  assign o[41890] = i[81];
  assign o[41891] = i[81];
  assign o[41892] = i[81];
  assign o[41893] = i[81];
  assign o[41894] = i[81];
  assign o[41895] = i[81];
  assign o[41896] = i[81];
  assign o[41897] = i[81];
  assign o[41898] = i[81];
  assign o[41899] = i[81];
  assign o[41900] = i[81];
  assign o[41901] = i[81];
  assign o[41902] = i[81];
  assign o[41903] = i[81];
  assign o[41904] = i[81];
  assign o[41905] = i[81];
  assign o[41906] = i[81];
  assign o[41907] = i[81];
  assign o[41908] = i[81];
  assign o[41909] = i[81];
  assign o[41910] = i[81];
  assign o[41911] = i[81];
  assign o[41912] = i[81];
  assign o[41913] = i[81];
  assign o[41914] = i[81];
  assign o[41915] = i[81];
  assign o[41916] = i[81];
  assign o[41917] = i[81];
  assign o[41918] = i[81];
  assign o[41919] = i[81];
  assign o[41920] = i[81];
  assign o[41921] = i[81];
  assign o[41922] = i[81];
  assign o[41923] = i[81];
  assign o[41924] = i[81];
  assign o[41925] = i[81];
  assign o[41926] = i[81];
  assign o[41927] = i[81];
  assign o[41928] = i[81];
  assign o[41929] = i[81];
  assign o[41930] = i[81];
  assign o[41931] = i[81];
  assign o[41932] = i[81];
  assign o[41933] = i[81];
  assign o[41934] = i[81];
  assign o[41935] = i[81];
  assign o[41936] = i[81];
  assign o[41937] = i[81];
  assign o[41938] = i[81];
  assign o[41939] = i[81];
  assign o[41940] = i[81];
  assign o[41941] = i[81];
  assign o[41942] = i[81];
  assign o[41943] = i[81];
  assign o[41944] = i[81];
  assign o[41945] = i[81];
  assign o[41946] = i[81];
  assign o[41947] = i[81];
  assign o[41948] = i[81];
  assign o[41949] = i[81];
  assign o[41950] = i[81];
  assign o[41951] = i[81];
  assign o[41952] = i[81];
  assign o[41953] = i[81];
  assign o[41954] = i[81];
  assign o[41955] = i[81];
  assign o[41956] = i[81];
  assign o[41957] = i[81];
  assign o[41958] = i[81];
  assign o[41959] = i[81];
  assign o[41960] = i[81];
  assign o[41961] = i[81];
  assign o[41962] = i[81];
  assign o[41963] = i[81];
  assign o[41964] = i[81];
  assign o[41965] = i[81];
  assign o[41966] = i[81];
  assign o[41967] = i[81];
  assign o[41968] = i[81];
  assign o[41969] = i[81];
  assign o[41970] = i[81];
  assign o[41971] = i[81];
  assign o[41972] = i[81];
  assign o[41973] = i[81];
  assign o[41974] = i[81];
  assign o[41975] = i[81];
  assign o[41976] = i[81];
  assign o[41977] = i[81];
  assign o[41978] = i[81];
  assign o[41979] = i[81];
  assign o[41980] = i[81];
  assign o[41981] = i[81];
  assign o[41982] = i[81];
  assign o[41983] = i[81];
  assign o[40960] = i[80];
  assign o[40961] = i[80];
  assign o[40962] = i[80];
  assign o[40963] = i[80];
  assign o[40964] = i[80];
  assign o[40965] = i[80];
  assign o[40966] = i[80];
  assign o[40967] = i[80];
  assign o[40968] = i[80];
  assign o[40969] = i[80];
  assign o[40970] = i[80];
  assign o[40971] = i[80];
  assign o[40972] = i[80];
  assign o[40973] = i[80];
  assign o[40974] = i[80];
  assign o[40975] = i[80];
  assign o[40976] = i[80];
  assign o[40977] = i[80];
  assign o[40978] = i[80];
  assign o[40979] = i[80];
  assign o[40980] = i[80];
  assign o[40981] = i[80];
  assign o[40982] = i[80];
  assign o[40983] = i[80];
  assign o[40984] = i[80];
  assign o[40985] = i[80];
  assign o[40986] = i[80];
  assign o[40987] = i[80];
  assign o[40988] = i[80];
  assign o[40989] = i[80];
  assign o[40990] = i[80];
  assign o[40991] = i[80];
  assign o[40992] = i[80];
  assign o[40993] = i[80];
  assign o[40994] = i[80];
  assign o[40995] = i[80];
  assign o[40996] = i[80];
  assign o[40997] = i[80];
  assign o[40998] = i[80];
  assign o[40999] = i[80];
  assign o[41000] = i[80];
  assign o[41001] = i[80];
  assign o[41002] = i[80];
  assign o[41003] = i[80];
  assign o[41004] = i[80];
  assign o[41005] = i[80];
  assign o[41006] = i[80];
  assign o[41007] = i[80];
  assign o[41008] = i[80];
  assign o[41009] = i[80];
  assign o[41010] = i[80];
  assign o[41011] = i[80];
  assign o[41012] = i[80];
  assign o[41013] = i[80];
  assign o[41014] = i[80];
  assign o[41015] = i[80];
  assign o[41016] = i[80];
  assign o[41017] = i[80];
  assign o[41018] = i[80];
  assign o[41019] = i[80];
  assign o[41020] = i[80];
  assign o[41021] = i[80];
  assign o[41022] = i[80];
  assign o[41023] = i[80];
  assign o[41024] = i[80];
  assign o[41025] = i[80];
  assign o[41026] = i[80];
  assign o[41027] = i[80];
  assign o[41028] = i[80];
  assign o[41029] = i[80];
  assign o[41030] = i[80];
  assign o[41031] = i[80];
  assign o[41032] = i[80];
  assign o[41033] = i[80];
  assign o[41034] = i[80];
  assign o[41035] = i[80];
  assign o[41036] = i[80];
  assign o[41037] = i[80];
  assign o[41038] = i[80];
  assign o[41039] = i[80];
  assign o[41040] = i[80];
  assign o[41041] = i[80];
  assign o[41042] = i[80];
  assign o[41043] = i[80];
  assign o[41044] = i[80];
  assign o[41045] = i[80];
  assign o[41046] = i[80];
  assign o[41047] = i[80];
  assign o[41048] = i[80];
  assign o[41049] = i[80];
  assign o[41050] = i[80];
  assign o[41051] = i[80];
  assign o[41052] = i[80];
  assign o[41053] = i[80];
  assign o[41054] = i[80];
  assign o[41055] = i[80];
  assign o[41056] = i[80];
  assign o[41057] = i[80];
  assign o[41058] = i[80];
  assign o[41059] = i[80];
  assign o[41060] = i[80];
  assign o[41061] = i[80];
  assign o[41062] = i[80];
  assign o[41063] = i[80];
  assign o[41064] = i[80];
  assign o[41065] = i[80];
  assign o[41066] = i[80];
  assign o[41067] = i[80];
  assign o[41068] = i[80];
  assign o[41069] = i[80];
  assign o[41070] = i[80];
  assign o[41071] = i[80];
  assign o[41072] = i[80];
  assign o[41073] = i[80];
  assign o[41074] = i[80];
  assign o[41075] = i[80];
  assign o[41076] = i[80];
  assign o[41077] = i[80];
  assign o[41078] = i[80];
  assign o[41079] = i[80];
  assign o[41080] = i[80];
  assign o[41081] = i[80];
  assign o[41082] = i[80];
  assign o[41083] = i[80];
  assign o[41084] = i[80];
  assign o[41085] = i[80];
  assign o[41086] = i[80];
  assign o[41087] = i[80];
  assign o[41088] = i[80];
  assign o[41089] = i[80];
  assign o[41090] = i[80];
  assign o[41091] = i[80];
  assign o[41092] = i[80];
  assign o[41093] = i[80];
  assign o[41094] = i[80];
  assign o[41095] = i[80];
  assign o[41096] = i[80];
  assign o[41097] = i[80];
  assign o[41098] = i[80];
  assign o[41099] = i[80];
  assign o[41100] = i[80];
  assign o[41101] = i[80];
  assign o[41102] = i[80];
  assign o[41103] = i[80];
  assign o[41104] = i[80];
  assign o[41105] = i[80];
  assign o[41106] = i[80];
  assign o[41107] = i[80];
  assign o[41108] = i[80];
  assign o[41109] = i[80];
  assign o[41110] = i[80];
  assign o[41111] = i[80];
  assign o[41112] = i[80];
  assign o[41113] = i[80];
  assign o[41114] = i[80];
  assign o[41115] = i[80];
  assign o[41116] = i[80];
  assign o[41117] = i[80];
  assign o[41118] = i[80];
  assign o[41119] = i[80];
  assign o[41120] = i[80];
  assign o[41121] = i[80];
  assign o[41122] = i[80];
  assign o[41123] = i[80];
  assign o[41124] = i[80];
  assign o[41125] = i[80];
  assign o[41126] = i[80];
  assign o[41127] = i[80];
  assign o[41128] = i[80];
  assign o[41129] = i[80];
  assign o[41130] = i[80];
  assign o[41131] = i[80];
  assign o[41132] = i[80];
  assign o[41133] = i[80];
  assign o[41134] = i[80];
  assign o[41135] = i[80];
  assign o[41136] = i[80];
  assign o[41137] = i[80];
  assign o[41138] = i[80];
  assign o[41139] = i[80];
  assign o[41140] = i[80];
  assign o[41141] = i[80];
  assign o[41142] = i[80];
  assign o[41143] = i[80];
  assign o[41144] = i[80];
  assign o[41145] = i[80];
  assign o[41146] = i[80];
  assign o[41147] = i[80];
  assign o[41148] = i[80];
  assign o[41149] = i[80];
  assign o[41150] = i[80];
  assign o[41151] = i[80];
  assign o[41152] = i[80];
  assign o[41153] = i[80];
  assign o[41154] = i[80];
  assign o[41155] = i[80];
  assign o[41156] = i[80];
  assign o[41157] = i[80];
  assign o[41158] = i[80];
  assign o[41159] = i[80];
  assign o[41160] = i[80];
  assign o[41161] = i[80];
  assign o[41162] = i[80];
  assign o[41163] = i[80];
  assign o[41164] = i[80];
  assign o[41165] = i[80];
  assign o[41166] = i[80];
  assign o[41167] = i[80];
  assign o[41168] = i[80];
  assign o[41169] = i[80];
  assign o[41170] = i[80];
  assign o[41171] = i[80];
  assign o[41172] = i[80];
  assign o[41173] = i[80];
  assign o[41174] = i[80];
  assign o[41175] = i[80];
  assign o[41176] = i[80];
  assign o[41177] = i[80];
  assign o[41178] = i[80];
  assign o[41179] = i[80];
  assign o[41180] = i[80];
  assign o[41181] = i[80];
  assign o[41182] = i[80];
  assign o[41183] = i[80];
  assign o[41184] = i[80];
  assign o[41185] = i[80];
  assign o[41186] = i[80];
  assign o[41187] = i[80];
  assign o[41188] = i[80];
  assign o[41189] = i[80];
  assign o[41190] = i[80];
  assign o[41191] = i[80];
  assign o[41192] = i[80];
  assign o[41193] = i[80];
  assign o[41194] = i[80];
  assign o[41195] = i[80];
  assign o[41196] = i[80];
  assign o[41197] = i[80];
  assign o[41198] = i[80];
  assign o[41199] = i[80];
  assign o[41200] = i[80];
  assign o[41201] = i[80];
  assign o[41202] = i[80];
  assign o[41203] = i[80];
  assign o[41204] = i[80];
  assign o[41205] = i[80];
  assign o[41206] = i[80];
  assign o[41207] = i[80];
  assign o[41208] = i[80];
  assign o[41209] = i[80];
  assign o[41210] = i[80];
  assign o[41211] = i[80];
  assign o[41212] = i[80];
  assign o[41213] = i[80];
  assign o[41214] = i[80];
  assign o[41215] = i[80];
  assign o[41216] = i[80];
  assign o[41217] = i[80];
  assign o[41218] = i[80];
  assign o[41219] = i[80];
  assign o[41220] = i[80];
  assign o[41221] = i[80];
  assign o[41222] = i[80];
  assign o[41223] = i[80];
  assign o[41224] = i[80];
  assign o[41225] = i[80];
  assign o[41226] = i[80];
  assign o[41227] = i[80];
  assign o[41228] = i[80];
  assign o[41229] = i[80];
  assign o[41230] = i[80];
  assign o[41231] = i[80];
  assign o[41232] = i[80];
  assign o[41233] = i[80];
  assign o[41234] = i[80];
  assign o[41235] = i[80];
  assign o[41236] = i[80];
  assign o[41237] = i[80];
  assign o[41238] = i[80];
  assign o[41239] = i[80];
  assign o[41240] = i[80];
  assign o[41241] = i[80];
  assign o[41242] = i[80];
  assign o[41243] = i[80];
  assign o[41244] = i[80];
  assign o[41245] = i[80];
  assign o[41246] = i[80];
  assign o[41247] = i[80];
  assign o[41248] = i[80];
  assign o[41249] = i[80];
  assign o[41250] = i[80];
  assign o[41251] = i[80];
  assign o[41252] = i[80];
  assign o[41253] = i[80];
  assign o[41254] = i[80];
  assign o[41255] = i[80];
  assign o[41256] = i[80];
  assign o[41257] = i[80];
  assign o[41258] = i[80];
  assign o[41259] = i[80];
  assign o[41260] = i[80];
  assign o[41261] = i[80];
  assign o[41262] = i[80];
  assign o[41263] = i[80];
  assign o[41264] = i[80];
  assign o[41265] = i[80];
  assign o[41266] = i[80];
  assign o[41267] = i[80];
  assign o[41268] = i[80];
  assign o[41269] = i[80];
  assign o[41270] = i[80];
  assign o[41271] = i[80];
  assign o[41272] = i[80];
  assign o[41273] = i[80];
  assign o[41274] = i[80];
  assign o[41275] = i[80];
  assign o[41276] = i[80];
  assign o[41277] = i[80];
  assign o[41278] = i[80];
  assign o[41279] = i[80];
  assign o[41280] = i[80];
  assign o[41281] = i[80];
  assign o[41282] = i[80];
  assign o[41283] = i[80];
  assign o[41284] = i[80];
  assign o[41285] = i[80];
  assign o[41286] = i[80];
  assign o[41287] = i[80];
  assign o[41288] = i[80];
  assign o[41289] = i[80];
  assign o[41290] = i[80];
  assign o[41291] = i[80];
  assign o[41292] = i[80];
  assign o[41293] = i[80];
  assign o[41294] = i[80];
  assign o[41295] = i[80];
  assign o[41296] = i[80];
  assign o[41297] = i[80];
  assign o[41298] = i[80];
  assign o[41299] = i[80];
  assign o[41300] = i[80];
  assign o[41301] = i[80];
  assign o[41302] = i[80];
  assign o[41303] = i[80];
  assign o[41304] = i[80];
  assign o[41305] = i[80];
  assign o[41306] = i[80];
  assign o[41307] = i[80];
  assign o[41308] = i[80];
  assign o[41309] = i[80];
  assign o[41310] = i[80];
  assign o[41311] = i[80];
  assign o[41312] = i[80];
  assign o[41313] = i[80];
  assign o[41314] = i[80];
  assign o[41315] = i[80];
  assign o[41316] = i[80];
  assign o[41317] = i[80];
  assign o[41318] = i[80];
  assign o[41319] = i[80];
  assign o[41320] = i[80];
  assign o[41321] = i[80];
  assign o[41322] = i[80];
  assign o[41323] = i[80];
  assign o[41324] = i[80];
  assign o[41325] = i[80];
  assign o[41326] = i[80];
  assign o[41327] = i[80];
  assign o[41328] = i[80];
  assign o[41329] = i[80];
  assign o[41330] = i[80];
  assign o[41331] = i[80];
  assign o[41332] = i[80];
  assign o[41333] = i[80];
  assign o[41334] = i[80];
  assign o[41335] = i[80];
  assign o[41336] = i[80];
  assign o[41337] = i[80];
  assign o[41338] = i[80];
  assign o[41339] = i[80];
  assign o[41340] = i[80];
  assign o[41341] = i[80];
  assign o[41342] = i[80];
  assign o[41343] = i[80];
  assign o[41344] = i[80];
  assign o[41345] = i[80];
  assign o[41346] = i[80];
  assign o[41347] = i[80];
  assign o[41348] = i[80];
  assign o[41349] = i[80];
  assign o[41350] = i[80];
  assign o[41351] = i[80];
  assign o[41352] = i[80];
  assign o[41353] = i[80];
  assign o[41354] = i[80];
  assign o[41355] = i[80];
  assign o[41356] = i[80];
  assign o[41357] = i[80];
  assign o[41358] = i[80];
  assign o[41359] = i[80];
  assign o[41360] = i[80];
  assign o[41361] = i[80];
  assign o[41362] = i[80];
  assign o[41363] = i[80];
  assign o[41364] = i[80];
  assign o[41365] = i[80];
  assign o[41366] = i[80];
  assign o[41367] = i[80];
  assign o[41368] = i[80];
  assign o[41369] = i[80];
  assign o[41370] = i[80];
  assign o[41371] = i[80];
  assign o[41372] = i[80];
  assign o[41373] = i[80];
  assign o[41374] = i[80];
  assign o[41375] = i[80];
  assign o[41376] = i[80];
  assign o[41377] = i[80];
  assign o[41378] = i[80];
  assign o[41379] = i[80];
  assign o[41380] = i[80];
  assign o[41381] = i[80];
  assign o[41382] = i[80];
  assign o[41383] = i[80];
  assign o[41384] = i[80];
  assign o[41385] = i[80];
  assign o[41386] = i[80];
  assign o[41387] = i[80];
  assign o[41388] = i[80];
  assign o[41389] = i[80];
  assign o[41390] = i[80];
  assign o[41391] = i[80];
  assign o[41392] = i[80];
  assign o[41393] = i[80];
  assign o[41394] = i[80];
  assign o[41395] = i[80];
  assign o[41396] = i[80];
  assign o[41397] = i[80];
  assign o[41398] = i[80];
  assign o[41399] = i[80];
  assign o[41400] = i[80];
  assign o[41401] = i[80];
  assign o[41402] = i[80];
  assign o[41403] = i[80];
  assign o[41404] = i[80];
  assign o[41405] = i[80];
  assign o[41406] = i[80];
  assign o[41407] = i[80];
  assign o[41408] = i[80];
  assign o[41409] = i[80];
  assign o[41410] = i[80];
  assign o[41411] = i[80];
  assign o[41412] = i[80];
  assign o[41413] = i[80];
  assign o[41414] = i[80];
  assign o[41415] = i[80];
  assign o[41416] = i[80];
  assign o[41417] = i[80];
  assign o[41418] = i[80];
  assign o[41419] = i[80];
  assign o[41420] = i[80];
  assign o[41421] = i[80];
  assign o[41422] = i[80];
  assign o[41423] = i[80];
  assign o[41424] = i[80];
  assign o[41425] = i[80];
  assign o[41426] = i[80];
  assign o[41427] = i[80];
  assign o[41428] = i[80];
  assign o[41429] = i[80];
  assign o[41430] = i[80];
  assign o[41431] = i[80];
  assign o[41432] = i[80];
  assign o[41433] = i[80];
  assign o[41434] = i[80];
  assign o[41435] = i[80];
  assign o[41436] = i[80];
  assign o[41437] = i[80];
  assign o[41438] = i[80];
  assign o[41439] = i[80];
  assign o[41440] = i[80];
  assign o[41441] = i[80];
  assign o[41442] = i[80];
  assign o[41443] = i[80];
  assign o[41444] = i[80];
  assign o[41445] = i[80];
  assign o[41446] = i[80];
  assign o[41447] = i[80];
  assign o[41448] = i[80];
  assign o[41449] = i[80];
  assign o[41450] = i[80];
  assign o[41451] = i[80];
  assign o[41452] = i[80];
  assign o[41453] = i[80];
  assign o[41454] = i[80];
  assign o[41455] = i[80];
  assign o[41456] = i[80];
  assign o[41457] = i[80];
  assign o[41458] = i[80];
  assign o[41459] = i[80];
  assign o[41460] = i[80];
  assign o[41461] = i[80];
  assign o[41462] = i[80];
  assign o[41463] = i[80];
  assign o[41464] = i[80];
  assign o[41465] = i[80];
  assign o[41466] = i[80];
  assign o[41467] = i[80];
  assign o[41468] = i[80];
  assign o[41469] = i[80];
  assign o[41470] = i[80];
  assign o[41471] = i[80];
  assign o[40448] = i[79];
  assign o[40449] = i[79];
  assign o[40450] = i[79];
  assign o[40451] = i[79];
  assign o[40452] = i[79];
  assign o[40453] = i[79];
  assign o[40454] = i[79];
  assign o[40455] = i[79];
  assign o[40456] = i[79];
  assign o[40457] = i[79];
  assign o[40458] = i[79];
  assign o[40459] = i[79];
  assign o[40460] = i[79];
  assign o[40461] = i[79];
  assign o[40462] = i[79];
  assign o[40463] = i[79];
  assign o[40464] = i[79];
  assign o[40465] = i[79];
  assign o[40466] = i[79];
  assign o[40467] = i[79];
  assign o[40468] = i[79];
  assign o[40469] = i[79];
  assign o[40470] = i[79];
  assign o[40471] = i[79];
  assign o[40472] = i[79];
  assign o[40473] = i[79];
  assign o[40474] = i[79];
  assign o[40475] = i[79];
  assign o[40476] = i[79];
  assign o[40477] = i[79];
  assign o[40478] = i[79];
  assign o[40479] = i[79];
  assign o[40480] = i[79];
  assign o[40481] = i[79];
  assign o[40482] = i[79];
  assign o[40483] = i[79];
  assign o[40484] = i[79];
  assign o[40485] = i[79];
  assign o[40486] = i[79];
  assign o[40487] = i[79];
  assign o[40488] = i[79];
  assign o[40489] = i[79];
  assign o[40490] = i[79];
  assign o[40491] = i[79];
  assign o[40492] = i[79];
  assign o[40493] = i[79];
  assign o[40494] = i[79];
  assign o[40495] = i[79];
  assign o[40496] = i[79];
  assign o[40497] = i[79];
  assign o[40498] = i[79];
  assign o[40499] = i[79];
  assign o[40500] = i[79];
  assign o[40501] = i[79];
  assign o[40502] = i[79];
  assign o[40503] = i[79];
  assign o[40504] = i[79];
  assign o[40505] = i[79];
  assign o[40506] = i[79];
  assign o[40507] = i[79];
  assign o[40508] = i[79];
  assign o[40509] = i[79];
  assign o[40510] = i[79];
  assign o[40511] = i[79];
  assign o[40512] = i[79];
  assign o[40513] = i[79];
  assign o[40514] = i[79];
  assign o[40515] = i[79];
  assign o[40516] = i[79];
  assign o[40517] = i[79];
  assign o[40518] = i[79];
  assign o[40519] = i[79];
  assign o[40520] = i[79];
  assign o[40521] = i[79];
  assign o[40522] = i[79];
  assign o[40523] = i[79];
  assign o[40524] = i[79];
  assign o[40525] = i[79];
  assign o[40526] = i[79];
  assign o[40527] = i[79];
  assign o[40528] = i[79];
  assign o[40529] = i[79];
  assign o[40530] = i[79];
  assign o[40531] = i[79];
  assign o[40532] = i[79];
  assign o[40533] = i[79];
  assign o[40534] = i[79];
  assign o[40535] = i[79];
  assign o[40536] = i[79];
  assign o[40537] = i[79];
  assign o[40538] = i[79];
  assign o[40539] = i[79];
  assign o[40540] = i[79];
  assign o[40541] = i[79];
  assign o[40542] = i[79];
  assign o[40543] = i[79];
  assign o[40544] = i[79];
  assign o[40545] = i[79];
  assign o[40546] = i[79];
  assign o[40547] = i[79];
  assign o[40548] = i[79];
  assign o[40549] = i[79];
  assign o[40550] = i[79];
  assign o[40551] = i[79];
  assign o[40552] = i[79];
  assign o[40553] = i[79];
  assign o[40554] = i[79];
  assign o[40555] = i[79];
  assign o[40556] = i[79];
  assign o[40557] = i[79];
  assign o[40558] = i[79];
  assign o[40559] = i[79];
  assign o[40560] = i[79];
  assign o[40561] = i[79];
  assign o[40562] = i[79];
  assign o[40563] = i[79];
  assign o[40564] = i[79];
  assign o[40565] = i[79];
  assign o[40566] = i[79];
  assign o[40567] = i[79];
  assign o[40568] = i[79];
  assign o[40569] = i[79];
  assign o[40570] = i[79];
  assign o[40571] = i[79];
  assign o[40572] = i[79];
  assign o[40573] = i[79];
  assign o[40574] = i[79];
  assign o[40575] = i[79];
  assign o[40576] = i[79];
  assign o[40577] = i[79];
  assign o[40578] = i[79];
  assign o[40579] = i[79];
  assign o[40580] = i[79];
  assign o[40581] = i[79];
  assign o[40582] = i[79];
  assign o[40583] = i[79];
  assign o[40584] = i[79];
  assign o[40585] = i[79];
  assign o[40586] = i[79];
  assign o[40587] = i[79];
  assign o[40588] = i[79];
  assign o[40589] = i[79];
  assign o[40590] = i[79];
  assign o[40591] = i[79];
  assign o[40592] = i[79];
  assign o[40593] = i[79];
  assign o[40594] = i[79];
  assign o[40595] = i[79];
  assign o[40596] = i[79];
  assign o[40597] = i[79];
  assign o[40598] = i[79];
  assign o[40599] = i[79];
  assign o[40600] = i[79];
  assign o[40601] = i[79];
  assign o[40602] = i[79];
  assign o[40603] = i[79];
  assign o[40604] = i[79];
  assign o[40605] = i[79];
  assign o[40606] = i[79];
  assign o[40607] = i[79];
  assign o[40608] = i[79];
  assign o[40609] = i[79];
  assign o[40610] = i[79];
  assign o[40611] = i[79];
  assign o[40612] = i[79];
  assign o[40613] = i[79];
  assign o[40614] = i[79];
  assign o[40615] = i[79];
  assign o[40616] = i[79];
  assign o[40617] = i[79];
  assign o[40618] = i[79];
  assign o[40619] = i[79];
  assign o[40620] = i[79];
  assign o[40621] = i[79];
  assign o[40622] = i[79];
  assign o[40623] = i[79];
  assign o[40624] = i[79];
  assign o[40625] = i[79];
  assign o[40626] = i[79];
  assign o[40627] = i[79];
  assign o[40628] = i[79];
  assign o[40629] = i[79];
  assign o[40630] = i[79];
  assign o[40631] = i[79];
  assign o[40632] = i[79];
  assign o[40633] = i[79];
  assign o[40634] = i[79];
  assign o[40635] = i[79];
  assign o[40636] = i[79];
  assign o[40637] = i[79];
  assign o[40638] = i[79];
  assign o[40639] = i[79];
  assign o[40640] = i[79];
  assign o[40641] = i[79];
  assign o[40642] = i[79];
  assign o[40643] = i[79];
  assign o[40644] = i[79];
  assign o[40645] = i[79];
  assign o[40646] = i[79];
  assign o[40647] = i[79];
  assign o[40648] = i[79];
  assign o[40649] = i[79];
  assign o[40650] = i[79];
  assign o[40651] = i[79];
  assign o[40652] = i[79];
  assign o[40653] = i[79];
  assign o[40654] = i[79];
  assign o[40655] = i[79];
  assign o[40656] = i[79];
  assign o[40657] = i[79];
  assign o[40658] = i[79];
  assign o[40659] = i[79];
  assign o[40660] = i[79];
  assign o[40661] = i[79];
  assign o[40662] = i[79];
  assign o[40663] = i[79];
  assign o[40664] = i[79];
  assign o[40665] = i[79];
  assign o[40666] = i[79];
  assign o[40667] = i[79];
  assign o[40668] = i[79];
  assign o[40669] = i[79];
  assign o[40670] = i[79];
  assign o[40671] = i[79];
  assign o[40672] = i[79];
  assign o[40673] = i[79];
  assign o[40674] = i[79];
  assign o[40675] = i[79];
  assign o[40676] = i[79];
  assign o[40677] = i[79];
  assign o[40678] = i[79];
  assign o[40679] = i[79];
  assign o[40680] = i[79];
  assign o[40681] = i[79];
  assign o[40682] = i[79];
  assign o[40683] = i[79];
  assign o[40684] = i[79];
  assign o[40685] = i[79];
  assign o[40686] = i[79];
  assign o[40687] = i[79];
  assign o[40688] = i[79];
  assign o[40689] = i[79];
  assign o[40690] = i[79];
  assign o[40691] = i[79];
  assign o[40692] = i[79];
  assign o[40693] = i[79];
  assign o[40694] = i[79];
  assign o[40695] = i[79];
  assign o[40696] = i[79];
  assign o[40697] = i[79];
  assign o[40698] = i[79];
  assign o[40699] = i[79];
  assign o[40700] = i[79];
  assign o[40701] = i[79];
  assign o[40702] = i[79];
  assign o[40703] = i[79];
  assign o[40704] = i[79];
  assign o[40705] = i[79];
  assign o[40706] = i[79];
  assign o[40707] = i[79];
  assign o[40708] = i[79];
  assign o[40709] = i[79];
  assign o[40710] = i[79];
  assign o[40711] = i[79];
  assign o[40712] = i[79];
  assign o[40713] = i[79];
  assign o[40714] = i[79];
  assign o[40715] = i[79];
  assign o[40716] = i[79];
  assign o[40717] = i[79];
  assign o[40718] = i[79];
  assign o[40719] = i[79];
  assign o[40720] = i[79];
  assign o[40721] = i[79];
  assign o[40722] = i[79];
  assign o[40723] = i[79];
  assign o[40724] = i[79];
  assign o[40725] = i[79];
  assign o[40726] = i[79];
  assign o[40727] = i[79];
  assign o[40728] = i[79];
  assign o[40729] = i[79];
  assign o[40730] = i[79];
  assign o[40731] = i[79];
  assign o[40732] = i[79];
  assign o[40733] = i[79];
  assign o[40734] = i[79];
  assign o[40735] = i[79];
  assign o[40736] = i[79];
  assign o[40737] = i[79];
  assign o[40738] = i[79];
  assign o[40739] = i[79];
  assign o[40740] = i[79];
  assign o[40741] = i[79];
  assign o[40742] = i[79];
  assign o[40743] = i[79];
  assign o[40744] = i[79];
  assign o[40745] = i[79];
  assign o[40746] = i[79];
  assign o[40747] = i[79];
  assign o[40748] = i[79];
  assign o[40749] = i[79];
  assign o[40750] = i[79];
  assign o[40751] = i[79];
  assign o[40752] = i[79];
  assign o[40753] = i[79];
  assign o[40754] = i[79];
  assign o[40755] = i[79];
  assign o[40756] = i[79];
  assign o[40757] = i[79];
  assign o[40758] = i[79];
  assign o[40759] = i[79];
  assign o[40760] = i[79];
  assign o[40761] = i[79];
  assign o[40762] = i[79];
  assign o[40763] = i[79];
  assign o[40764] = i[79];
  assign o[40765] = i[79];
  assign o[40766] = i[79];
  assign o[40767] = i[79];
  assign o[40768] = i[79];
  assign o[40769] = i[79];
  assign o[40770] = i[79];
  assign o[40771] = i[79];
  assign o[40772] = i[79];
  assign o[40773] = i[79];
  assign o[40774] = i[79];
  assign o[40775] = i[79];
  assign o[40776] = i[79];
  assign o[40777] = i[79];
  assign o[40778] = i[79];
  assign o[40779] = i[79];
  assign o[40780] = i[79];
  assign o[40781] = i[79];
  assign o[40782] = i[79];
  assign o[40783] = i[79];
  assign o[40784] = i[79];
  assign o[40785] = i[79];
  assign o[40786] = i[79];
  assign o[40787] = i[79];
  assign o[40788] = i[79];
  assign o[40789] = i[79];
  assign o[40790] = i[79];
  assign o[40791] = i[79];
  assign o[40792] = i[79];
  assign o[40793] = i[79];
  assign o[40794] = i[79];
  assign o[40795] = i[79];
  assign o[40796] = i[79];
  assign o[40797] = i[79];
  assign o[40798] = i[79];
  assign o[40799] = i[79];
  assign o[40800] = i[79];
  assign o[40801] = i[79];
  assign o[40802] = i[79];
  assign o[40803] = i[79];
  assign o[40804] = i[79];
  assign o[40805] = i[79];
  assign o[40806] = i[79];
  assign o[40807] = i[79];
  assign o[40808] = i[79];
  assign o[40809] = i[79];
  assign o[40810] = i[79];
  assign o[40811] = i[79];
  assign o[40812] = i[79];
  assign o[40813] = i[79];
  assign o[40814] = i[79];
  assign o[40815] = i[79];
  assign o[40816] = i[79];
  assign o[40817] = i[79];
  assign o[40818] = i[79];
  assign o[40819] = i[79];
  assign o[40820] = i[79];
  assign o[40821] = i[79];
  assign o[40822] = i[79];
  assign o[40823] = i[79];
  assign o[40824] = i[79];
  assign o[40825] = i[79];
  assign o[40826] = i[79];
  assign o[40827] = i[79];
  assign o[40828] = i[79];
  assign o[40829] = i[79];
  assign o[40830] = i[79];
  assign o[40831] = i[79];
  assign o[40832] = i[79];
  assign o[40833] = i[79];
  assign o[40834] = i[79];
  assign o[40835] = i[79];
  assign o[40836] = i[79];
  assign o[40837] = i[79];
  assign o[40838] = i[79];
  assign o[40839] = i[79];
  assign o[40840] = i[79];
  assign o[40841] = i[79];
  assign o[40842] = i[79];
  assign o[40843] = i[79];
  assign o[40844] = i[79];
  assign o[40845] = i[79];
  assign o[40846] = i[79];
  assign o[40847] = i[79];
  assign o[40848] = i[79];
  assign o[40849] = i[79];
  assign o[40850] = i[79];
  assign o[40851] = i[79];
  assign o[40852] = i[79];
  assign o[40853] = i[79];
  assign o[40854] = i[79];
  assign o[40855] = i[79];
  assign o[40856] = i[79];
  assign o[40857] = i[79];
  assign o[40858] = i[79];
  assign o[40859] = i[79];
  assign o[40860] = i[79];
  assign o[40861] = i[79];
  assign o[40862] = i[79];
  assign o[40863] = i[79];
  assign o[40864] = i[79];
  assign o[40865] = i[79];
  assign o[40866] = i[79];
  assign o[40867] = i[79];
  assign o[40868] = i[79];
  assign o[40869] = i[79];
  assign o[40870] = i[79];
  assign o[40871] = i[79];
  assign o[40872] = i[79];
  assign o[40873] = i[79];
  assign o[40874] = i[79];
  assign o[40875] = i[79];
  assign o[40876] = i[79];
  assign o[40877] = i[79];
  assign o[40878] = i[79];
  assign o[40879] = i[79];
  assign o[40880] = i[79];
  assign o[40881] = i[79];
  assign o[40882] = i[79];
  assign o[40883] = i[79];
  assign o[40884] = i[79];
  assign o[40885] = i[79];
  assign o[40886] = i[79];
  assign o[40887] = i[79];
  assign o[40888] = i[79];
  assign o[40889] = i[79];
  assign o[40890] = i[79];
  assign o[40891] = i[79];
  assign o[40892] = i[79];
  assign o[40893] = i[79];
  assign o[40894] = i[79];
  assign o[40895] = i[79];
  assign o[40896] = i[79];
  assign o[40897] = i[79];
  assign o[40898] = i[79];
  assign o[40899] = i[79];
  assign o[40900] = i[79];
  assign o[40901] = i[79];
  assign o[40902] = i[79];
  assign o[40903] = i[79];
  assign o[40904] = i[79];
  assign o[40905] = i[79];
  assign o[40906] = i[79];
  assign o[40907] = i[79];
  assign o[40908] = i[79];
  assign o[40909] = i[79];
  assign o[40910] = i[79];
  assign o[40911] = i[79];
  assign o[40912] = i[79];
  assign o[40913] = i[79];
  assign o[40914] = i[79];
  assign o[40915] = i[79];
  assign o[40916] = i[79];
  assign o[40917] = i[79];
  assign o[40918] = i[79];
  assign o[40919] = i[79];
  assign o[40920] = i[79];
  assign o[40921] = i[79];
  assign o[40922] = i[79];
  assign o[40923] = i[79];
  assign o[40924] = i[79];
  assign o[40925] = i[79];
  assign o[40926] = i[79];
  assign o[40927] = i[79];
  assign o[40928] = i[79];
  assign o[40929] = i[79];
  assign o[40930] = i[79];
  assign o[40931] = i[79];
  assign o[40932] = i[79];
  assign o[40933] = i[79];
  assign o[40934] = i[79];
  assign o[40935] = i[79];
  assign o[40936] = i[79];
  assign o[40937] = i[79];
  assign o[40938] = i[79];
  assign o[40939] = i[79];
  assign o[40940] = i[79];
  assign o[40941] = i[79];
  assign o[40942] = i[79];
  assign o[40943] = i[79];
  assign o[40944] = i[79];
  assign o[40945] = i[79];
  assign o[40946] = i[79];
  assign o[40947] = i[79];
  assign o[40948] = i[79];
  assign o[40949] = i[79];
  assign o[40950] = i[79];
  assign o[40951] = i[79];
  assign o[40952] = i[79];
  assign o[40953] = i[79];
  assign o[40954] = i[79];
  assign o[40955] = i[79];
  assign o[40956] = i[79];
  assign o[40957] = i[79];
  assign o[40958] = i[79];
  assign o[40959] = i[79];
  assign o[39936] = i[78];
  assign o[39937] = i[78];
  assign o[39938] = i[78];
  assign o[39939] = i[78];
  assign o[39940] = i[78];
  assign o[39941] = i[78];
  assign o[39942] = i[78];
  assign o[39943] = i[78];
  assign o[39944] = i[78];
  assign o[39945] = i[78];
  assign o[39946] = i[78];
  assign o[39947] = i[78];
  assign o[39948] = i[78];
  assign o[39949] = i[78];
  assign o[39950] = i[78];
  assign o[39951] = i[78];
  assign o[39952] = i[78];
  assign o[39953] = i[78];
  assign o[39954] = i[78];
  assign o[39955] = i[78];
  assign o[39956] = i[78];
  assign o[39957] = i[78];
  assign o[39958] = i[78];
  assign o[39959] = i[78];
  assign o[39960] = i[78];
  assign o[39961] = i[78];
  assign o[39962] = i[78];
  assign o[39963] = i[78];
  assign o[39964] = i[78];
  assign o[39965] = i[78];
  assign o[39966] = i[78];
  assign o[39967] = i[78];
  assign o[39968] = i[78];
  assign o[39969] = i[78];
  assign o[39970] = i[78];
  assign o[39971] = i[78];
  assign o[39972] = i[78];
  assign o[39973] = i[78];
  assign o[39974] = i[78];
  assign o[39975] = i[78];
  assign o[39976] = i[78];
  assign o[39977] = i[78];
  assign o[39978] = i[78];
  assign o[39979] = i[78];
  assign o[39980] = i[78];
  assign o[39981] = i[78];
  assign o[39982] = i[78];
  assign o[39983] = i[78];
  assign o[39984] = i[78];
  assign o[39985] = i[78];
  assign o[39986] = i[78];
  assign o[39987] = i[78];
  assign o[39988] = i[78];
  assign o[39989] = i[78];
  assign o[39990] = i[78];
  assign o[39991] = i[78];
  assign o[39992] = i[78];
  assign o[39993] = i[78];
  assign o[39994] = i[78];
  assign o[39995] = i[78];
  assign o[39996] = i[78];
  assign o[39997] = i[78];
  assign o[39998] = i[78];
  assign o[39999] = i[78];
  assign o[40000] = i[78];
  assign o[40001] = i[78];
  assign o[40002] = i[78];
  assign o[40003] = i[78];
  assign o[40004] = i[78];
  assign o[40005] = i[78];
  assign o[40006] = i[78];
  assign o[40007] = i[78];
  assign o[40008] = i[78];
  assign o[40009] = i[78];
  assign o[40010] = i[78];
  assign o[40011] = i[78];
  assign o[40012] = i[78];
  assign o[40013] = i[78];
  assign o[40014] = i[78];
  assign o[40015] = i[78];
  assign o[40016] = i[78];
  assign o[40017] = i[78];
  assign o[40018] = i[78];
  assign o[40019] = i[78];
  assign o[40020] = i[78];
  assign o[40021] = i[78];
  assign o[40022] = i[78];
  assign o[40023] = i[78];
  assign o[40024] = i[78];
  assign o[40025] = i[78];
  assign o[40026] = i[78];
  assign o[40027] = i[78];
  assign o[40028] = i[78];
  assign o[40029] = i[78];
  assign o[40030] = i[78];
  assign o[40031] = i[78];
  assign o[40032] = i[78];
  assign o[40033] = i[78];
  assign o[40034] = i[78];
  assign o[40035] = i[78];
  assign o[40036] = i[78];
  assign o[40037] = i[78];
  assign o[40038] = i[78];
  assign o[40039] = i[78];
  assign o[40040] = i[78];
  assign o[40041] = i[78];
  assign o[40042] = i[78];
  assign o[40043] = i[78];
  assign o[40044] = i[78];
  assign o[40045] = i[78];
  assign o[40046] = i[78];
  assign o[40047] = i[78];
  assign o[40048] = i[78];
  assign o[40049] = i[78];
  assign o[40050] = i[78];
  assign o[40051] = i[78];
  assign o[40052] = i[78];
  assign o[40053] = i[78];
  assign o[40054] = i[78];
  assign o[40055] = i[78];
  assign o[40056] = i[78];
  assign o[40057] = i[78];
  assign o[40058] = i[78];
  assign o[40059] = i[78];
  assign o[40060] = i[78];
  assign o[40061] = i[78];
  assign o[40062] = i[78];
  assign o[40063] = i[78];
  assign o[40064] = i[78];
  assign o[40065] = i[78];
  assign o[40066] = i[78];
  assign o[40067] = i[78];
  assign o[40068] = i[78];
  assign o[40069] = i[78];
  assign o[40070] = i[78];
  assign o[40071] = i[78];
  assign o[40072] = i[78];
  assign o[40073] = i[78];
  assign o[40074] = i[78];
  assign o[40075] = i[78];
  assign o[40076] = i[78];
  assign o[40077] = i[78];
  assign o[40078] = i[78];
  assign o[40079] = i[78];
  assign o[40080] = i[78];
  assign o[40081] = i[78];
  assign o[40082] = i[78];
  assign o[40083] = i[78];
  assign o[40084] = i[78];
  assign o[40085] = i[78];
  assign o[40086] = i[78];
  assign o[40087] = i[78];
  assign o[40088] = i[78];
  assign o[40089] = i[78];
  assign o[40090] = i[78];
  assign o[40091] = i[78];
  assign o[40092] = i[78];
  assign o[40093] = i[78];
  assign o[40094] = i[78];
  assign o[40095] = i[78];
  assign o[40096] = i[78];
  assign o[40097] = i[78];
  assign o[40098] = i[78];
  assign o[40099] = i[78];
  assign o[40100] = i[78];
  assign o[40101] = i[78];
  assign o[40102] = i[78];
  assign o[40103] = i[78];
  assign o[40104] = i[78];
  assign o[40105] = i[78];
  assign o[40106] = i[78];
  assign o[40107] = i[78];
  assign o[40108] = i[78];
  assign o[40109] = i[78];
  assign o[40110] = i[78];
  assign o[40111] = i[78];
  assign o[40112] = i[78];
  assign o[40113] = i[78];
  assign o[40114] = i[78];
  assign o[40115] = i[78];
  assign o[40116] = i[78];
  assign o[40117] = i[78];
  assign o[40118] = i[78];
  assign o[40119] = i[78];
  assign o[40120] = i[78];
  assign o[40121] = i[78];
  assign o[40122] = i[78];
  assign o[40123] = i[78];
  assign o[40124] = i[78];
  assign o[40125] = i[78];
  assign o[40126] = i[78];
  assign o[40127] = i[78];
  assign o[40128] = i[78];
  assign o[40129] = i[78];
  assign o[40130] = i[78];
  assign o[40131] = i[78];
  assign o[40132] = i[78];
  assign o[40133] = i[78];
  assign o[40134] = i[78];
  assign o[40135] = i[78];
  assign o[40136] = i[78];
  assign o[40137] = i[78];
  assign o[40138] = i[78];
  assign o[40139] = i[78];
  assign o[40140] = i[78];
  assign o[40141] = i[78];
  assign o[40142] = i[78];
  assign o[40143] = i[78];
  assign o[40144] = i[78];
  assign o[40145] = i[78];
  assign o[40146] = i[78];
  assign o[40147] = i[78];
  assign o[40148] = i[78];
  assign o[40149] = i[78];
  assign o[40150] = i[78];
  assign o[40151] = i[78];
  assign o[40152] = i[78];
  assign o[40153] = i[78];
  assign o[40154] = i[78];
  assign o[40155] = i[78];
  assign o[40156] = i[78];
  assign o[40157] = i[78];
  assign o[40158] = i[78];
  assign o[40159] = i[78];
  assign o[40160] = i[78];
  assign o[40161] = i[78];
  assign o[40162] = i[78];
  assign o[40163] = i[78];
  assign o[40164] = i[78];
  assign o[40165] = i[78];
  assign o[40166] = i[78];
  assign o[40167] = i[78];
  assign o[40168] = i[78];
  assign o[40169] = i[78];
  assign o[40170] = i[78];
  assign o[40171] = i[78];
  assign o[40172] = i[78];
  assign o[40173] = i[78];
  assign o[40174] = i[78];
  assign o[40175] = i[78];
  assign o[40176] = i[78];
  assign o[40177] = i[78];
  assign o[40178] = i[78];
  assign o[40179] = i[78];
  assign o[40180] = i[78];
  assign o[40181] = i[78];
  assign o[40182] = i[78];
  assign o[40183] = i[78];
  assign o[40184] = i[78];
  assign o[40185] = i[78];
  assign o[40186] = i[78];
  assign o[40187] = i[78];
  assign o[40188] = i[78];
  assign o[40189] = i[78];
  assign o[40190] = i[78];
  assign o[40191] = i[78];
  assign o[40192] = i[78];
  assign o[40193] = i[78];
  assign o[40194] = i[78];
  assign o[40195] = i[78];
  assign o[40196] = i[78];
  assign o[40197] = i[78];
  assign o[40198] = i[78];
  assign o[40199] = i[78];
  assign o[40200] = i[78];
  assign o[40201] = i[78];
  assign o[40202] = i[78];
  assign o[40203] = i[78];
  assign o[40204] = i[78];
  assign o[40205] = i[78];
  assign o[40206] = i[78];
  assign o[40207] = i[78];
  assign o[40208] = i[78];
  assign o[40209] = i[78];
  assign o[40210] = i[78];
  assign o[40211] = i[78];
  assign o[40212] = i[78];
  assign o[40213] = i[78];
  assign o[40214] = i[78];
  assign o[40215] = i[78];
  assign o[40216] = i[78];
  assign o[40217] = i[78];
  assign o[40218] = i[78];
  assign o[40219] = i[78];
  assign o[40220] = i[78];
  assign o[40221] = i[78];
  assign o[40222] = i[78];
  assign o[40223] = i[78];
  assign o[40224] = i[78];
  assign o[40225] = i[78];
  assign o[40226] = i[78];
  assign o[40227] = i[78];
  assign o[40228] = i[78];
  assign o[40229] = i[78];
  assign o[40230] = i[78];
  assign o[40231] = i[78];
  assign o[40232] = i[78];
  assign o[40233] = i[78];
  assign o[40234] = i[78];
  assign o[40235] = i[78];
  assign o[40236] = i[78];
  assign o[40237] = i[78];
  assign o[40238] = i[78];
  assign o[40239] = i[78];
  assign o[40240] = i[78];
  assign o[40241] = i[78];
  assign o[40242] = i[78];
  assign o[40243] = i[78];
  assign o[40244] = i[78];
  assign o[40245] = i[78];
  assign o[40246] = i[78];
  assign o[40247] = i[78];
  assign o[40248] = i[78];
  assign o[40249] = i[78];
  assign o[40250] = i[78];
  assign o[40251] = i[78];
  assign o[40252] = i[78];
  assign o[40253] = i[78];
  assign o[40254] = i[78];
  assign o[40255] = i[78];
  assign o[40256] = i[78];
  assign o[40257] = i[78];
  assign o[40258] = i[78];
  assign o[40259] = i[78];
  assign o[40260] = i[78];
  assign o[40261] = i[78];
  assign o[40262] = i[78];
  assign o[40263] = i[78];
  assign o[40264] = i[78];
  assign o[40265] = i[78];
  assign o[40266] = i[78];
  assign o[40267] = i[78];
  assign o[40268] = i[78];
  assign o[40269] = i[78];
  assign o[40270] = i[78];
  assign o[40271] = i[78];
  assign o[40272] = i[78];
  assign o[40273] = i[78];
  assign o[40274] = i[78];
  assign o[40275] = i[78];
  assign o[40276] = i[78];
  assign o[40277] = i[78];
  assign o[40278] = i[78];
  assign o[40279] = i[78];
  assign o[40280] = i[78];
  assign o[40281] = i[78];
  assign o[40282] = i[78];
  assign o[40283] = i[78];
  assign o[40284] = i[78];
  assign o[40285] = i[78];
  assign o[40286] = i[78];
  assign o[40287] = i[78];
  assign o[40288] = i[78];
  assign o[40289] = i[78];
  assign o[40290] = i[78];
  assign o[40291] = i[78];
  assign o[40292] = i[78];
  assign o[40293] = i[78];
  assign o[40294] = i[78];
  assign o[40295] = i[78];
  assign o[40296] = i[78];
  assign o[40297] = i[78];
  assign o[40298] = i[78];
  assign o[40299] = i[78];
  assign o[40300] = i[78];
  assign o[40301] = i[78];
  assign o[40302] = i[78];
  assign o[40303] = i[78];
  assign o[40304] = i[78];
  assign o[40305] = i[78];
  assign o[40306] = i[78];
  assign o[40307] = i[78];
  assign o[40308] = i[78];
  assign o[40309] = i[78];
  assign o[40310] = i[78];
  assign o[40311] = i[78];
  assign o[40312] = i[78];
  assign o[40313] = i[78];
  assign o[40314] = i[78];
  assign o[40315] = i[78];
  assign o[40316] = i[78];
  assign o[40317] = i[78];
  assign o[40318] = i[78];
  assign o[40319] = i[78];
  assign o[40320] = i[78];
  assign o[40321] = i[78];
  assign o[40322] = i[78];
  assign o[40323] = i[78];
  assign o[40324] = i[78];
  assign o[40325] = i[78];
  assign o[40326] = i[78];
  assign o[40327] = i[78];
  assign o[40328] = i[78];
  assign o[40329] = i[78];
  assign o[40330] = i[78];
  assign o[40331] = i[78];
  assign o[40332] = i[78];
  assign o[40333] = i[78];
  assign o[40334] = i[78];
  assign o[40335] = i[78];
  assign o[40336] = i[78];
  assign o[40337] = i[78];
  assign o[40338] = i[78];
  assign o[40339] = i[78];
  assign o[40340] = i[78];
  assign o[40341] = i[78];
  assign o[40342] = i[78];
  assign o[40343] = i[78];
  assign o[40344] = i[78];
  assign o[40345] = i[78];
  assign o[40346] = i[78];
  assign o[40347] = i[78];
  assign o[40348] = i[78];
  assign o[40349] = i[78];
  assign o[40350] = i[78];
  assign o[40351] = i[78];
  assign o[40352] = i[78];
  assign o[40353] = i[78];
  assign o[40354] = i[78];
  assign o[40355] = i[78];
  assign o[40356] = i[78];
  assign o[40357] = i[78];
  assign o[40358] = i[78];
  assign o[40359] = i[78];
  assign o[40360] = i[78];
  assign o[40361] = i[78];
  assign o[40362] = i[78];
  assign o[40363] = i[78];
  assign o[40364] = i[78];
  assign o[40365] = i[78];
  assign o[40366] = i[78];
  assign o[40367] = i[78];
  assign o[40368] = i[78];
  assign o[40369] = i[78];
  assign o[40370] = i[78];
  assign o[40371] = i[78];
  assign o[40372] = i[78];
  assign o[40373] = i[78];
  assign o[40374] = i[78];
  assign o[40375] = i[78];
  assign o[40376] = i[78];
  assign o[40377] = i[78];
  assign o[40378] = i[78];
  assign o[40379] = i[78];
  assign o[40380] = i[78];
  assign o[40381] = i[78];
  assign o[40382] = i[78];
  assign o[40383] = i[78];
  assign o[40384] = i[78];
  assign o[40385] = i[78];
  assign o[40386] = i[78];
  assign o[40387] = i[78];
  assign o[40388] = i[78];
  assign o[40389] = i[78];
  assign o[40390] = i[78];
  assign o[40391] = i[78];
  assign o[40392] = i[78];
  assign o[40393] = i[78];
  assign o[40394] = i[78];
  assign o[40395] = i[78];
  assign o[40396] = i[78];
  assign o[40397] = i[78];
  assign o[40398] = i[78];
  assign o[40399] = i[78];
  assign o[40400] = i[78];
  assign o[40401] = i[78];
  assign o[40402] = i[78];
  assign o[40403] = i[78];
  assign o[40404] = i[78];
  assign o[40405] = i[78];
  assign o[40406] = i[78];
  assign o[40407] = i[78];
  assign o[40408] = i[78];
  assign o[40409] = i[78];
  assign o[40410] = i[78];
  assign o[40411] = i[78];
  assign o[40412] = i[78];
  assign o[40413] = i[78];
  assign o[40414] = i[78];
  assign o[40415] = i[78];
  assign o[40416] = i[78];
  assign o[40417] = i[78];
  assign o[40418] = i[78];
  assign o[40419] = i[78];
  assign o[40420] = i[78];
  assign o[40421] = i[78];
  assign o[40422] = i[78];
  assign o[40423] = i[78];
  assign o[40424] = i[78];
  assign o[40425] = i[78];
  assign o[40426] = i[78];
  assign o[40427] = i[78];
  assign o[40428] = i[78];
  assign o[40429] = i[78];
  assign o[40430] = i[78];
  assign o[40431] = i[78];
  assign o[40432] = i[78];
  assign o[40433] = i[78];
  assign o[40434] = i[78];
  assign o[40435] = i[78];
  assign o[40436] = i[78];
  assign o[40437] = i[78];
  assign o[40438] = i[78];
  assign o[40439] = i[78];
  assign o[40440] = i[78];
  assign o[40441] = i[78];
  assign o[40442] = i[78];
  assign o[40443] = i[78];
  assign o[40444] = i[78];
  assign o[40445] = i[78];
  assign o[40446] = i[78];
  assign o[40447] = i[78];
  assign o[39424] = i[77];
  assign o[39425] = i[77];
  assign o[39426] = i[77];
  assign o[39427] = i[77];
  assign o[39428] = i[77];
  assign o[39429] = i[77];
  assign o[39430] = i[77];
  assign o[39431] = i[77];
  assign o[39432] = i[77];
  assign o[39433] = i[77];
  assign o[39434] = i[77];
  assign o[39435] = i[77];
  assign o[39436] = i[77];
  assign o[39437] = i[77];
  assign o[39438] = i[77];
  assign o[39439] = i[77];
  assign o[39440] = i[77];
  assign o[39441] = i[77];
  assign o[39442] = i[77];
  assign o[39443] = i[77];
  assign o[39444] = i[77];
  assign o[39445] = i[77];
  assign o[39446] = i[77];
  assign o[39447] = i[77];
  assign o[39448] = i[77];
  assign o[39449] = i[77];
  assign o[39450] = i[77];
  assign o[39451] = i[77];
  assign o[39452] = i[77];
  assign o[39453] = i[77];
  assign o[39454] = i[77];
  assign o[39455] = i[77];
  assign o[39456] = i[77];
  assign o[39457] = i[77];
  assign o[39458] = i[77];
  assign o[39459] = i[77];
  assign o[39460] = i[77];
  assign o[39461] = i[77];
  assign o[39462] = i[77];
  assign o[39463] = i[77];
  assign o[39464] = i[77];
  assign o[39465] = i[77];
  assign o[39466] = i[77];
  assign o[39467] = i[77];
  assign o[39468] = i[77];
  assign o[39469] = i[77];
  assign o[39470] = i[77];
  assign o[39471] = i[77];
  assign o[39472] = i[77];
  assign o[39473] = i[77];
  assign o[39474] = i[77];
  assign o[39475] = i[77];
  assign o[39476] = i[77];
  assign o[39477] = i[77];
  assign o[39478] = i[77];
  assign o[39479] = i[77];
  assign o[39480] = i[77];
  assign o[39481] = i[77];
  assign o[39482] = i[77];
  assign o[39483] = i[77];
  assign o[39484] = i[77];
  assign o[39485] = i[77];
  assign o[39486] = i[77];
  assign o[39487] = i[77];
  assign o[39488] = i[77];
  assign o[39489] = i[77];
  assign o[39490] = i[77];
  assign o[39491] = i[77];
  assign o[39492] = i[77];
  assign o[39493] = i[77];
  assign o[39494] = i[77];
  assign o[39495] = i[77];
  assign o[39496] = i[77];
  assign o[39497] = i[77];
  assign o[39498] = i[77];
  assign o[39499] = i[77];
  assign o[39500] = i[77];
  assign o[39501] = i[77];
  assign o[39502] = i[77];
  assign o[39503] = i[77];
  assign o[39504] = i[77];
  assign o[39505] = i[77];
  assign o[39506] = i[77];
  assign o[39507] = i[77];
  assign o[39508] = i[77];
  assign o[39509] = i[77];
  assign o[39510] = i[77];
  assign o[39511] = i[77];
  assign o[39512] = i[77];
  assign o[39513] = i[77];
  assign o[39514] = i[77];
  assign o[39515] = i[77];
  assign o[39516] = i[77];
  assign o[39517] = i[77];
  assign o[39518] = i[77];
  assign o[39519] = i[77];
  assign o[39520] = i[77];
  assign o[39521] = i[77];
  assign o[39522] = i[77];
  assign o[39523] = i[77];
  assign o[39524] = i[77];
  assign o[39525] = i[77];
  assign o[39526] = i[77];
  assign o[39527] = i[77];
  assign o[39528] = i[77];
  assign o[39529] = i[77];
  assign o[39530] = i[77];
  assign o[39531] = i[77];
  assign o[39532] = i[77];
  assign o[39533] = i[77];
  assign o[39534] = i[77];
  assign o[39535] = i[77];
  assign o[39536] = i[77];
  assign o[39537] = i[77];
  assign o[39538] = i[77];
  assign o[39539] = i[77];
  assign o[39540] = i[77];
  assign o[39541] = i[77];
  assign o[39542] = i[77];
  assign o[39543] = i[77];
  assign o[39544] = i[77];
  assign o[39545] = i[77];
  assign o[39546] = i[77];
  assign o[39547] = i[77];
  assign o[39548] = i[77];
  assign o[39549] = i[77];
  assign o[39550] = i[77];
  assign o[39551] = i[77];
  assign o[39552] = i[77];
  assign o[39553] = i[77];
  assign o[39554] = i[77];
  assign o[39555] = i[77];
  assign o[39556] = i[77];
  assign o[39557] = i[77];
  assign o[39558] = i[77];
  assign o[39559] = i[77];
  assign o[39560] = i[77];
  assign o[39561] = i[77];
  assign o[39562] = i[77];
  assign o[39563] = i[77];
  assign o[39564] = i[77];
  assign o[39565] = i[77];
  assign o[39566] = i[77];
  assign o[39567] = i[77];
  assign o[39568] = i[77];
  assign o[39569] = i[77];
  assign o[39570] = i[77];
  assign o[39571] = i[77];
  assign o[39572] = i[77];
  assign o[39573] = i[77];
  assign o[39574] = i[77];
  assign o[39575] = i[77];
  assign o[39576] = i[77];
  assign o[39577] = i[77];
  assign o[39578] = i[77];
  assign o[39579] = i[77];
  assign o[39580] = i[77];
  assign o[39581] = i[77];
  assign o[39582] = i[77];
  assign o[39583] = i[77];
  assign o[39584] = i[77];
  assign o[39585] = i[77];
  assign o[39586] = i[77];
  assign o[39587] = i[77];
  assign o[39588] = i[77];
  assign o[39589] = i[77];
  assign o[39590] = i[77];
  assign o[39591] = i[77];
  assign o[39592] = i[77];
  assign o[39593] = i[77];
  assign o[39594] = i[77];
  assign o[39595] = i[77];
  assign o[39596] = i[77];
  assign o[39597] = i[77];
  assign o[39598] = i[77];
  assign o[39599] = i[77];
  assign o[39600] = i[77];
  assign o[39601] = i[77];
  assign o[39602] = i[77];
  assign o[39603] = i[77];
  assign o[39604] = i[77];
  assign o[39605] = i[77];
  assign o[39606] = i[77];
  assign o[39607] = i[77];
  assign o[39608] = i[77];
  assign o[39609] = i[77];
  assign o[39610] = i[77];
  assign o[39611] = i[77];
  assign o[39612] = i[77];
  assign o[39613] = i[77];
  assign o[39614] = i[77];
  assign o[39615] = i[77];
  assign o[39616] = i[77];
  assign o[39617] = i[77];
  assign o[39618] = i[77];
  assign o[39619] = i[77];
  assign o[39620] = i[77];
  assign o[39621] = i[77];
  assign o[39622] = i[77];
  assign o[39623] = i[77];
  assign o[39624] = i[77];
  assign o[39625] = i[77];
  assign o[39626] = i[77];
  assign o[39627] = i[77];
  assign o[39628] = i[77];
  assign o[39629] = i[77];
  assign o[39630] = i[77];
  assign o[39631] = i[77];
  assign o[39632] = i[77];
  assign o[39633] = i[77];
  assign o[39634] = i[77];
  assign o[39635] = i[77];
  assign o[39636] = i[77];
  assign o[39637] = i[77];
  assign o[39638] = i[77];
  assign o[39639] = i[77];
  assign o[39640] = i[77];
  assign o[39641] = i[77];
  assign o[39642] = i[77];
  assign o[39643] = i[77];
  assign o[39644] = i[77];
  assign o[39645] = i[77];
  assign o[39646] = i[77];
  assign o[39647] = i[77];
  assign o[39648] = i[77];
  assign o[39649] = i[77];
  assign o[39650] = i[77];
  assign o[39651] = i[77];
  assign o[39652] = i[77];
  assign o[39653] = i[77];
  assign o[39654] = i[77];
  assign o[39655] = i[77];
  assign o[39656] = i[77];
  assign o[39657] = i[77];
  assign o[39658] = i[77];
  assign o[39659] = i[77];
  assign o[39660] = i[77];
  assign o[39661] = i[77];
  assign o[39662] = i[77];
  assign o[39663] = i[77];
  assign o[39664] = i[77];
  assign o[39665] = i[77];
  assign o[39666] = i[77];
  assign o[39667] = i[77];
  assign o[39668] = i[77];
  assign o[39669] = i[77];
  assign o[39670] = i[77];
  assign o[39671] = i[77];
  assign o[39672] = i[77];
  assign o[39673] = i[77];
  assign o[39674] = i[77];
  assign o[39675] = i[77];
  assign o[39676] = i[77];
  assign o[39677] = i[77];
  assign o[39678] = i[77];
  assign o[39679] = i[77];
  assign o[39680] = i[77];
  assign o[39681] = i[77];
  assign o[39682] = i[77];
  assign o[39683] = i[77];
  assign o[39684] = i[77];
  assign o[39685] = i[77];
  assign o[39686] = i[77];
  assign o[39687] = i[77];
  assign o[39688] = i[77];
  assign o[39689] = i[77];
  assign o[39690] = i[77];
  assign o[39691] = i[77];
  assign o[39692] = i[77];
  assign o[39693] = i[77];
  assign o[39694] = i[77];
  assign o[39695] = i[77];
  assign o[39696] = i[77];
  assign o[39697] = i[77];
  assign o[39698] = i[77];
  assign o[39699] = i[77];
  assign o[39700] = i[77];
  assign o[39701] = i[77];
  assign o[39702] = i[77];
  assign o[39703] = i[77];
  assign o[39704] = i[77];
  assign o[39705] = i[77];
  assign o[39706] = i[77];
  assign o[39707] = i[77];
  assign o[39708] = i[77];
  assign o[39709] = i[77];
  assign o[39710] = i[77];
  assign o[39711] = i[77];
  assign o[39712] = i[77];
  assign o[39713] = i[77];
  assign o[39714] = i[77];
  assign o[39715] = i[77];
  assign o[39716] = i[77];
  assign o[39717] = i[77];
  assign o[39718] = i[77];
  assign o[39719] = i[77];
  assign o[39720] = i[77];
  assign o[39721] = i[77];
  assign o[39722] = i[77];
  assign o[39723] = i[77];
  assign o[39724] = i[77];
  assign o[39725] = i[77];
  assign o[39726] = i[77];
  assign o[39727] = i[77];
  assign o[39728] = i[77];
  assign o[39729] = i[77];
  assign o[39730] = i[77];
  assign o[39731] = i[77];
  assign o[39732] = i[77];
  assign o[39733] = i[77];
  assign o[39734] = i[77];
  assign o[39735] = i[77];
  assign o[39736] = i[77];
  assign o[39737] = i[77];
  assign o[39738] = i[77];
  assign o[39739] = i[77];
  assign o[39740] = i[77];
  assign o[39741] = i[77];
  assign o[39742] = i[77];
  assign o[39743] = i[77];
  assign o[39744] = i[77];
  assign o[39745] = i[77];
  assign o[39746] = i[77];
  assign o[39747] = i[77];
  assign o[39748] = i[77];
  assign o[39749] = i[77];
  assign o[39750] = i[77];
  assign o[39751] = i[77];
  assign o[39752] = i[77];
  assign o[39753] = i[77];
  assign o[39754] = i[77];
  assign o[39755] = i[77];
  assign o[39756] = i[77];
  assign o[39757] = i[77];
  assign o[39758] = i[77];
  assign o[39759] = i[77];
  assign o[39760] = i[77];
  assign o[39761] = i[77];
  assign o[39762] = i[77];
  assign o[39763] = i[77];
  assign o[39764] = i[77];
  assign o[39765] = i[77];
  assign o[39766] = i[77];
  assign o[39767] = i[77];
  assign o[39768] = i[77];
  assign o[39769] = i[77];
  assign o[39770] = i[77];
  assign o[39771] = i[77];
  assign o[39772] = i[77];
  assign o[39773] = i[77];
  assign o[39774] = i[77];
  assign o[39775] = i[77];
  assign o[39776] = i[77];
  assign o[39777] = i[77];
  assign o[39778] = i[77];
  assign o[39779] = i[77];
  assign o[39780] = i[77];
  assign o[39781] = i[77];
  assign o[39782] = i[77];
  assign o[39783] = i[77];
  assign o[39784] = i[77];
  assign o[39785] = i[77];
  assign o[39786] = i[77];
  assign o[39787] = i[77];
  assign o[39788] = i[77];
  assign o[39789] = i[77];
  assign o[39790] = i[77];
  assign o[39791] = i[77];
  assign o[39792] = i[77];
  assign o[39793] = i[77];
  assign o[39794] = i[77];
  assign o[39795] = i[77];
  assign o[39796] = i[77];
  assign o[39797] = i[77];
  assign o[39798] = i[77];
  assign o[39799] = i[77];
  assign o[39800] = i[77];
  assign o[39801] = i[77];
  assign o[39802] = i[77];
  assign o[39803] = i[77];
  assign o[39804] = i[77];
  assign o[39805] = i[77];
  assign o[39806] = i[77];
  assign o[39807] = i[77];
  assign o[39808] = i[77];
  assign o[39809] = i[77];
  assign o[39810] = i[77];
  assign o[39811] = i[77];
  assign o[39812] = i[77];
  assign o[39813] = i[77];
  assign o[39814] = i[77];
  assign o[39815] = i[77];
  assign o[39816] = i[77];
  assign o[39817] = i[77];
  assign o[39818] = i[77];
  assign o[39819] = i[77];
  assign o[39820] = i[77];
  assign o[39821] = i[77];
  assign o[39822] = i[77];
  assign o[39823] = i[77];
  assign o[39824] = i[77];
  assign o[39825] = i[77];
  assign o[39826] = i[77];
  assign o[39827] = i[77];
  assign o[39828] = i[77];
  assign o[39829] = i[77];
  assign o[39830] = i[77];
  assign o[39831] = i[77];
  assign o[39832] = i[77];
  assign o[39833] = i[77];
  assign o[39834] = i[77];
  assign o[39835] = i[77];
  assign o[39836] = i[77];
  assign o[39837] = i[77];
  assign o[39838] = i[77];
  assign o[39839] = i[77];
  assign o[39840] = i[77];
  assign o[39841] = i[77];
  assign o[39842] = i[77];
  assign o[39843] = i[77];
  assign o[39844] = i[77];
  assign o[39845] = i[77];
  assign o[39846] = i[77];
  assign o[39847] = i[77];
  assign o[39848] = i[77];
  assign o[39849] = i[77];
  assign o[39850] = i[77];
  assign o[39851] = i[77];
  assign o[39852] = i[77];
  assign o[39853] = i[77];
  assign o[39854] = i[77];
  assign o[39855] = i[77];
  assign o[39856] = i[77];
  assign o[39857] = i[77];
  assign o[39858] = i[77];
  assign o[39859] = i[77];
  assign o[39860] = i[77];
  assign o[39861] = i[77];
  assign o[39862] = i[77];
  assign o[39863] = i[77];
  assign o[39864] = i[77];
  assign o[39865] = i[77];
  assign o[39866] = i[77];
  assign o[39867] = i[77];
  assign o[39868] = i[77];
  assign o[39869] = i[77];
  assign o[39870] = i[77];
  assign o[39871] = i[77];
  assign o[39872] = i[77];
  assign o[39873] = i[77];
  assign o[39874] = i[77];
  assign o[39875] = i[77];
  assign o[39876] = i[77];
  assign o[39877] = i[77];
  assign o[39878] = i[77];
  assign o[39879] = i[77];
  assign o[39880] = i[77];
  assign o[39881] = i[77];
  assign o[39882] = i[77];
  assign o[39883] = i[77];
  assign o[39884] = i[77];
  assign o[39885] = i[77];
  assign o[39886] = i[77];
  assign o[39887] = i[77];
  assign o[39888] = i[77];
  assign o[39889] = i[77];
  assign o[39890] = i[77];
  assign o[39891] = i[77];
  assign o[39892] = i[77];
  assign o[39893] = i[77];
  assign o[39894] = i[77];
  assign o[39895] = i[77];
  assign o[39896] = i[77];
  assign o[39897] = i[77];
  assign o[39898] = i[77];
  assign o[39899] = i[77];
  assign o[39900] = i[77];
  assign o[39901] = i[77];
  assign o[39902] = i[77];
  assign o[39903] = i[77];
  assign o[39904] = i[77];
  assign o[39905] = i[77];
  assign o[39906] = i[77];
  assign o[39907] = i[77];
  assign o[39908] = i[77];
  assign o[39909] = i[77];
  assign o[39910] = i[77];
  assign o[39911] = i[77];
  assign o[39912] = i[77];
  assign o[39913] = i[77];
  assign o[39914] = i[77];
  assign o[39915] = i[77];
  assign o[39916] = i[77];
  assign o[39917] = i[77];
  assign o[39918] = i[77];
  assign o[39919] = i[77];
  assign o[39920] = i[77];
  assign o[39921] = i[77];
  assign o[39922] = i[77];
  assign o[39923] = i[77];
  assign o[39924] = i[77];
  assign o[39925] = i[77];
  assign o[39926] = i[77];
  assign o[39927] = i[77];
  assign o[39928] = i[77];
  assign o[39929] = i[77];
  assign o[39930] = i[77];
  assign o[39931] = i[77];
  assign o[39932] = i[77];
  assign o[39933] = i[77];
  assign o[39934] = i[77];
  assign o[39935] = i[77];
  assign o[38912] = i[76];
  assign o[38913] = i[76];
  assign o[38914] = i[76];
  assign o[38915] = i[76];
  assign o[38916] = i[76];
  assign o[38917] = i[76];
  assign o[38918] = i[76];
  assign o[38919] = i[76];
  assign o[38920] = i[76];
  assign o[38921] = i[76];
  assign o[38922] = i[76];
  assign o[38923] = i[76];
  assign o[38924] = i[76];
  assign o[38925] = i[76];
  assign o[38926] = i[76];
  assign o[38927] = i[76];
  assign o[38928] = i[76];
  assign o[38929] = i[76];
  assign o[38930] = i[76];
  assign o[38931] = i[76];
  assign o[38932] = i[76];
  assign o[38933] = i[76];
  assign o[38934] = i[76];
  assign o[38935] = i[76];
  assign o[38936] = i[76];
  assign o[38937] = i[76];
  assign o[38938] = i[76];
  assign o[38939] = i[76];
  assign o[38940] = i[76];
  assign o[38941] = i[76];
  assign o[38942] = i[76];
  assign o[38943] = i[76];
  assign o[38944] = i[76];
  assign o[38945] = i[76];
  assign o[38946] = i[76];
  assign o[38947] = i[76];
  assign o[38948] = i[76];
  assign o[38949] = i[76];
  assign o[38950] = i[76];
  assign o[38951] = i[76];
  assign o[38952] = i[76];
  assign o[38953] = i[76];
  assign o[38954] = i[76];
  assign o[38955] = i[76];
  assign o[38956] = i[76];
  assign o[38957] = i[76];
  assign o[38958] = i[76];
  assign o[38959] = i[76];
  assign o[38960] = i[76];
  assign o[38961] = i[76];
  assign o[38962] = i[76];
  assign o[38963] = i[76];
  assign o[38964] = i[76];
  assign o[38965] = i[76];
  assign o[38966] = i[76];
  assign o[38967] = i[76];
  assign o[38968] = i[76];
  assign o[38969] = i[76];
  assign o[38970] = i[76];
  assign o[38971] = i[76];
  assign o[38972] = i[76];
  assign o[38973] = i[76];
  assign o[38974] = i[76];
  assign o[38975] = i[76];
  assign o[38976] = i[76];
  assign o[38977] = i[76];
  assign o[38978] = i[76];
  assign o[38979] = i[76];
  assign o[38980] = i[76];
  assign o[38981] = i[76];
  assign o[38982] = i[76];
  assign o[38983] = i[76];
  assign o[38984] = i[76];
  assign o[38985] = i[76];
  assign o[38986] = i[76];
  assign o[38987] = i[76];
  assign o[38988] = i[76];
  assign o[38989] = i[76];
  assign o[38990] = i[76];
  assign o[38991] = i[76];
  assign o[38992] = i[76];
  assign o[38993] = i[76];
  assign o[38994] = i[76];
  assign o[38995] = i[76];
  assign o[38996] = i[76];
  assign o[38997] = i[76];
  assign o[38998] = i[76];
  assign o[38999] = i[76];
  assign o[39000] = i[76];
  assign o[39001] = i[76];
  assign o[39002] = i[76];
  assign o[39003] = i[76];
  assign o[39004] = i[76];
  assign o[39005] = i[76];
  assign o[39006] = i[76];
  assign o[39007] = i[76];
  assign o[39008] = i[76];
  assign o[39009] = i[76];
  assign o[39010] = i[76];
  assign o[39011] = i[76];
  assign o[39012] = i[76];
  assign o[39013] = i[76];
  assign o[39014] = i[76];
  assign o[39015] = i[76];
  assign o[39016] = i[76];
  assign o[39017] = i[76];
  assign o[39018] = i[76];
  assign o[39019] = i[76];
  assign o[39020] = i[76];
  assign o[39021] = i[76];
  assign o[39022] = i[76];
  assign o[39023] = i[76];
  assign o[39024] = i[76];
  assign o[39025] = i[76];
  assign o[39026] = i[76];
  assign o[39027] = i[76];
  assign o[39028] = i[76];
  assign o[39029] = i[76];
  assign o[39030] = i[76];
  assign o[39031] = i[76];
  assign o[39032] = i[76];
  assign o[39033] = i[76];
  assign o[39034] = i[76];
  assign o[39035] = i[76];
  assign o[39036] = i[76];
  assign o[39037] = i[76];
  assign o[39038] = i[76];
  assign o[39039] = i[76];
  assign o[39040] = i[76];
  assign o[39041] = i[76];
  assign o[39042] = i[76];
  assign o[39043] = i[76];
  assign o[39044] = i[76];
  assign o[39045] = i[76];
  assign o[39046] = i[76];
  assign o[39047] = i[76];
  assign o[39048] = i[76];
  assign o[39049] = i[76];
  assign o[39050] = i[76];
  assign o[39051] = i[76];
  assign o[39052] = i[76];
  assign o[39053] = i[76];
  assign o[39054] = i[76];
  assign o[39055] = i[76];
  assign o[39056] = i[76];
  assign o[39057] = i[76];
  assign o[39058] = i[76];
  assign o[39059] = i[76];
  assign o[39060] = i[76];
  assign o[39061] = i[76];
  assign o[39062] = i[76];
  assign o[39063] = i[76];
  assign o[39064] = i[76];
  assign o[39065] = i[76];
  assign o[39066] = i[76];
  assign o[39067] = i[76];
  assign o[39068] = i[76];
  assign o[39069] = i[76];
  assign o[39070] = i[76];
  assign o[39071] = i[76];
  assign o[39072] = i[76];
  assign o[39073] = i[76];
  assign o[39074] = i[76];
  assign o[39075] = i[76];
  assign o[39076] = i[76];
  assign o[39077] = i[76];
  assign o[39078] = i[76];
  assign o[39079] = i[76];
  assign o[39080] = i[76];
  assign o[39081] = i[76];
  assign o[39082] = i[76];
  assign o[39083] = i[76];
  assign o[39084] = i[76];
  assign o[39085] = i[76];
  assign o[39086] = i[76];
  assign o[39087] = i[76];
  assign o[39088] = i[76];
  assign o[39089] = i[76];
  assign o[39090] = i[76];
  assign o[39091] = i[76];
  assign o[39092] = i[76];
  assign o[39093] = i[76];
  assign o[39094] = i[76];
  assign o[39095] = i[76];
  assign o[39096] = i[76];
  assign o[39097] = i[76];
  assign o[39098] = i[76];
  assign o[39099] = i[76];
  assign o[39100] = i[76];
  assign o[39101] = i[76];
  assign o[39102] = i[76];
  assign o[39103] = i[76];
  assign o[39104] = i[76];
  assign o[39105] = i[76];
  assign o[39106] = i[76];
  assign o[39107] = i[76];
  assign o[39108] = i[76];
  assign o[39109] = i[76];
  assign o[39110] = i[76];
  assign o[39111] = i[76];
  assign o[39112] = i[76];
  assign o[39113] = i[76];
  assign o[39114] = i[76];
  assign o[39115] = i[76];
  assign o[39116] = i[76];
  assign o[39117] = i[76];
  assign o[39118] = i[76];
  assign o[39119] = i[76];
  assign o[39120] = i[76];
  assign o[39121] = i[76];
  assign o[39122] = i[76];
  assign o[39123] = i[76];
  assign o[39124] = i[76];
  assign o[39125] = i[76];
  assign o[39126] = i[76];
  assign o[39127] = i[76];
  assign o[39128] = i[76];
  assign o[39129] = i[76];
  assign o[39130] = i[76];
  assign o[39131] = i[76];
  assign o[39132] = i[76];
  assign o[39133] = i[76];
  assign o[39134] = i[76];
  assign o[39135] = i[76];
  assign o[39136] = i[76];
  assign o[39137] = i[76];
  assign o[39138] = i[76];
  assign o[39139] = i[76];
  assign o[39140] = i[76];
  assign o[39141] = i[76];
  assign o[39142] = i[76];
  assign o[39143] = i[76];
  assign o[39144] = i[76];
  assign o[39145] = i[76];
  assign o[39146] = i[76];
  assign o[39147] = i[76];
  assign o[39148] = i[76];
  assign o[39149] = i[76];
  assign o[39150] = i[76];
  assign o[39151] = i[76];
  assign o[39152] = i[76];
  assign o[39153] = i[76];
  assign o[39154] = i[76];
  assign o[39155] = i[76];
  assign o[39156] = i[76];
  assign o[39157] = i[76];
  assign o[39158] = i[76];
  assign o[39159] = i[76];
  assign o[39160] = i[76];
  assign o[39161] = i[76];
  assign o[39162] = i[76];
  assign o[39163] = i[76];
  assign o[39164] = i[76];
  assign o[39165] = i[76];
  assign o[39166] = i[76];
  assign o[39167] = i[76];
  assign o[39168] = i[76];
  assign o[39169] = i[76];
  assign o[39170] = i[76];
  assign o[39171] = i[76];
  assign o[39172] = i[76];
  assign o[39173] = i[76];
  assign o[39174] = i[76];
  assign o[39175] = i[76];
  assign o[39176] = i[76];
  assign o[39177] = i[76];
  assign o[39178] = i[76];
  assign o[39179] = i[76];
  assign o[39180] = i[76];
  assign o[39181] = i[76];
  assign o[39182] = i[76];
  assign o[39183] = i[76];
  assign o[39184] = i[76];
  assign o[39185] = i[76];
  assign o[39186] = i[76];
  assign o[39187] = i[76];
  assign o[39188] = i[76];
  assign o[39189] = i[76];
  assign o[39190] = i[76];
  assign o[39191] = i[76];
  assign o[39192] = i[76];
  assign o[39193] = i[76];
  assign o[39194] = i[76];
  assign o[39195] = i[76];
  assign o[39196] = i[76];
  assign o[39197] = i[76];
  assign o[39198] = i[76];
  assign o[39199] = i[76];
  assign o[39200] = i[76];
  assign o[39201] = i[76];
  assign o[39202] = i[76];
  assign o[39203] = i[76];
  assign o[39204] = i[76];
  assign o[39205] = i[76];
  assign o[39206] = i[76];
  assign o[39207] = i[76];
  assign o[39208] = i[76];
  assign o[39209] = i[76];
  assign o[39210] = i[76];
  assign o[39211] = i[76];
  assign o[39212] = i[76];
  assign o[39213] = i[76];
  assign o[39214] = i[76];
  assign o[39215] = i[76];
  assign o[39216] = i[76];
  assign o[39217] = i[76];
  assign o[39218] = i[76];
  assign o[39219] = i[76];
  assign o[39220] = i[76];
  assign o[39221] = i[76];
  assign o[39222] = i[76];
  assign o[39223] = i[76];
  assign o[39224] = i[76];
  assign o[39225] = i[76];
  assign o[39226] = i[76];
  assign o[39227] = i[76];
  assign o[39228] = i[76];
  assign o[39229] = i[76];
  assign o[39230] = i[76];
  assign o[39231] = i[76];
  assign o[39232] = i[76];
  assign o[39233] = i[76];
  assign o[39234] = i[76];
  assign o[39235] = i[76];
  assign o[39236] = i[76];
  assign o[39237] = i[76];
  assign o[39238] = i[76];
  assign o[39239] = i[76];
  assign o[39240] = i[76];
  assign o[39241] = i[76];
  assign o[39242] = i[76];
  assign o[39243] = i[76];
  assign o[39244] = i[76];
  assign o[39245] = i[76];
  assign o[39246] = i[76];
  assign o[39247] = i[76];
  assign o[39248] = i[76];
  assign o[39249] = i[76];
  assign o[39250] = i[76];
  assign o[39251] = i[76];
  assign o[39252] = i[76];
  assign o[39253] = i[76];
  assign o[39254] = i[76];
  assign o[39255] = i[76];
  assign o[39256] = i[76];
  assign o[39257] = i[76];
  assign o[39258] = i[76];
  assign o[39259] = i[76];
  assign o[39260] = i[76];
  assign o[39261] = i[76];
  assign o[39262] = i[76];
  assign o[39263] = i[76];
  assign o[39264] = i[76];
  assign o[39265] = i[76];
  assign o[39266] = i[76];
  assign o[39267] = i[76];
  assign o[39268] = i[76];
  assign o[39269] = i[76];
  assign o[39270] = i[76];
  assign o[39271] = i[76];
  assign o[39272] = i[76];
  assign o[39273] = i[76];
  assign o[39274] = i[76];
  assign o[39275] = i[76];
  assign o[39276] = i[76];
  assign o[39277] = i[76];
  assign o[39278] = i[76];
  assign o[39279] = i[76];
  assign o[39280] = i[76];
  assign o[39281] = i[76];
  assign o[39282] = i[76];
  assign o[39283] = i[76];
  assign o[39284] = i[76];
  assign o[39285] = i[76];
  assign o[39286] = i[76];
  assign o[39287] = i[76];
  assign o[39288] = i[76];
  assign o[39289] = i[76];
  assign o[39290] = i[76];
  assign o[39291] = i[76];
  assign o[39292] = i[76];
  assign o[39293] = i[76];
  assign o[39294] = i[76];
  assign o[39295] = i[76];
  assign o[39296] = i[76];
  assign o[39297] = i[76];
  assign o[39298] = i[76];
  assign o[39299] = i[76];
  assign o[39300] = i[76];
  assign o[39301] = i[76];
  assign o[39302] = i[76];
  assign o[39303] = i[76];
  assign o[39304] = i[76];
  assign o[39305] = i[76];
  assign o[39306] = i[76];
  assign o[39307] = i[76];
  assign o[39308] = i[76];
  assign o[39309] = i[76];
  assign o[39310] = i[76];
  assign o[39311] = i[76];
  assign o[39312] = i[76];
  assign o[39313] = i[76];
  assign o[39314] = i[76];
  assign o[39315] = i[76];
  assign o[39316] = i[76];
  assign o[39317] = i[76];
  assign o[39318] = i[76];
  assign o[39319] = i[76];
  assign o[39320] = i[76];
  assign o[39321] = i[76];
  assign o[39322] = i[76];
  assign o[39323] = i[76];
  assign o[39324] = i[76];
  assign o[39325] = i[76];
  assign o[39326] = i[76];
  assign o[39327] = i[76];
  assign o[39328] = i[76];
  assign o[39329] = i[76];
  assign o[39330] = i[76];
  assign o[39331] = i[76];
  assign o[39332] = i[76];
  assign o[39333] = i[76];
  assign o[39334] = i[76];
  assign o[39335] = i[76];
  assign o[39336] = i[76];
  assign o[39337] = i[76];
  assign o[39338] = i[76];
  assign o[39339] = i[76];
  assign o[39340] = i[76];
  assign o[39341] = i[76];
  assign o[39342] = i[76];
  assign o[39343] = i[76];
  assign o[39344] = i[76];
  assign o[39345] = i[76];
  assign o[39346] = i[76];
  assign o[39347] = i[76];
  assign o[39348] = i[76];
  assign o[39349] = i[76];
  assign o[39350] = i[76];
  assign o[39351] = i[76];
  assign o[39352] = i[76];
  assign o[39353] = i[76];
  assign o[39354] = i[76];
  assign o[39355] = i[76];
  assign o[39356] = i[76];
  assign o[39357] = i[76];
  assign o[39358] = i[76];
  assign o[39359] = i[76];
  assign o[39360] = i[76];
  assign o[39361] = i[76];
  assign o[39362] = i[76];
  assign o[39363] = i[76];
  assign o[39364] = i[76];
  assign o[39365] = i[76];
  assign o[39366] = i[76];
  assign o[39367] = i[76];
  assign o[39368] = i[76];
  assign o[39369] = i[76];
  assign o[39370] = i[76];
  assign o[39371] = i[76];
  assign o[39372] = i[76];
  assign o[39373] = i[76];
  assign o[39374] = i[76];
  assign o[39375] = i[76];
  assign o[39376] = i[76];
  assign o[39377] = i[76];
  assign o[39378] = i[76];
  assign o[39379] = i[76];
  assign o[39380] = i[76];
  assign o[39381] = i[76];
  assign o[39382] = i[76];
  assign o[39383] = i[76];
  assign o[39384] = i[76];
  assign o[39385] = i[76];
  assign o[39386] = i[76];
  assign o[39387] = i[76];
  assign o[39388] = i[76];
  assign o[39389] = i[76];
  assign o[39390] = i[76];
  assign o[39391] = i[76];
  assign o[39392] = i[76];
  assign o[39393] = i[76];
  assign o[39394] = i[76];
  assign o[39395] = i[76];
  assign o[39396] = i[76];
  assign o[39397] = i[76];
  assign o[39398] = i[76];
  assign o[39399] = i[76];
  assign o[39400] = i[76];
  assign o[39401] = i[76];
  assign o[39402] = i[76];
  assign o[39403] = i[76];
  assign o[39404] = i[76];
  assign o[39405] = i[76];
  assign o[39406] = i[76];
  assign o[39407] = i[76];
  assign o[39408] = i[76];
  assign o[39409] = i[76];
  assign o[39410] = i[76];
  assign o[39411] = i[76];
  assign o[39412] = i[76];
  assign o[39413] = i[76];
  assign o[39414] = i[76];
  assign o[39415] = i[76];
  assign o[39416] = i[76];
  assign o[39417] = i[76];
  assign o[39418] = i[76];
  assign o[39419] = i[76];
  assign o[39420] = i[76];
  assign o[39421] = i[76];
  assign o[39422] = i[76];
  assign o[39423] = i[76];
  assign o[38400] = i[75];
  assign o[38401] = i[75];
  assign o[38402] = i[75];
  assign o[38403] = i[75];
  assign o[38404] = i[75];
  assign o[38405] = i[75];
  assign o[38406] = i[75];
  assign o[38407] = i[75];
  assign o[38408] = i[75];
  assign o[38409] = i[75];
  assign o[38410] = i[75];
  assign o[38411] = i[75];
  assign o[38412] = i[75];
  assign o[38413] = i[75];
  assign o[38414] = i[75];
  assign o[38415] = i[75];
  assign o[38416] = i[75];
  assign o[38417] = i[75];
  assign o[38418] = i[75];
  assign o[38419] = i[75];
  assign o[38420] = i[75];
  assign o[38421] = i[75];
  assign o[38422] = i[75];
  assign o[38423] = i[75];
  assign o[38424] = i[75];
  assign o[38425] = i[75];
  assign o[38426] = i[75];
  assign o[38427] = i[75];
  assign o[38428] = i[75];
  assign o[38429] = i[75];
  assign o[38430] = i[75];
  assign o[38431] = i[75];
  assign o[38432] = i[75];
  assign o[38433] = i[75];
  assign o[38434] = i[75];
  assign o[38435] = i[75];
  assign o[38436] = i[75];
  assign o[38437] = i[75];
  assign o[38438] = i[75];
  assign o[38439] = i[75];
  assign o[38440] = i[75];
  assign o[38441] = i[75];
  assign o[38442] = i[75];
  assign o[38443] = i[75];
  assign o[38444] = i[75];
  assign o[38445] = i[75];
  assign o[38446] = i[75];
  assign o[38447] = i[75];
  assign o[38448] = i[75];
  assign o[38449] = i[75];
  assign o[38450] = i[75];
  assign o[38451] = i[75];
  assign o[38452] = i[75];
  assign o[38453] = i[75];
  assign o[38454] = i[75];
  assign o[38455] = i[75];
  assign o[38456] = i[75];
  assign o[38457] = i[75];
  assign o[38458] = i[75];
  assign o[38459] = i[75];
  assign o[38460] = i[75];
  assign o[38461] = i[75];
  assign o[38462] = i[75];
  assign o[38463] = i[75];
  assign o[38464] = i[75];
  assign o[38465] = i[75];
  assign o[38466] = i[75];
  assign o[38467] = i[75];
  assign o[38468] = i[75];
  assign o[38469] = i[75];
  assign o[38470] = i[75];
  assign o[38471] = i[75];
  assign o[38472] = i[75];
  assign o[38473] = i[75];
  assign o[38474] = i[75];
  assign o[38475] = i[75];
  assign o[38476] = i[75];
  assign o[38477] = i[75];
  assign o[38478] = i[75];
  assign o[38479] = i[75];
  assign o[38480] = i[75];
  assign o[38481] = i[75];
  assign o[38482] = i[75];
  assign o[38483] = i[75];
  assign o[38484] = i[75];
  assign o[38485] = i[75];
  assign o[38486] = i[75];
  assign o[38487] = i[75];
  assign o[38488] = i[75];
  assign o[38489] = i[75];
  assign o[38490] = i[75];
  assign o[38491] = i[75];
  assign o[38492] = i[75];
  assign o[38493] = i[75];
  assign o[38494] = i[75];
  assign o[38495] = i[75];
  assign o[38496] = i[75];
  assign o[38497] = i[75];
  assign o[38498] = i[75];
  assign o[38499] = i[75];
  assign o[38500] = i[75];
  assign o[38501] = i[75];
  assign o[38502] = i[75];
  assign o[38503] = i[75];
  assign o[38504] = i[75];
  assign o[38505] = i[75];
  assign o[38506] = i[75];
  assign o[38507] = i[75];
  assign o[38508] = i[75];
  assign o[38509] = i[75];
  assign o[38510] = i[75];
  assign o[38511] = i[75];
  assign o[38512] = i[75];
  assign o[38513] = i[75];
  assign o[38514] = i[75];
  assign o[38515] = i[75];
  assign o[38516] = i[75];
  assign o[38517] = i[75];
  assign o[38518] = i[75];
  assign o[38519] = i[75];
  assign o[38520] = i[75];
  assign o[38521] = i[75];
  assign o[38522] = i[75];
  assign o[38523] = i[75];
  assign o[38524] = i[75];
  assign o[38525] = i[75];
  assign o[38526] = i[75];
  assign o[38527] = i[75];
  assign o[38528] = i[75];
  assign o[38529] = i[75];
  assign o[38530] = i[75];
  assign o[38531] = i[75];
  assign o[38532] = i[75];
  assign o[38533] = i[75];
  assign o[38534] = i[75];
  assign o[38535] = i[75];
  assign o[38536] = i[75];
  assign o[38537] = i[75];
  assign o[38538] = i[75];
  assign o[38539] = i[75];
  assign o[38540] = i[75];
  assign o[38541] = i[75];
  assign o[38542] = i[75];
  assign o[38543] = i[75];
  assign o[38544] = i[75];
  assign o[38545] = i[75];
  assign o[38546] = i[75];
  assign o[38547] = i[75];
  assign o[38548] = i[75];
  assign o[38549] = i[75];
  assign o[38550] = i[75];
  assign o[38551] = i[75];
  assign o[38552] = i[75];
  assign o[38553] = i[75];
  assign o[38554] = i[75];
  assign o[38555] = i[75];
  assign o[38556] = i[75];
  assign o[38557] = i[75];
  assign o[38558] = i[75];
  assign o[38559] = i[75];
  assign o[38560] = i[75];
  assign o[38561] = i[75];
  assign o[38562] = i[75];
  assign o[38563] = i[75];
  assign o[38564] = i[75];
  assign o[38565] = i[75];
  assign o[38566] = i[75];
  assign o[38567] = i[75];
  assign o[38568] = i[75];
  assign o[38569] = i[75];
  assign o[38570] = i[75];
  assign o[38571] = i[75];
  assign o[38572] = i[75];
  assign o[38573] = i[75];
  assign o[38574] = i[75];
  assign o[38575] = i[75];
  assign o[38576] = i[75];
  assign o[38577] = i[75];
  assign o[38578] = i[75];
  assign o[38579] = i[75];
  assign o[38580] = i[75];
  assign o[38581] = i[75];
  assign o[38582] = i[75];
  assign o[38583] = i[75];
  assign o[38584] = i[75];
  assign o[38585] = i[75];
  assign o[38586] = i[75];
  assign o[38587] = i[75];
  assign o[38588] = i[75];
  assign o[38589] = i[75];
  assign o[38590] = i[75];
  assign o[38591] = i[75];
  assign o[38592] = i[75];
  assign o[38593] = i[75];
  assign o[38594] = i[75];
  assign o[38595] = i[75];
  assign o[38596] = i[75];
  assign o[38597] = i[75];
  assign o[38598] = i[75];
  assign o[38599] = i[75];
  assign o[38600] = i[75];
  assign o[38601] = i[75];
  assign o[38602] = i[75];
  assign o[38603] = i[75];
  assign o[38604] = i[75];
  assign o[38605] = i[75];
  assign o[38606] = i[75];
  assign o[38607] = i[75];
  assign o[38608] = i[75];
  assign o[38609] = i[75];
  assign o[38610] = i[75];
  assign o[38611] = i[75];
  assign o[38612] = i[75];
  assign o[38613] = i[75];
  assign o[38614] = i[75];
  assign o[38615] = i[75];
  assign o[38616] = i[75];
  assign o[38617] = i[75];
  assign o[38618] = i[75];
  assign o[38619] = i[75];
  assign o[38620] = i[75];
  assign o[38621] = i[75];
  assign o[38622] = i[75];
  assign o[38623] = i[75];
  assign o[38624] = i[75];
  assign o[38625] = i[75];
  assign o[38626] = i[75];
  assign o[38627] = i[75];
  assign o[38628] = i[75];
  assign o[38629] = i[75];
  assign o[38630] = i[75];
  assign o[38631] = i[75];
  assign o[38632] = i[75];
  assign o[38633] = i[75];
  assign o[38634] = i[75];
  assign o[38635] = i[75];
  assign o[38636] = i[75];
  assign o[38637] = i[75];
  assign o[38638] = i[75];
  assign o[38639] = i[75];
  assign o[38640] = i[75];
  assign o[38641] = i[75];
  assign o[38642] = i[75];
  assign o[38643] = i[75];
  assign o[38644] = i[75];
  assign o[38645] = i[75];
  assign o[38646] = i[75];
  assign o[38647] = i[75];
  assign o[38648] = i[75];
  assign o[38649] = i[75];
  assign o[38650] = i[75];
  assign o[38651] = i[75];
  assign o[38652] = i[75];
  assign o[38653] = i[75];
  assign o[38654] = i[75];
  assign o[38655] = i[75];
  assign o[38656] = i[75];
  assign o[38657] = i[75];
  assign o[38658] = i[75];
  assign o[38659] = i[75];
  assign o[38660] = i[75];
  assign o[38661] = i[75];
  assign o[38662] = i[75];
  assign o[38663] = i[75];
  assign o[38664] = i[75];
  assign o[38665] = i[75];
  assign o[38666] = i[75];
  assign o[38667] = i[75];
  assign o[38668] = i[75];
  assign o[38669] = i[75];
  assign o[38670] = i[75];
  assign o[38671] = i[75];
  assign o[38672] = i[75];
  assign o[38673] = i[75];
  assign o[38674] = i[75];
  assign o[38675] = i[75];
  assign o[38676] = i[75];
  assign o[38677] = i[75];
  assign o[38678] = i[75];
  assign o[38679] = i[75];
  assign o[38680] = i[75];
  assign o[38681] = i[75];
  assign o[38682] = i[75];
  assign o[38683] = i[75];
  assign o[38684] = i[75];
  assign o[38685] = i[75];
  assign o[38686] = i[75];
  assign o[38687] = i[75];
  assign o[38688] = i[75];
  assign o[38689] = i[75];
  assign o[38690] = i[75];
  assign o[38691] = i[75];
  assign o[38692] = i[75];
  assign o[38693] = i[75];
  assign o[38694] = i[75];
  assign o[38695] = i[75];
  assign o[38696] = i[75];
  assign o[38697] = i[75];
  assign o[38698] = i[75];
  assign o[38699] = i[75];
  assign o[38700] = i[75];
  assign o[38701] = i[75];
  assign o[38702] = i[75];
  assign o[38703] = i[75];
  assign o[38704] = i[75];
  assign o[38705] = i[75];
  assign o[38706] = i[75];
  assign o[38707] = i[75];
  assign o[38708] = i[75];
  assign o[38709] = i[75];
  assign o[38710] = i[75];
  assign o[38711] = i[75];
  assign o[38712] = i[75];
  assign o[38713] = i[75];
  assign o[38714] = i[75];
  assign o[38715] = i[75];
  assign o[38716] = i[75];
  assign o[38717] = i[75];
  assign o[38718] = i[75];
  assign o[38719] = i[75];
  assign o[38720] = i[75];
  assign o[38721] = i[75];
  assign o[38722] = i[75];
  assign o[38723] = i[75];
  assign o[38724] = i[75];
  assign o[38725] = i[75];
  assign o[38726] = i[75];
  assign o[38727] = i[75];
  assign o[38728] = i[75];
  assign o[38729] = i[75];
  assign o[38730] = i[75];
  assign o[38731] = i[75];
  assign o[38732] = i[75];
  assign o[38733] = i[75];
  assign o[38734] = i[75];
  assign o[38735] = i[75];
  assign o[38736] = i[75];
  assign o[38737] = i[75];
  assign o[38738] = i[75];
  assign o[38739] = i[75];
  assign o[38740] = i[75];
  assign o[38741] = i[75];
  assign o[38742] = i[75];
  assign o[38743] = i[75];
  assign o[38744] = i[75];
  assign o[38745] = i[75];
  assign o[38746] = i[75];
  assign o[38747] = i[75];
  assign o[38748] = i[75];
  assign o[38749] = i[75];
  assign o[38750] = i[75];
  assign o[38751] = i[75];
  assign o[38752] = i[75];
  assign o[38753] = i[75];
  assign o[38754] = i[75];
  assign o[38755] = i[75];
  assign o[38756] = i[75];
  assign o[38757] = i[75];
  assign o[38758] = i[75];
  assign o[38759] = i[75];
  assign o[38760] = i[75];
  assign o[38761] = i[75];
  assign o[38762] = i[75];
  assign o[38763] = i[75];
  assign o[38764] = i[75];
  assign o[38765] = i[75];
  assign o[38766] = i[75];
  assign o[38767] = i[75];
  assign o[38768] = i[75];
  assign o[38769] = i[75];
  assign o[38770] = i[75];
  assign o[38771] = i[75];
  assign o[38772] = i[75];
  assign o[38773] = i[75];
  assign o[38774] = i[75];
  assign o[38775] = i[75];
  assign o[38776] = i[75];
  assign o[38777] = i[75];
  assign o[38778] = i[75];
  assign o[38779] = i[75];
  assign o[38780] = i[75];
  assign o[38781] = i[75];
  assign o[38782] = i[75];
  assign o[38783] = i[75];
  assign o[38784] = i[75];
  assign o[38785] = i[75];
  assign o[38786] = i[75];
  assign o[38787] = i[75];
  assign o[38788] = i[75];
  assign o[38789] = i[75];
  assign o[38790] = i[75];
  assign o[38791] = i[75];
  assign o[38792] = i[75];
  assign o[38793] = i[75];
  assign o[38794] = i[75];
  assign o[38795] = i[75];
  assign o[38796] = i[75];
  assign o[38797] = i[75];
  assign o[38798] = i[75];
  assign o[38799] = i[75];
  assign o[38800] = i[75];
  assign o[38801] = i[75];
  assign o[38802] = i[75];
  assign o[38803] = i[75];
  assign o[38804] = i[75];
  assign o[38805] = i[75];
  assign o[38806] = i[75];
  assign o[38807] = i[75];
  assign o[38808] = i[75];
  assign o[38809] = i[75];
  assign o[38810] = i[75];
  assign o[38811] = i[75];
  assign o[38812] = i[75];
  assign o[38813] = i[75];
  assign o[38814] = i[75];
  assign o[38815] = i[75];
  assign o[38816] = i[75];
  assign o[38817] = i[75];
  assign o[38818] = i[75];
  assign o[38819] = i[75];
  assign o[38820] = i[75];
  assign o[38821] = i[75];
  assign o[38822] = i[75];
  assign o[38823] = i[75];
  assign o[38824] = i[75];
  assign o[38825] = i[75];
  assign o[38826] = i[75];
  assign o[38827] = i[75];
  assign o[38828] = i[75];
  assign o[38829] = i[75];
  assign o[38830] = i[75];
  assign o[38831] = i[75];
  assign o[38832] = i[75];
  assign o[38833] = i[75];
  assign o[38834] = i[75];
  assign o[38835] = i[75];
  assign o[38836] = i[75];
  assign o[38837] = i[75];
  assign o[38838] = i[75];
  assign o[38839] = i[75];
  assign o[38840] = i[75];
  assign o[38841] = i[75];
  assign o[38842] = i[75];
  assign o[38843] = i[75];
  assign o[38844] = i[75];
  assign o[38845] = i[75];
  assign o[38846] = i[75];
  assign o[38847] = i[75];
  assign o[38848] = i[75];
  assign o[38849] = i[75];
  assign o[38850] = i[75];
  assign o[38851] = i[75];
  assign o[38852] = i[75];
  assign o[38853] = i[75];
  assign o[38854] = i[75];
  assign o[38855] = i[75];
  assign o[38856] = i[75];
  assign o[38857] = i[75];
  assign o[38858] = i[75];
  assign o[38859] = i[75];
  assign o[38860] = i[75];
  assign o[38861] = i[75];
  assign o[38862] = i[75];
  assign o[38863] = i[75];
  assign o[38864] = i[75];
  assign o[38865] = i[75];
  assign o[38866] = i[75];
  assign o[38867] = i[75];
  assign o[38868] = i[75];
  assign o[38869] = i[75];
  assign o[38870] = i[75];
  assign o[38871] = i[75];
  assign o[38872] = i[75];
  assign o[38873] = i[75];
  assign o[38874] = i[75];
  assign o[38875] = i[75];
  assign o[38876] = i[75];
  assign o[38877] = i[75];
  assign o[38878] = i[75];
  assign o[38879] = i[75];
  assign o[38880] = i[75];
  assign o[38881] = i[75];
  assign o[38882] = i[75];
  assign o[38883] = i[75];
  assign o[38884] = i[75];
  assign o[38885] = i[75];
  assign o[38886] = i[75];
  assign o[38887] = i[75];
  assign o[38888] = i[75];
  assign o[38889] = i[75];
  assign o[38890] = i[75];
  assign o[38891] = i[75];
  assign o[38892] = i[75];
  assign o[38893] = i[75];
  assign o[38894] = i[75];
  assign o[38895] = i[75];
  assign o[38896] = i[75];
  assign o[38897] = i[75];
  assign o[38898] = i[75];
  assign o[38899] = i[75];
  assign o[38900] = i[75];
  assign o[38901] = i[75];
  assign o[38902] = i[75];
  assign o[38903] = i[75];
  assign o[38904] = i[75];
  assign o[38905] = i[75];
  assign o[38906] = i[75];
  assign o[38907] = i[75];
  assign o[38908] = i[75];
  assign o[38909] = i[75];
  assign o[38910] = i[75];
  assign o[38911] = i[75];
  assign o[37888] = i[74];
  assign o[37889] = i[74];
  assign o[37890] = i[74];
  assign o[37891] = i[74];
  assign o[37892] = i[74];
  assign o[37893] = i[74];
  assign o[37894] = i[74];
  assign o[37895] = i[74];
  assign o[37896] = i[74];
  assign o[37897] = i[74];
  assign o[37898] = i[74];
  assign o[37899] = i[74];
  assign o[37900] = i[74];
  assign o[37901] = i[74];
  assign o[37902] = i[74];
  assign o[37903] = i[74];
  assign o[37904] = i[74];
  assign o[37905] = i[74];
  assign o[37906] = i[74];
  assign o[37907] = i[74];
  assign o[37908] = i[74];
  assign o[37909] = i[74];
  assign o[37910] = i[74];
  assign o[37911] = i[74];
  assign o[37912] = i[74];
  assign o[37913] = i[74];
  assign o[37914] = i[74];
  assign o[37915] = i[74];
  assign o[37916] = i[74];
  assign o[37917] = i[74];
  assign o[37918] = i[74];
  assign o[37919] = i[74];
  assign o[37920] = i[74];
  assign o[37921] = i[74];
  assign o[37922] = i[74];
  assign o[37923] = i[74];
  assign o[37924] = i[74];
  assign o[37925] = i[74];
  assign o[37926] = i[74];
  assign o[37927] = i[74];
  assign o[37928] = i[74];
  assign o[37929] = i[74];
  assign o[37930] = i[74];
  assign o[37931] = i[74];
  assign o[37932] = i[74];
  assign o[37933] = i[74];
  assign o[37934] = i[74];
  assign o[37935] = i[74];
  assign o[37936] = i[74];
  assign o[37937] = i[74];
  assign o[37938] = i[74];
  assign o[37939] = i[74];
  assign o[37940] = i[74];
  assign o[37941] = i[74];
  assign o[37942] = i[74];
  assign o[37943] = i[74];
  assign o[37944] = i[74];
  assign o[37945] = i[74];
  assign o[37946] = i[74];
  assign o[37947] = i[74];
  assign o[37948] = i[74];
  assign o[37949] = i[74];
  assign o[37950] = i[74];
  assign o[37951] = i[74];
  assign o[37952] = i[74];
  assign o[37953] = i[74];
  assign o[37954] = i[74];
  assign o[37955] = i[74];
  assign o[37956] = i[74];
  assign o[37957] = i[74];
  assign o[37958] = i[74];
  assign o[37959] = i[74];
  assign o[37960] = i[74];
  assign o[37961] = i[74];
  assign o[37962] = i[74];
  assign o[37963] = i[74];
  assign o[37964] = i[74];
  assign o[37965] = i[74];
  assign o[37966] = i[74];
  assign o[37967] = i[74];
  assign o[37968] = i[74];
  assign o[37969] = i[74];
  assign o[37970] = i[74];
  assign o[37971] = i[74];
  assign o[37972] = i[74];
  assign o[37973] = i[74];
  assign o[37974] = i[74];
  assign o[37975] = i[74];
  assign o[37976] = i[74];
  assign o[37977] = i[74];
  assign o[37978] = i[74];
  assign o[37979] = i[74];
  assign o[37980] = i[74];
  assign o[37981] = i[74];
  assign o[37982] = i[74];
  assign o[37983] = i[74];
  assign o[37984] = i[74];
  assign o[37985] = i[74];
  assign o[37986] = i[74];
  assign o[37987] = i[74];
  assign o[37988] = i[74];
  assign o[37989] = i[74];
  assign o[37990] = i[74];
  assign o[37991] = i[74];
  assign o[37992] = i[74];
  assign o[37993] = i[74];
  assign o[37994] = i[74];
  assign o[37995] = i[74];
  assign o[37996] = i[74];
  assign o[37997] = i[74];
  assign o[37998] = i[74];
  assign o[37999] = i[74];
  assign o[38000] = i[74];
  assign o[38001] = i[74];
  assign o[38002] = i[74];
  assign o[38003] = i[74];
  assign o[38004] = i[74];
  assign o[38005] = i[74];
  assign o[38006] = i[74];
  assign o[38007] = i[74];
  assign o[38008] = i[74];
  assign o[38009] = i[74];
  assign o[38010] = i[74];
  assign o[38011] = i[74];
  assign o[38012] = i[74];
  assign o[38013] = i[74];
  assign o[38014] = i[74];
  assign o[38015] = i[74];
  assign o[38016] = i[74];
  assign o[38017] = i[74];
  assign o[38018] = i[74];
  assign o[38019] = i[74];
  assign o[38020] = i[74];
  assign o[38021] = i[74];
  assign o[38022] = i[74];
  assign o[38023] = i[74];
  assign o[38024] = i[74];
  assign o[38025] = i[74];
  assign o[38026] = i[74];
  assign o[38027] = i[74];
  assign o[38028] = i[74];
  assign o[38029] = i[74];
  assign o[38030] = i[74];
  assign o[38031] = i[74];
  assign o[38032] = i[74];
  assign o[38033] = i[74];
  assign o[38034] = i[74];
  assign o[38035] = i[74];
  assign o[38036] = i[74];
  assign o[38037] = i[74];
  assign o[38038] = i[74];
  assign o[38039] = i[74];
  assign o[38040] = i[74];
  assign o[38041] = i[74];
  assign o[38042] = i[74];
  assign o[38043] = i[74];
  assign o[38044] = i[74];
  assign o[38045] = i[74];
  assign o[38046] = i[74];
  assign o[38047] = i[74];
  assign o[38048] = i[74];
  assign o[38049] = i[74];
  assign o[38050] = i[74];
  assign o[38051] = i[74];
  assign o[38052] = i[74];
  assign o[38053] = i[74];
  assign o[38054] = i[74];
  assign o[38055] = i[74];
  assign o[38056] = i[74];
  assign o[38057] = i[74];
  assign o[38058] = i[74];
  assign o[38059] = i[74];
  assign o[38060] = i[74];
  assign o[38061] = i[74];
  assign o[38062] = i[74];
  assign o[38063] = i[74];
  assign o[38064] = i[74];
  assign o[38065] = i[74];
  assign o[38066] = i[74];
  assign o[38067] = i[74];
  assign o[38068] = i[74];
  assign o[38069] = i[74];
  assign o[38070] = i[74];
  assign o[38071] = i[74];
  assign o[38072] = i[74];
  assign o[38073] = i[74];
  assign o[38074] = i[74];
  assign o[38075] = i[74];
  assign o[38076] = i[74];
  assign o[38077] = i[74];
  assign o[38078] = i[74];
  assign o[38079] = i[74];
  assign o[38080] = i[74];
  assign o[38081] = i[74];
  assign o[38082] = i[74];
  assign o[38083] = i[74];
  assign o[38084] = i[74];
  assign o[38085] = i[74];
  assign o[38086] = i[74];
  assign o[38087] = i[74];
  assign o[38088] = i[74];
  assign o[38089] = i[74];
  assign o[38090] = i[74];
  assign o[38091] = i[74];
  assign o[38092] = i[74];
  assign o[38093] = i[74];
  assign o[38094] = i[74];
  assign o[38095] = i[74];
  assign o[38096] = i[74];
  assign o[38097] = i[74];
  assign o[38098] = i[74];
  assign o[38099] = i[74];
  assign o[38100] = i[74];
  assign o[38101] = i[74];
  assign o[38102] = i[74];
  assign o[38103] = i[74];
  assign o[38104] = i[74];
  assign o[38105] = i[74];
  assign o[38106] = i[74];
  assign o[38107] = i[74];
  assign o[38108] = i[74];
  assign o[38109] = i[74];
  assign o[38110] = i[74];
  assign o[38111] = i[74];
  assign o[38112] = i[74];
  assign o[38113] = i[74];
  assign o[38114] = i[74];
  assign o[38115] = i[74];
  assign o[38116] = i[74];
  assign o[38117] = i[74];
  assign o[38118] = i[74];
  assign o[38119] = i[74];
  assign o[38120] = i[74];
  assign o[38121] = i[74];
  assign o[38122] = i[74];
  assign o[38123] = i[74];
  assign o[38124] = i[74];
  assign o[38125] = i[74];
  assign o[38126] = i[74];
  assign o[38127] = i[74];
  assign o[38128] = i[74];
  assign o[38129] = i[74];
  assign o[38130] = i[74];
  assign o[38131] = i[74];
  assign o[38132] = i[74];
  assign o[38133] = i[74];
  assign o[38134] = i[74];
  assign o[38135] = i[74];
  assign o[38136] = i[74];
  assign o[38137] = i[74];
  assign o[38138] = i[74];
  assign o[38139] = i[74];
  assign o[38140] = i[74];
  assign o[38141] = i[74];
  assign o[38142] = i[74];
  assign o[38143] = i[74];
  assign o[38144] = i[74];
  assign o[38145] = i[74];
  assign o[38146] = i[74];
  assign o[38147] = i[74];
  assign o[38148] = i[74];
  assign o[38149] = i[74];
  assign o[38150] = i[74];
  assign o[38151] = i[74];
  assign o[38152] = i[74];
  assign o[38153] = i[74];
  assign o[38154] = i[74];
  assign o[38155] = i[74];
  assign o[38156] = i[74];
  assign o[38157] = i[74];
  assign o[38158] = i[74];
  assign o[38159] = i[74];
  assign o[38160] = i[74];
  assign o[38161] = i[74];
  assign o[38162] = i[74];
  assign o[38163] = i[74];
  assign o[38164] = i[74];
  assign o[38165] = i[74];
  assign o[38166] = i[74];
  assign o[38167] = i[74];
  assign o[38168] = i[74];
  assign o[38169] = i[74];
  assign o[38170] = i[74];
  assign o[38171] = i[74];
  assign o[38172] = i[74];
  assign o[38173] = i[74];
  assign o[38174] = i[74];
  assign o[38175] = i[74];
  assign o[38176] = i[74];
  assign o[38177] = i[74];
  assign o[38178] = i[74];
  assign o[38179] = i[74];
  assign o[38180] = i[74];
  assign o[38181] = i[74];
  assign o[38182] = i[74];
  assign o[38183] = i[74];
  assign o[38184] = i[74];
  assign o[38185] = i[74];
  assign o[38186] = i[74];
  assign o[38187] = i[74];
  assign o[38188] = i[74];
  assign o[38189] = i[74];
  assign o[38190] = i[74];
  assign o[38191] = i[74];
  assign o[38192] = i[74];
  assign o[38193] = i[74];
  assign o[38194] = i[74];
  assign o[38195] = i[74];
  assign o[38196] = i[74];
  assign o[38197] = i[74];
  assign o[38198] = i[74];
  assign o[38199] = i[74];
  assign o[38200] = i[74];
  assign o[38201] = i[74];
  assign o[38202] = i[74];
  assign o[38203] = i[74];
  assign o[38204] = i[74];
  assign o[38205] = i[74];
  assign o[38206] = i[74];
  assign o[38207] = i[74];
  assign o[38208] = i[74];
  assign o[38209] = i[74];
  assign o[38210] = i[74];
  assign o[38211] = i[74];
  assign o[38212] = i[74];
  assign o[38213] = i[74];
  assign o[38214] = i[74];
  assign o[38215] = i[74];
  assign o[38216] = i[74];
  assign o[38217] = i[74];
  assign o[38218] = i[74];
  assign o[38219] = i[74];
  assign o[38220] = i[74];
  assign o[38221] = i[74];
  assign o[38222] = i[74];
  assign o[38223] = i[74];
  assign o[38224] = i[74];
  assign o[38225] = i[74];
  assign o[38226] = i[74];
  assign o[38227] = i[74];
  assign o[38228] = i[74];
  assign o[38229] = i[74];
  assign o[38230] = i[74];
  assign o[38231] = i[74];
  assign o[38232] = i[74];
  assign o[38233] = i[74];
  assign o[38234] = i[74];
  assign o[38235] = i[74];
  assign o[38236] = i[74];
  assign o[38237] = i[74];
  assign o[38238] = i[74];
  assign o[38239] = i[74];
  assign o[38240] = i[74];
  assign o[38241] = i[74];
  assign o[38242] = i[74];
  assign o[38243] = i[74];
  assign o[38244] = i[74];
  assign o[38245] = i[74];
  assign o[38246] = i[74];
  assign o[38247] = i[74];
  assign o[38248] = i[74];
  assign o[38249] = i[74];
  assign o[38250] = i[74];
  assign o[38251] = i[74];
  assign o[38252] = i[74];
  assign o[38253] = i[74];
  assign o[38254] = i[74];
  assign o[38255] = i[74];
  assign o[38256] = i[74];
  assign o[38257] = i[74];
  assign o[38258] = i[74];
  assign o[38259] = i[74];
  assign o[38260] = i[74];
  assign o[38261] = i[74];
  assign o[38262] = i[74];
  assign o[38263] = i[74];
  assign o[38264] = i[74];
  assign o[38265] = i[74];
  assign o[38266] = i[74];
  assign o[38267] = i[74];
  assign o[38268] = i[74];
  assign o[38269] = i[74];
  assign o[38270] = i[74];
  assign o[38271] = i[74];
  assign o[38272] = i[74];
  assign o[38273] = i[74];
  assign o[38274] = i[74];
  assign o[38275] = i[74];
  assign o[38276] = i[74];
  assign o[38277] = i[74];
  assign o[38278] = i[74];
  assign o[38279] = i[74];
  assign o[38280] = i[74];
  assign o[38281] = i[74];
  assign o[38282] = i[74];
  assign o[38283] = i[74];
  assign o[38284] = i[74];
  assign o[38285] = i[74];
  assign o[38286] = i[74];
  assign o[38287] = i[74];
  assign o[38288] = i[74];
  assign o[38289] = i[74];
  assign o[38290] = i[74];
  assign o[38291] = i[74];
  assign o[38292] = i[74];
  assign o[38293] = i[74];
  assign o[38294] = i[74];
  assign o[38295] = i[74];
  assign o[38296] = i[74];
  assign o[38297] = i[74];
  assign o[38298] = i[74];
  assign o[38299] = i[74];
  assign o[38300] = i[74];
  assign o[38301] = i[74];
  assign o[38302] = i[74];
  assign o[38303] = i[74];
  assign o[38304] = i[74];
  assign o[38305] = i[74];
  assign o[38306] = i[74];
  assign o[38307] = i[74];
  assign o[38308] = i[74];
  assign o[38309] = i[74];
  assign o[38310] = i[74];
  assign o[38311] = i[74];
  assign o[38312] = i[74];
  assign o[38313] = i[74];
  assign o[38314] = i[74];
  assign o[38315] = i[74];
  assign o[38316] = i[74];
  assign o[38317] = i[74];
  assign o[38318] = i[74];
  assign o[38319] = i[74];
  assign o[38320] = i[74];
  assign o[38321] = i[74];
  assign o[38322] = i[74];
  assign o[38323] = i[74];
  assign o[38324] = i[74];
  assign o[38325] = i[74];
  assign o[38326] = i[74];
  assign o[38327] = i[74];
  assign o[38328] = i[74];
  assign o[38329] = i[74];
  assign o[38330] = i[74];
  assign o[38331] = i[74];
  assign o[38332] = i[74];
  assign o[38333] = i[74];
  assign o[38334] = i[74];
  assign o[38335] = i[74];
  assign o[38336] = i[74];
  assign o[38337] = i[74];
  assign o[38338] = i[74];
  assign o[38339] = i[74];
  assign o[38340] = i[74];
  assign o[38341] = i[74];
  assign o[38342] = i[74];
  assign o[38343] = i[74];
  assign o[38344] = i[74];
  assign o[38345] = i[74];
  assign o[38346] = i[74];
  assign o[38347] = i[74];
  assign o[38348] = i[74];
  assign o[38349] = i[74];
  assign o[38350] = i[74];
  assign o[38351] = i[74];
  assign o[38352] = i[74];
  assign o[38353] = i[74];
  assign o[38354] = i[74];
  assign o[38355] = i[74];
  assign o[38356] = i[74];
  assign o[38357] = i[74];
  assign o[38358] = i[74];
  assign o[38359] = i[74];
  assign o[38360] = i[74];
  assign o[38361] = i[74];
  assign o[38362] = i[74];
  assign o[38363] = i[74];
  assign o[38364] = i[74];
  assign o[38365] = i[74];
  assign o[38366] = i[74];
  assign o[38367] = i[74];
  assign o[38368] = i[74];
  assign o[38369] = i[74];
  assign o[38370] = i[74];
  assign o[38371] = i[74];
  assign o[38372] = i[74];
  assign o[38373] = i[74];
  assign o[38374] = i[74];
  assign o[38375] = i[74];
  assign o[38376] = i[74];
  assign o[38377] = i[74];
  assign o[38378] = i[74];
  assign o[38379] = i[74];
  assign o[38380] = i[74];
  assign o[38381] = i[74];
  assign o[38382] = i[74];
  assign o[38383] = i[74];
  assign o[38384] = i[74];
  assign o[38385] = i[74];
  assign o[38386] = i[74];
  assign o[38387] = i[74];
  assign o[38388] = i[74];
  assign o[38389] = i[74];
  assign o[38390] = i[74];
  assign o[38391] = i[74];
  assign o[38392] = i[74];
  assign o[38393] = i[74];
  assign o[38394] = i[74];
  assign o[38395] = i[74];
  assign o[38396] = i[74];
  assign o[38397] = i[74];
  assign o[38398] = i[74];
  assign o[38399] = i[74];
  assign o[37376] = i[73];
  assign o[37377] = i[73];
  assign o[37378] = i[73];
  assign o[37379] = i[73];
  assign o[37380] = i[73];
  assign o[37381] = i[73];
  assign o[37382] = i[73];
  assign o[37383] = i[73];
  assign o[37384] = i[73];
  assign o[37385] = i[73];
  assign o[37386] = i[73];
  assign o[37387] = i[73];
  assign o[37388] = i[73];
  assign o[37389] = i[73];
  assign o[37390] = i[73];
  assign o[37391] = i[73];
  assign o[37392] = i[73];
  assign o[37393] = i[73];
  assign o[37394] = i[73];
  assign o[37395] = i[73];
  assign o[37396] = i[73];
  assign o[37397] = i[73];
  assign o[37398] = i[73];
  assign o[37399] = i[73];
  assign o[37400] = i[73];
  assign o[37401] = i[73];
  assign o[37402] = i[73];
  assign o[37403] = i[73];
  assign o[37404] = i[73];
  assign o[37405] = i[73];
  assign o[37406] = i[73];
  assign o[37407] = i[73];
  assign o[37408] = i[73];
  assign o[37409] = i[73];
  assign o[37410] = i[73];
  assign o[37411] = i[73];
  assign o[37412] = i[73];
  assign o[37413] = i[73];
  assign o[37414] = i[73];
  assign o[37415] = i[73];
  assign o[37416] = i[73];
  assign o[37417] = i[73];
  assign o[37418] = i[73];
  assign o[37419] = i[73];
  assign o[37420] = i[73];
  assign o[37421] = i[73];
  assign o[37422] = i[73];
  assign o[37423] = i[73];
  assign o[37424] = i[73];
  assign o[37425] = i[73];
  assign o[37426] = i[73];
  assign o[37427] = i[73];
  assign o[37428] = i[73];
  assign o[37429] = i[73];
  assign o[37430] = i[73];
  assign o[37431] = i[73];
  assign o[37432] = i[73];
  assign o[37433] = i[73];
  assign o[37434] = i[73];
  assign o[37435] = i[73];
  assign o[37436] = i[73];
  assign o[37437] = i[73];
  assign o[37438] = i[73];
  assign o[37439] = i[73];
  assign o[37440] = i[73];
  assign o[37441] = i[73];
  assign o[37442] = i[73];
  assign o[37443] = i[73];
  assign o[37444] = i[73];
  assign o[37445] = i[73];
  assign o[37446] = i[73];
  assign o[37447] = i[73];
  assign o[37448] = i[73];
  assign o[37449] = i[73];
  assign o[37450] = i[73];
  assign o[37451] = i[73];
  assign o[37452] = i[73];
  assign o[37453] = i[73];
  assign o[37454] = i[73];
  assign o[37455] = i[73];
  assign o[37456] = i[73];
  assign o[37457] = i[73];
  assign o[37458] = i[73];
  assign o[37459] = i[73];
  assign o[37460] = i[73];
  assign o[37461] = i[73];
  assign o[37462] = i[73];
  assign o[37463] = i[73];
  assign o[37464] = i[73];
  assign o[37465] = i[73];
  assign o[37466] = i[73];
  assign o[37467] = i[73];
  assign o[37468] = i[73];
  assign o[37469] = i[73];
  assign o[37470] = i[73];
  assign o[37471] = i[73];
  assign o[37472] = i[73];
  assign o[37473] = i[73];
  assign o[37474] = i[73];
  assign o[37475] = i[73];
  assign o[37476] = i[73];
  assign o[37477] = i[73];
  assign o[37478] = i[73];
  assign o[37479] = i[73];
  assign o[37480] = i[73];
  assign o[37481] = i[73];
  assign o[37482] = i[73];
  assign o[37483] = i[73];
  assign o[37484] = i[73];
  assign o[37485] = i[73];
  assign o[37486] = i[73];
  assign o[37487] = i[73];
  assign o[37488] = i[73];
  assign o[37489] = i[73];
  assign o[37490] = i[73];
  assign o[37491] = i[73];
  assign o[37492] = i[73];
  assign o[37493] = i[73];
  assign o[37494] = i[73];
  assign o[37495] = i[73];
  assign o[37496] = i[73];
  assign o[37497] = i[73];
  assign o[37498] = i[73];
  assign o[37499] = i[73];
  assign o[37500] = i[73];
  assign o[37501] = i[73];
  assign o[37502] = i[73];
  assign o[37503] = i[73];
  assign o[37504] = i[73];
  assign o[37505] = i[73];
  assign o[37506] = i[73];
  assign o[37507] = i[73];
  assign o[37508] = i[73];
  assign o[37509] = i[73];
  assign o[37510] = i[73];
  assign o[37511] = i[73];
  assign o[37512] = i[73];
  assign o[37513] = i[73];
  assign o[37514] = i[73];
  assign o[37515] = i[73];
  assign o[37516] = i[73];
  assign o[37517] = i[73];
  assign o[37518] = i[73];
  assign o[37519] = i[73];
  assign o[37520] = i[73];
  assign o[37521] = i[73];
  assign o[37522] = i[73];
  assign o[37523] = i[73];
  assign o[37524] = i[73];
  assign o[37525] = i[73];
  assign o[37526] = i[73];
  assign o[37527] = i[73];
  assign o[37528] = i[73];
  assign o[37529] = i[73];
  assign o[37530] = i[73];
  assign o[37531] = i[73];
  assign o[37532] = i[73];
  assign o[37533] = i[73];
  assign o[37534] = i[73];
  assign o[37535] = i[73];
  assign o[37536] = i[73];
  assign o[37537] = i[73];
  assign o[37538] = i[73];
  assign o[37539] = i[73];
  assign o[37540] = i[73];
  assign o[37541] = i[73];
  assign o[37542] = i[73];
  assign o[37543] = i[73];
  assign o[37544] = i[73];
  assign o[37545] = i[73];
  assign o[37546] = i[73];
  assign o[37547] = i[73];
  assign o[37548] = i[73];
  assign o[37549] = i[73];
  assign o[37550] = i[73];
  assign o[37551] = i[73];
  assign o[37552] = i[73];
  assign o[37553] = i[73];
  assign o[37554] = i[73];
  assign o[37555] = i[73];
  assign o[37556] = i[73];
  assign o[37557] = i[73];
  assign o[37558] = i[73];
  assign o[37559] = i[73];
  assign o[37560] = i[73];
  assign o[37561] = i[73];
  assign o[37562] = i[73];
  assign o[37563] = i[73];
  assign o[37564] = i[73];
  assign o[37565] = i[73];
  assign o[37566] = i[73];
  assign o[37567] = i[73];
  assign o[37568] = i[73];
  assign o[37569] = i[73];
  assign o[37570] = i[73];
  assign o[37571] = i[73];
  assign o[37572] = i[73];
  assign o[37573] = i[73];
  assign o[37574] = i[73];
  assign o[37575] = i[73];
  assign o[37576] = i[73];
  assign o[37577] = i[73];
  assign o[37578] = i[73];
  assign o[37579] = i[73];
  assign o[37580] = i[73];
  assign o[37581] = i[73];
  assign o[37582] = i[73];
  assign o[37583] = i[73];
  assign o[37584] = i[73];
  assign o[37585] = i[73];
  assign o[37586] = i[73];
  assign o[37587] = i[73];
  assign o[37588] = i[73];
  assign o[37589] = i[73];
  assign o[37590] = i[73];
  assign o[37591] = i[73];
  assign o[37592] = i[73];
  assign o[37593] = i[73];
  assign o[37594] = i[73];
  assign o[37595] = i[73];
  assign o[37596] = i[73];
  assign o[37597] = i[73];
  assign o[37598] = i[73];
  assign o[37599] = i[73];
  assign o[37600] = i[73];
  assign o[37601] = i[73];
  assign o[37602] = i[73];
  assign o[37603] = i[73];
  assign o[37604] = i[73];
  assign o[37605] = i[73];
  assign o[37606] = i[73];
  assign o[37607] = i[73];
  assign o[37608] = i[73];
  assign o[37609] = i[73];
  assign o[37610] = i[73];
  assign o[37611] = i[73];
  assign o[37612] = i[73];
  assign o[37613] = i[73];
  assign o[37614] = i[73];
  assign o[37615] = i[73];
  assign o[37616] = i[73];
  assign o[37617] = i[73];
  assign o[37618] = i[73];
  assign o[37619] = i[73];
  assign o[37620] = i[73];
  assign o[37621] = i[73];
  assign o[37622] = i[73];
  assign o[37623] = i[73];
  assign o[37624] = i[73];
  assign o[37625] = i[73];
  assign o[37626] = i[73];
  assign o[37627] = i[73];
  assign o[37628] = i[73];
  assign o[37629] = i[73];
  assign o[37630] = i[73];
  assign o[37631] = i[73];
  assign o[37632] = i[73];
  assign o[37633] = i[73];
  assign o[37634] = i[73];
  assign o[37635] = i[73];
  assign o[37636] = i[73];
  assign o[37637] = i[73];
  assign o[37638] = i[73];
  assign o[37639] = i[73];
  assign o[37640] = i[73];
  assign o[37641] = i[73];
  assign o[37642] = i[73];
  assign o[37643] = i[73];
  assign o[37644] = i[73];
  assign o[37645] = i[73];
  assign o[37646] = i[73];
  assign o[37647] = i[73];
  assign o[37648] = i[73];
  assign o[37649] = i[73];
  assign o[37650] = i[73];
  assign o[37651] = i[73];
  assign o[37652] = i[73];
  assign o[37653] = i[73];
  assign o[37654] = i[73];
  assign o[37655] = i[73];
  assign o[37656] = i[73];
  assign o[37657] = i[73];
  assign o[37658] = i[73];
  assign o[37659] = i[73];
  assign o[37660] = i[73];
  assign o[37661] = i[73];
  assign o[37662] = i[73];
  assign o[37663] = i[73];
  assign o[37664] = i[73];
  assign o[37665] = i[73];
  assign o[37666] = i[73];
  assign o[37667] = i[73];
  assign o[37668] = i[73];
  assign o[37669] = i[73];
  assign o[37670] = i[73];
  assign o[37671] = i[73];
  assign o[37672] = i[73];
  assign o[37673] = i[73];
  assign o[37674] = i[73];
  assign o[37675] = i[73];
  assign o[37676] = i[73];
  assign o[37677] = i[73];
  assign o[37678] = i[73];
  assign o[37679] = i[73];
  assign o[37680] = i[73];
  assign o[37681] = i[73];
  assign o[37682] = i[73];
  assign o[37683] = i[73];
  assign o[37684] = i[73];
  assign o[37685] = i[73];
  assign o[37686] = i[73];
  assign o[37687] = i[73];
  assign o[37688] = i[73];
  assign o[37689] = i[73];
  assign o[37690] = i[73];
  assign o[37691] = i[73];
  assign o[37692] = i[73];
  assign o[37693] = i[73];
  assign o[37694] = i[73];
  assign o[37695] = i[73];
  assign o[37696] = i[73];
  assign o[37697] = i[73];
  assign o[37698] = i[73];
  assign o[37699] = i[73];
  assign o[37700] = i[73];
  assign o[37701] = i[73];
  assign o[37702] = i[73];
  assign o[37703] = i[73];
  assign o[37704] = i[73];
  assign o[37705] = i[73];
  assign o[37706] = i[73];
  assign o[37707] = i[73];
  assign o[37708] = i[73];
  assign o[37709] = i[73];
  assign o[37710] = i[73];
  assign o[37711] = i[73];
  assign o[37712] = i[73];
  assign o[37713] = i[73];
  assign o[37714] = i[73];
  assign o[37715] = i[73];
  assign o[37716] = i[73];
  assign o[37717] = i[73];
  assign o[37718] = i[73];
  assign o[37719] = i[73];
  assign o[37720] = i[73];
  assign o[37721] = i[73];
  assign o[37722] = i[73];
  assign o[37723] = i[73];
  assign o[37724] = i[73];
  assign o[37725] = i[73];
  assign o[37726] = i[73];
  assign o[37727] = i[73];
  assign o[37728] = i[73];
  assign o[37729] = i[73];
  assign o[37730] = i[73];
  assign o[37731] = i[73];
  assign o[37732] = i[73];
  assign o[37733] = i[73];
  assign o[37734] = i[73];
  assign o[37735] = i[73];
  assign o[37736] = i[73];
  assign o[37737] = i[73];
  assign o[37738] = i[73];
  assign o[37739] = i[73];
  assign o[37740] = i[73];
  assign o[37741] = i[73];
  assign o[37742] = i[73];
  assign o[37743] = i[73];
  assign o[37744] = i[73];
  assign o[37745] = i[73];
  assign o[37746] = i[73];
  assign o[37747] = i[73];
  assign o[37748] = i[73];
  assign o[37749] = i[73];
  assign o[37750] = i[73];
  assign o[37751] = i[73];
  assign o[37752] = i[73];
  assign o[37753] = i[73];
  assign o[37754] = i[73];
  assign o[37755] = i[73];
  assign o[37756] = i[73];
  assign o[37757] = i[73];
  assign o[37758] = i[73];
  assign o[37759] = i[73];
  assign o[37760] = i[73];
  assign o[37761] = i[73];
  assign o[37762] = i[73];
  assign o[37763] = i[73];
  assign o[37764] = i[73];
  assign o[37765] = i[73];
  assign o[37766] = i[73];
  assign o[37767] = i[73];
  assign o[37768] = i[73];
  assign o[37769] = i[73];
  assign o[37770] = i[73];
  assign o[37771] = i[73];
  assign o[37772] = i[73];
  assign o[37773] = i[73];
  assign o[37774] = i[73];
  assign o[37775] = i[73];
  assign o[37776] = i[73];
  assign o[37777] = i[73];
  assign o[37778] = i[73];
  assign o[37779] = i[73];
  assign o[37780] = i[73];
  assign o[37781] = i[73];
  assign o[37782] = i[73];
  assign o[37783] = i[73];
  assign o[37784] = i[73];
  assign o[37785] = i[73];
  assign o[37786] = i[73];
  assign o[37787] = i[73];
  assign o[37788] = i[73];
  assign o[37789] = i[73];
  assign o[37790] = i[73];
  assign o[37791] = i[73];
  assign o[37792] = i[73];
  assign o[37793] = i[73];
  assign o[37794] = i[73];
  assign o[37795] = i[73];
  assign o[37796] = i[73];
  assign o[37797] = i[73];
  assign o[37798] = i[73];
  assign o[37799] = i[73];
  assign o[37800] = i[73];
  assign o[37801] = i[73];
  assign o[37802] = i[73];
  assign o[37803] = i[73];
  assign o[37804] = i[73];
  assign o[37805] = i[73];
  assign o[37806] = i[73];
  assign o[37807] = i[73];
  assign o[37808] = i[73];
  assign o[37809] = i[73];
  assign o[37810] = i[73];
  assign o[37811] = i[73];
  assign o[37812] = i[73];
  assign o[37813] = i[73];
  assign o[37814] = i[73];
  assign o[37815] = i[73];
  assign o[37816] = i[73];
  assign o[37817] = i[73];
  assign o[37818] = i[73];
  assign o[37819] = i[73];
  assign o[37820] = i[73];
  assign o[37821] = i[73];
  assign o[37822] = i[73];
  assign o[37823] = i[73];
  assign o[37824] = i[73];
  assign o[37825] = i[73];
  assign o[37826] = i[73];
  assign o[37827] = i[73];
  assign o[37828] = i[73];
  assign o[37829] = i[73];
  assign o[37830] = i[73];
  assign o[37831] = i[73];
  assign o[37832] = i[73];
  assign o[37833] = i[73];
  assign o[37834] = i[73];
  assign o[37835] = i[73];
  assign o[37836] = i[73];
  assign o[37837] = i[73];
  assign o[37838] = i[73];
  assign o[37839] = i[73];
  assign o[37840] = i[73];
  assign o[37841] = i[73];
  assign o[37842] = i[73];
  assign o[37843] = i[73];
  assign o[37844] = i[73];
  assign o[37845] = i[73];
  assign o[37846] = i[73];
  assign o[37847] = i[73];
  assign o[37848] = i[73];
  assign o[37849] = i[73];
  assign o[37850] = i[73];
  assign o[37851] = i[73];
  assign o[37852] = i[73];
  assign o[37853] = i[73];
  assign o[37854] = i[73];
  assign o[37855] = i[73];
  assign o[37856] = i[73];
  assign o[37857] = i[73];
  assign o[37858] = i[73];
  assign o[37859] = i[73];
  assign o[37860] = i[73];
  assign o[37861] = i[73];
  assign o[37862] = i[73];
  assign o[37863] = i[73];
  assign o[37864] = i[73];
  assign o[37865] = i[73];
  assign o[37866] = i[73];
  assign o[37867] = i[73];
  assign o[37868] = i[73];
  assign o[37869] = i[73];
  assign o[37870] = i[73];
  assign o[37871] = i[73];
  assign o[37872] = i[73];
  assign o[37873] = i[73];
  assign o[37874] = i[73];
  assign o[37875] = i[73];
  assign o[37876] = i[73];
  assign o[37877] = i[73];
  assign o[37878] = i[73];
  assign o[37879] = i[73];
  assign o[37880] = i[73];
  assign o[37881] = i[73];
  assign o[37882] = i[73];
  assign o[37883] = i[73];
  assign o[37884] = i[73];
  assign o[37885] = i[73];
  assign o[37886] = i[73];
  assign o[37887] = i[73];
  assign o[36864] = i[72];
  assign o[36865] = i[72];
  assign o[36866] = i[72];
  assign o[36867] = i[72];
  assign o[36868] = i[72];
  assign o[36869] = i[72];
  assign o[36870] = i[72];
  assign o[36871] = i[72];
  assign o[36872] = i[72];
  assign o[36873] = i[72];
  assign o[36874] = i[72];
  assign o[36875] = i[72];
  assign o[36876] = i[72];
  assign o[36877] = i[72];
  assign o[36878] = i[72];
  assign o[36879] = i[72];
  assign o[36880] = i[72];
  assign o[36881] = i[72];
  assign o[36882] = i[72];
  assign o[36883] = i[72];
  assign o[36884] = i[72];
  assign o[36885] = i[72];
  assign o[36886] = i[72];
  assign o[36887] = i[72];
  assign o[36888] = i[72];
  assign o[36889] = i[72];
  assign o[36890] = i[72];
  assign o[36891] = i[72];
  assign o[36892] = i[72];
  assign o[36893] = i[72];
  assign o[36894] = i[72];
  assign o[36895] = i[72];
  assign o[36896] = i[72];
  assign o[36897] = i[72];
  assign o[36898] = i[72];
  assign o[36899] = i[72];
  assign o[36900] = i[72];
  assign o[36901] = i[72];
  assign o[36902] = i[72];
  assign o[36903] = i[72];
  assign o[36904] = i[72];
  assign o[36905] = i[72];
  assign o[36906] = i[72];
  assign o[36907] = i[72];
  assign o[36908] = i[72];
  assign o[36909] = i[72];
  assign o[36910] = i[72];
  assign o[36911] = i[72];
  assign o[36912] = i[72];
  assign o[36913] = i[72];
  assign o[36914] = i[72];
  assign o[36915] = i[72];
  assign o[36916] = i[72];
  assign o[36917] = i[72];
  assign o[36918] = i[72];
  assign o[36919] = i[72];
  assign o[36920] = i[72];
  assign o[36921] = i[72];
  assign o[36922] = i[72];
  assign o[36923] = i[72];
  assign o[36924] = i[72];
  assign o[36925] = i[72];
  assign o[36926] = i[72];
  assign o[36927] = i[72];
  assign o[36928] = i[72];
  assign o[36929] = i[72];
  assign o[36930] = i[72];
  assign o[36931] = i[72];
  assign o[36932] = i[72];
  assign o[36933] = i[72];
  assign o[36934] = i[72];
  assign o[36935] = i[72];
  assign o[36936] = i[72];
  assign o[36937] = i[72];
  assign o[36938] = i[72];
  assign o[36939] = i[72];
  assign o[36940] = i[72];
  assign o[36941] = i[72];
  assign o[36942] = i[72];
  assign o[36943] = i[72];
  assign o[36944] = i[72];
  assign o[36945] = i[72];
  assign o[36946] = i[72];
  assign o[36947] = i[72];
  assign o[36948] = i[72];
  assign o[36949] = i[72];
  assign o[36950] = i[72];
  assign o[36951] = i[72];
  assign o[36952] = i[72];
  assign o[36953] = i[72];
  assign o[36954] = i[72];
  assign o[36955] = i[72];
  assign o[36956] = i[72];
  assign o[36957] = i[72];
  assign o[36958] = i[72];
  assign o[36959] = i[72];
  assign o[36960] = i[72];
  assign o[36961] = i[72];
  assign o[36962] = i[72];
  assign o[36963] = i[72];
  assign o[36964] = i[72];
  assign o[36965] = i[72];
  assign o[36966] = i[72];
  assign o[36967] = i[72];
  assign o[36968] = i[72];
  assign o[36969] = i[72];
  assign o[36970] = i[72];
  assign o[36971] = i[72];
  assign o[36972] = i[72];
  assign o[36973] = i[72];
  assign o[36974] = i[72];
  assign o[36975] = i[72];
  assign o[36976] = i[72];
  assign o[36977] = i[72];
  assign o[36978] = i[72];
  assign o[36979] = i[72];
  assign o[36980] = i[72];
  assign o[36981] = i[72];
  assign o[36982] = i[72];
  assign o[36983] = i[72];
  assign o[36984] = i[72];
  assign o[36985] = i[72];
  assign o[36986] = i[72];
  assign o[36987] = i[72];
  assign o[36988] = i[72];
  assign o[36989] = i[72];
  assign o[36990] = i[72];
  assign o[36991] = i[72];
  assign o[36992] = i[72];
  assign o[36993] = i[72];
  assign o[36994] = i[72];
  assign o[36995] = i[72];
  assign o[36996] = i[72];
  assign o[36997] = i[72];
  assign o[36998] = i[72];
  assign o[36999] = i[72];
  assign o[37000] = i[72];
  assign o[37001] = i[72];
  assign o[37002] = i[72];
  assign o[37003] = i[72];
  assign o[37004] = i[72];
  assign o[37005] = i[72];
  assign o[37006] = i[72];
  assign o[37007] = i[72];
  assign o[37008] = i[72];
  assign o[37009] = i[72];
  assign o[37010] = i[72];
  assign o[37011] = i[72];
  assign o[37012] = i[72];
  assign o[37013] = i[72];
  assign o[37014] = i[72];
  assign o[37015] = i[72];
  assign o[37016] = i[72];
  assign o[37017] = i[72];
  assign o[37018] = i[72];
  assign o[37019] = i[72];
  assign o[37020] = i[72];
  assign o[37021] = i[72];
  assign o[37022] = i[72];
  assign o[37023] = i[72];
  assign o[37024] = i[72];
  assign o[37025] = i[72];
  assign o[37026] = i[72];
  assign o[37027] = i[72];
  assign o[37028] = i[72];
  assign o[37029] = i[72];
  assign o[37030] = i[72];
  assign o[37031] = i[72];
  assign o[37032] = i[72];
  assign o[37033] = i[72];
  assign o[37034] = i[72];
  assign o[37035] = i[72];
  assign o[37036] = i[72];
  assign o[37037] = i[72];
  assign o[37038] = i[72];
  assign o[37039] = i[72];
  assign o[37040] = i[72];
  assign o[37041] = i[72];
  assign o[37042] = i[72];
  assign o[37043] = i[72];
  assign o[37044] = i[72];
  assign o[37045] = i[72];
  assign o[37046] = i[72];
  assign o[37047] = i[72];
  assign o[37048] = i[72];
  assign o[37049] = i[72];
  assign o[37050] = i[72];
  assign o[37051] = i[72];
  assign o[37052] = i[72];
  assign o[37053] = i[72];
  assign o[37054] = i[72];
  assign o[37055] = i[72];
  assign o[37056] = i[72];
  assign o[37057] = i[72];
  assign o[37058] = i[72];
  assign o[37059] = i[72];
  assign o[37060] = i[72];
  assign o[37061] = i[72];
  assign o[37062] = i[72];
  assign o[37063] = i[72];
  assign o[37064] = i[72];
  assign o[37065] = i[72];
  assign o[37066] = i[72];
  assign o[37067] = i[72];
  assign o[37068] = i[72];
  assign o[37069] = i[72];
  assign o[37070] = i[72];
  assign o[37071] = i[72];
  assign o[37072] = i[72];
  assign o[37073] = i[72];
  assign o[37074] = i[72];
  assign o[37075] = i[72];
  assign o[37076] = i[72];
  assign o[37077] = i[72];
  assign o[37078] = i[72];
  assign o[37079] = i[72];
  assign o[37080] = i[72];
  assign o[37081] = i[72];
  assign o[37082] = i[72];
  assign o[37083] = i[72];
  assign o[37084] = i[72];
  assign o[37085] = i[72];
  assign o[37086] = i[72];
  assign o[37087] = i[72];
  assign o[37088] = i[72];
  assign o[37089] = i[72];
  assign o[37090] = i[72];
  assign o[37091] = i[72];
  assign o[37092] = i[72];
  assign o[37093] = i[72];
  assign o[37094] = i[72];
  assign o[37095] = i[72];
  assign o[37096] = i[72];
  assign o[37097] = i[72];
  assign o[37098] = i[72];
  assign o[37099] = i[72];
  assign o[37100] = i[72];
  assign o[37101] = i[72];
  assign o[37102] = i[72];
  assign o[37103] = i[72];
  assign o[37104] = i[72];
  assign o[37105] = i[72];
  assign o[37106] = i[72];
  assign o[37107] = i[72];
  assign o[37108] = i[72];
  assign o[37109] = i[72];
  assign o[37110] = i[72];
  assign o[37111] = i[72];
  assign o[37112] = i[72];
  assign o[37113] = i[72];
  assign o[37114] = i[72];
  assign o[37115] = i[72];
  assign o[37116] = i[72];
  assign o[37117] = i[72];
  assign o[37118] = i[72];
  assign o[37119] = i[72];
  assign o[37120] = i[72];
  assign o[37121] = i[72];
  assign o[37122] = i[72];
  assign o[37123] = i[72];
  assign o[37124] = i[72];
  assign o[37125] = i[72];
  assign o[37126] = i[72];
  assign o[37127] = i[72];
  assign o[37128] = i[72];
  assign o[37129] = i[72];
  assign o[37130] = i[72];
  assign o[37131] = i[72];
  assign o[37132] = i[72];
  assign o[37133] = i[72];
  assign o[37134] = i[72];
  assign o[37135] = i[72];
  assign o[37136] = i[72];
  assign o[37137] = i[72];
  assign o[37138] = i[72];
  assign o[37139] = i[72];
  assign o[37140] = i[72];
  assign o[37141] = i[72];
  assign o[37142] = i[72];
  assign o[37143] = i[72];
  assign o[37144] = i[72];
  assign o[37145] = i[72];
  assign o[37146] = i[72];
  assign o[37147] = i[72];
  assign o[37148] = i[72];
  assign o[37149] = i[72];
  assign o[37150] = i[72];
  assign o[37151] = i[72];
  assign o[37152] = i[72];
  assign o[37153] = i[72];
  assign o[37154] = i[72];
  assign o[37155] = i[72];
  assign o[37156] = i[72];
  assign o[37157] = i[72];
  assign o[37158] = i[72];
  assign o[37159] = i[72];
  assign o[37160] = i[72];
  assign o[37161] = i[72];
  assign o[37162] = i[72];
  assign o[37163] = i[72];
  assign o[37164] = i[72];
  assign o[37165] = i[72];
  assign o[37166] = i[72];
  assign o[37167] = i[72];
  assign o[37168] = i[72];
  assign o[37169] = i[72];
  assign o[37170] = i[72];
  assign o[37171] = i[72];
  assign o[37172] = i[72];
  assign o[37173] = i[72];
  assign o[37174] = i[72];
  assign o[37175] = i[72];
  assign o[37176] = i[72];
  assign o[37177] = i[72];
  assign o[37178] = i[72];
  assign o[37179] = i[72];
  assign o[37180] = i[72];
  assign o[37181] = i[72];
  assign o[37182] = i[72];
  assign o[37183] = i[72];
  assign o[37184] = i[72];
  assign o[37185] = i[72];
  assign o[37186] = i[72];
  assign o[37187] = i[72];
  assign o[37188] = i[72];
  assign o[37189] = i[72];
  assign o[37190] = i[72];
  assign o[37191] = i[72];
  assign o[37192] = i[72];
  assign o[37193] = i[72];
  assign o[37194] = i[72];
  assign o[37195] = i[72];
  assign o[37196] = i[72];
  assign o[37197] = i[72];
  assign o[37198] = i[72];
  assign o[37199] = i[72];
  assign o[37200] = i[72];
  assign o[37201] = i[72];
  assign o[37202] = i[72];
  assign o[37203] = i[72];
  assign o[37204] = i[72];
  assign o[37205] = i[72];
  assign o[37206] = i[72];
  assign o[37207] = i[72];
  assign o[37208] = i[72];
  assign o[37209] = i[72];
  assign o[37210] = i[72];
  assign o[37211] = i[72];
  assign o[37212] = i[72];
  assign o[37213] = i[72];
  assign o[37214] = i[72];
  assign o[37215] = i[72];
  assign o[37216] = i[72];
  assign o[37217] = i[72];
  assign o[37218] = i[72];
  assign o[37219] = i[72];
  assign o[37220] = i[72];
  assign o[37221] = i[72];
  assign o[37222] = i[72];
  assign o[37223] = i[72];
  assign o[37224] = i[72];
  assign o[37225] = i[72];
  assign o[37226] = i[72];
  assign o[37227] = i[72];
  assign o[37228] = i[72];
  assign o[37229] = i[72];
  assign o[37230] = i[72];
  assign o[37231] = i[72];
  assign o[37232] = i[72];
  assign o[37233] = i[72];
  assign o[37234] = i[72];
  assign o[37235] = i[72];
  assign o[37236] = i[72];
  assign o[37237] = i[72];
  assign o[37238] = i[72];
  assign o[37239] = i[72];
  assign o[37240] = i[72];
  assign o[37241] = i[72];
  assign o[37242] = i[72];
  assign o[37243] = i[72];
  assign o[37244] = i[72];
  assign o[37245] = i[72];
  assign o[37246] = i[72];
  assign o[37247] = i[72];
  assign o[37248] = i[72];
  assign o[37249] = i[72];
  assign o[37250] = i[72];
  assign o[37251] = i[72];
  assign o[37252] = i[72];
  assign o[37253] = i[72];
  assign o[37254] = i[72];
  assign o[37255] = i[72];
  assign o[37256] = i[72];
  assign o[37257] = i[72];
  assign o[37258] = i[72];
  assign o[37259] = i[72];
  assign o[37260] = i[72];
  assign o[37261] = i[72];
  assign o[37262] = i[72];
  assign o[37263] = i[72];
  assign o[37264] = i[72];
  assign o[37265] = i[72];
  assign o[37266] = i[72];
  assign o[37267] = i[72];
  assign o[37268] = i[72];
  assign o[37269] = i[72];
  assign o[37270] = i[72];
  assign o[37271] = i[72];
  assign o[37272] = i[72];
  assign o[37273] = i[72];
  assign o[37274] = i[72];
  assign o[37275] = i[72];
  assign o[37276] = i[72];
  assign o[37277] = i[72];
  assign o[37278] = i[72];
  assign o[37279] = i[72];
  assign o[37280] = i[72];
  assign o[37281] = i[72];
  assign o[37282] = i[72];
  assign o[37283] = i[72];
  assign o[37284] = i[72];
  assign o[37285] = i[72];
  assign o[37286] = i[72];
  assign o[37287] = i[72];
  assign o[37288] = i[72];
  assign o[37289] = i[72];
  assign o[37290] = i[72];
  assign o[37291] = i[72];
  assign o[37292] = i[72];
  assign o[37293] = i[72];
  assign o[37294] = i[72];
  assign o[37295] = i[72];
  assign o[37296] = i[72];
  assign o[37297] = i[72];
  assign o[37298] = i[72];
  assign o[37299] = i[72];
  assign o[37300] = i[72];
  assign o[37301] = i[72];
  assign o[37302] = i[72];
  assign o[37303] = i[72];
  assign o[37304] = i[72];
  assign o[37305] = i[72];
  assign o[37306] = i[72];
  assign o[37307] = i[72];
  assign o[37308] = i[72];
  assign o[37309] = i[72];
  assign o[37310] = i[72];
  assign o[37311] = i[72];
  assign o[37312] = i[72];
  assign o[37313] = i[72];
  assign o[37314] = i[72];
  assign o[37315] = i[72];
  assign o[37316] = i[72];
  assign o[37317] = i[72];
  assign o[37318] = i[72];
  assign o[37319] = i[72];
  assign o[37320] = i[72];
  assign o[37321] = i[72];
  assign o[37322] = i[72];
  assign o[37323] = i[72];
  assign o[37324] = i[72];
  assign o[37325] = i[72];
  assign o[37326] = i[72];
  assign o[37327] = i[72];
  assign o[37328] = i[72];
  assign o[37329] = i[72];
  assign o[37330] = i[72];
  assign o[37331] = i[72];
  assign o[37332] = i[72];
  assign o[37333] = i[72];
  assign o[37334] = i[72];
  assign o[37335] = i[72];
  assign o[37336] = i[72];
  assign o[37337] = i[72];
  assign o[37338] = i[72];
  assign o[37339] = i[72];
  assign o[37340] = i[72];
  assign o[37341] = i[72];
  assign o[37342] = i[72];
  assign o[37343] = i[72];
  assign o[37344] = i[72];
  assign o[37345] = i[72];
  assign o[37346] = i[72];
  assign o[37347] = i[72];
  assign o[37348] = i[72];
  assign o[37349] = i[72];
  assign o[37350] = i[72];
  assign o[37351] = i[72];
  assign o[37352] = i[72];
  assign o[37353] = i[72];
  assign o[37354] = i[72];
  assign o[37355] = i[72];
  assign o[37356] = i[72];
  assign o[37357] = i[72];
  assign o[37358] = i[72];
  assign o[37359] = i[72];
  assign o[37360] = i[72];
  assign o[37361] = i[72];
  assign o[37362] = i[72];
  assign o[37363] = i[72];
  assign o[37364] = i[72];
  assign o[37365] = i[72];
  assign o[37366] = i[72];
  assign o[37367] = i[72];
  assign o[37368] = i[72];
  assign o[37369] = i[72];
  assign o[37370] = i[72];
  assign o[37371] = i[72];
  assign o[37372] = i[72];
  assign o[37373] = i[72];
  assign o[37374] = i[72];
  assign o[37375] = i[72];
  assign o[36352] = i[71];
  assign o[36353] = i[71];
  assign o[36354] = i[71];
  assign o[36355] = i[71];
  assign o[36356] = i[71];
  assign o[36357] = i[71];
  assign o[36358] = i[71];
  assign o[36359] = i[71];
  assign o[36360] = i[71];
  assign o[36361] = i[71];
  assign o[36362] = i[71];
  assign o[36363] = i[71];
  assign o[36364] = i[71];
  assign o[36365] = i[71];
  assign o[36366] = i[71];
  assign o[36367] = i[71];
  assign o[36368] = i[71];
  assign o[36369] = i[71];
  assign o[36370] = i[71];
  assign o[36371] = i[71];
  assign o[36372] = i[71];
  assign o[36373] = i[71];
  assign o[36374] = i[71];
  assign o[36375] = i[71];
  assign o[36376] = i[71];
  assign o[36377] = i[71];
  assign o[36378] = i[71];
  assign o[36379] = i[71];
  assign o[36380] = i[71];
  assign o[36381] = i[71];
  assign o[36382] = i[71];
  assign o[36383] = i[71];
  assign o[36384] = i[71];
  assign o[36385] = i[71];
  assign o[36386] = i[71];
  assign o[36387] = i[71];
  assign o[36388] = i[71];
  assign o[36389] = i[71];
  assign o[36390] = i[71];
  assign o[36391] = i[71];
  assign o[36392] = i[71];
  assign o[36393] = i[71];
  assign o[36394] = i[71];
  assign o[36395] = i[71];
  assign o[36396] = i[71];
  assign o[36397] = i[71];
  assign o[36398] = i[71];
  assign o[36399] = i[71];
  assign o[36400] = i[71];
  assign o[36401] = i[71];
  assign o[36402] = i[71];
  assign o[36403] = i[71];
  assign o[36404] = i[71];
  assign o[36405] = i[71];
  assign o[36406] = i[71];
  assign o[36407] = i[71];
  assign o[36408] = i[71];
  assign o[36409] = i[71];
  assign o[36410] = i[71];
  assign o[36411] = i[71];
  assign o[36412] = i[71];
  assign o[36413] = i[71];
  assign o[36414] = i[71];
  assign o[36415] = i[71];
  assign o[36416] = i[71];
  assign o[36417] = i[71];
  assign o[36418] = i[71];
  assign o[36419] = i[71];
  assign o[36420] = i[71];
  assign o[36421] = i[71];
  assign o[36422] = i[71];
  assign o[36423] = i[71];
  assign o[36424] = i[71];
  assign o[36425] = i[71];
  assign o[36426] = i[71];
  assign o[36427] = i[71];
  assign o[36428] = i[71];
  assign o[36429] = i[71];
  assign o[36430] = i[71];
  assign o[36431] = i[71];
  assign o[36432] = i[71];
  assign o[36433] = i[71];
  assign o[36434] = i[71];
  assign o[36435] = i[71];
  assign o[36436] = i[71];
  assign o[36437] = i[71];
  assign o[36438] = i[71];
  assign o[36439] = i[71];
  assign o[36440] = i[71];
  assign o[36441] = i[71];
  assign o[36442] = i[71];
  assign o[36443] = i[71];
  assign o[36444] = i[71];
  assign o[36445] = i[71];
  assign o[36446] = i[71];
  assign o[36447] = i[71];
  assign o[36448] = i[71];
  assign o[36449] = i[71];
  assign o[36450] = i[71];
  assign o[36451] = i[71];
  assign o[36452] = i[71];
  assign o[36453] = i[71];
  assign o[36454] = i[71];
  assign o[36455] = i[71];
  assign o[36456] = i[71];
  assign o[36457] = i[71];
  assign o[36458] = i[71];
  assign o[36459] = i[71];
  assign o[36460] = i[71];
  assign o[36461] = i[71];
  assign o[36462] = i[71];
  assign o[36463] = i[71];
  assign o[36464] = i[71];
  assign o[36465] = i[71];
  assign o[36466] = i[71];
  assign o[36467] = i[71];
  assign o[36468] = i[71];
  assign o[36469] = i[71];
  assign o[36470] = i[71];
  assign o[36471] = i[71];
  assign o[36472] = i[71];
  assign o[36473] = i[71];
  assign o[36474] = i[71];
  assign o[36475] = i[71];
  assign o[36476] = i[71];
  assign o[36477] = i[71];
  assign o[36478] = i[71];
  assign o[36479] = i[71];
  assign o[36480] = i[71];
  assign o[36481] = i[71];
  assign o[36482] = i[71];
  assign o[36483] = i[71];
  assign o[36484] = i[71];
  assign o[36485] = i[71];
  assign o[36486] = i[71];
  assign o[36487] = i[71];
  assign o[36488] = i[71];
  assign o[36489] = i[71];
  assign o[36490] = i[71];
  assign o[36491] = i[71];
  assign o[36492] = i[71];
  assign o[36493] = i[71];
  assign o[36494] = i[71];
  assign o[36495] = i[71];
  assign o[36496] = i[71];
  assign o[36497] = i[71];
  assign o[36498] = i[71];
  assign o[36499] = i[71];
  assign o[36500] = i[71];
  assign o[36501] = i[71];
  assign o[36502] = i[71];
  assign o[36503] = i[71];
  assign o[36504] = i[71];
  assign o[36505] = i[71];
  assign o[36506] = i[71];
  assign o[36507] = i[71];
  assign o[36508] = i[71];
  assign o[36509] = i[71];
  assign o[36510] = i[71];
  assign o[36511] = i[71];
  assign o[36512] = i[71];
  assign o[36513] = i[71];
  assign o[36514] = i[71];
  assign o[36515] = i[71];
  assign o[36516] = i[71];
  assign o[36517] = i[71];
  assign o[36518] = i[71];
  assign o[36519] = i[71];
  assign o[36520] = i[71];
  assign o[36521] = i[71];
  assign o[36522] = i[71];
  assign o[36523] = i[71];
  assign o[36524] = i[71];
  assign o[36525] = i[71];
  assign o[36526] = i[71];
  assign o[36527] = i[71];
  assign o[36528] = i[71];
  assign o[36529] = i[71];
  assign o[36530] = i[71];
  assign o[36531] = i[71];
  assign o[36532] = i[71];
  assign o[36533] = i[71];
  assign o[36534] = i[71];
  assign o[36535] = i[71];
  assign o[36536] = i[71];
  assign o[36537] = i[71];
  assign o[36538] = i[71];
  assign o[36539] = i[71];
  assign o[36540] = i[71];
  assign o[36541] = i[71];
  assign o[36542] = i[71];
  assign o[36543] = i[71];
  assign o[36544] = i[71];
  assign o[36545] = i[71];
  assign o[36546] = i[71];
  assign o[36547] = i[71];
  assign o[36548] = i[71];
  assign o[36549] = i[71];
  assign o[36550] = i[71];
  assign o[36551] = i[71];
  assign o[36552] = i[71];
  assign o[36553] = i[71];
  assign o[36554] = i[71];
  assign o[36555] = i[71];
  assign o[36556] = i[71];
  assign o[36557] = i[71];
  assign o[36558] = i[71];
  assign o[36559] = i[71];
  assign o[36560] = i[71];
  assign o[36561] = i[71];
  assign o[36562] = i[71];
  assign o[36563] = i[71];
  assign o[36564] = i[71];
  assign o[36565] = i[71];
  assign o[36566] = i[71];
  assign o[36567] = i[71];
  assign o[36568] = i[71];
  assign o[36569] = i[71];
  assign o[36570] = i[71];
  assign o[36571] = i[71];
  assign o[36572] = i[71];
  assign o[36573] = i[71];
  assign o[36574] = i[71];
  assign o[36575] = i[71];
  assign o[36576] = i[71];
  assign o[36577] = i[71];
  assign o[36578] = i[71];
  assign o[36579] = i[71];
  assign o[36580] = i[71];
  assign o[36581] = i[71];
  assign o[36582] = i[71];
  assign o[36583] = i[71];
  assign o[36584] = i[71];
  assign o[36585] = i[71];
  assign o[36586] = i[71];
  assign o[36587] = i[71];
  assign o[36588] = i[71];
  assign o[36589] = i[71];
  assign o[36590] = i[71];
  assign o[36591] = i[71];
  assign o[36592] = i[71];
  assign o[36593] = i[71];
  assign o[36594] = i[71];
  assign o[36595] = i[71];
  assign o[36596] = i[71];
  assign o[36597] = i[71];
  assign o[36598] = i[71];
  assign o[36599] = i[71];
  assign o[36600] = i[71];
  assign o[36601] = i[71];
  assign o[36602] = i[71];
  assign o[36603] = i[71];
  assign o[36604] = i[71];
  assign o[36605] = i[71];
  assign o[36606] = i[71];
  assign o[36607] = i[71];
  assign o[36608] = i[71];
  assign o[36609] = i[71];
  assign o[36610] = i[71];
  assign o[36611] = i[71];
  assign o[36612] = i[71];
  assign o[36613] = i[71];
  assign o[36614] = i[71];
  assign o[36615] = i[71];
  assign o[36616] = i[71];
  assign o[36617] = i[71];
  assign o[36618] = i[71];
  assign o[36619] = i[71];
  assign o[36620] = i[71];
  assign o[36621] = i[71];
  assign o[36622] = i[71];
  assign o[36623] = i[71];
  assign o[36624] = i[71];
  assign o[36625] = i[71];
  assign o[36626] = i[71];
  assign o[36627] = i[71];
  assign o[36628] = i[71];
  assign o[36629] = i[71];
  assign o[36630] = i[71];
  assign o[36631] = i[71];
  assign o[36632] = i[71];
  assign o[36633] = i[71];
  assign o[36634] = i[71];
  assign o[36635] = i[71];
  assign o[36636] = i[71];
  assign o[36637] = i[71];
  assign o[36638] = i[71];
  assign o[36639] = i[71];
  assign o[36640] = i[71];
  assign o[36641] = i[71];
  assign o[36642] = i[71];
  assign o[36643] = i[71];
  assign o[36644] = i[71];
  assign o[36645] = i[71];
  assign o[36646] = i[71];
  assign o[36647] = i[71];
  assign o[36648] = i[71];
  assign o[36649] = i[71];
  assign o[36650] = i[71];
  assign o[36651] = i[71];
  assign o[36652] = i[71];
  assign o[36653] = i[71];
  assign o[36654] = i[71];
  assign o[36655] = i[71];
  assign o[36656] = i[71];
  assign o[36657] = i[71];
  assign o[36658] = i[71];
  assign o[36659] = i[71];
  assign o[36660] = i[71];
  assign o[36661] = i[71];
  assign o[36662] = i[71];
  assign o[36663] = i[71];
  assign o[36664] = i[71];
  assign o[36665] = i[71];
  assign o[36666] = i[71];
  assign o[36667] = i[71];
  assign o[36668] = i[71];
  assign o[36669] = i[71];
  assign o[36670] = i[71];
  assign o[36671] = i[71];
  assign o[36672] = i[71];
  assign o[36673] = i[71];
  assign o[36674] = i[71];
  assign o[36675] = i[71];
  assign o[36676] = i[71];
  assign o[36677] = i[71];
  assign o[36678] = i[71];
  assign o[36679] = i[71];
  assign o[36680] = i[71];
  assign o[36681] = i[71];
  assign o[36682] = i[71];
  assign o[36683] = i[71];
  assign o[36684] = i[71];
  assign o[36685] = i[71];
  assign o[36686] = i[71];
  assign o[36687] = i[71];
  assign o[36688] = i[71];
  assign o[36689] = i[71];
  assign o[36690] = i[71];
  assign o[36691] = i[71];
  assign o[36692] = i[71];
  assign o[36693] = i[71];
  assign o[36694] = i[71];
  assign o[36695] = i[71];
  assign o[36696] = i[71];
  assign o[36697] = i[71];
  assign o[36698] = i[71];
  assign o[36699] = i[71];
  assign o[36700] = i[71];
  assign o[36701] = i[71];
  assign o[36702] = i[71];
  assign o[36703] = i[71];
  assign o[36704] = i[71];
  assign o[36705] = i[71];
  assign o[36706] = i[71];
  assign o[36707] = i[71];
  assign o[36708] = i[71];
  assign o[36709] = i[71];
  assign o[36710] = i[71];
  assign o[36711] = i[71];
  assign o[36712] = i[71];
  assign o[36713] = i[71];
  assign o[36714] = i[71];
  assign o[36715] = i[71];
  assign o[36716] = i[71];
  assign o[36717] = i[71];
  assign o[36718] = i[71];
  assign o[36719] = i[71];
  assign o[36720] = i[71];
  assign o[36721] = i[71];
  assign o[36722] = i[71];
  assign o[36723] = i[71];
  assign o[36724] = i[71];
  assign o[36725] = i[71];
  assign o[36726] = i[71];
  assign o[36727] = i[71];
  assign o[36728] = i[71];
  assign o[36729] = i[71];
  assign o[36730] = i[71];
  assign o[36731] = i[71];
  assign o[36732] = i[71];
  assign o[36733] = i[71];
  assign o[36734] = i[71];
  assign o[36735] = i[71];
  assign o[36736] = i[71];
  assign o[36737] = i[71];
  assign o[36738] = i[71];
  assign o[36739] = i[71];
  assign o[36740] = i[71];
  assign o[36741] = i[71];
  assign o[36742] = i[71];
  assign o[36743] = i[71];
  assign o[36744] = i[71];
  assign o[36745] = i[71];
  assign o[36746] = i[71];
  assign o[36747] = i[71];
  assign o[36748] = i[71];
  assign o[36749] = i[71];
  assign o[36750] = i[71];
  assign o[36751] = i[71];
  assign o[36752] = i[71];
  assign o[36753] = i[71];
  assign o[36754] = i[71];
  assign o[36755] = i[71];
  assign o[36756] = i[71];
  assign o[36757] = i[71];
  assign o[36758] = i[71];
  assign o[36759] = i[71];
  assign o[36760] = i[71];
  assign o[36761] = i[71];
  assign o[36762] = i[71];
  assign o[36763] = i[71];
  assign o[36764] = i[71];
  assign o[36765] = i[71];
  assign o[36766] = i[71];
  assign o[36767] = i[71];
  assign o[36768] = i[71];
  assign o[36769] = i[71];
  assign o[36770] = i[71];
  assign o[36771] = i[71];
  assign o[36772] = i[71];
  assign o[36773] = i[71];
  assign o[36774] = i[71];
  assign o[36775] = i[71];
  assign o[36776] = i[71];
  assign o[36777] = i[71];
  assign o[36778] = i[71];
  assign o[36779] = i[71];
  assign o[36780] = i[71];
  assign o[36781] = i[71];
  assign o[36782] = i[71];
  assign o[36783] = i[71];
  assign o[36784] = i[71];
  assign o[36785] = i[71];
  assign o[36786] = i[71];
  assign o[36787] = i[71];
  assign o[36788] = i[71];
  assign o[36789] = i[71];
  assign o[36790] = i[71];
  assign o[36791] = i[71];
  assign o[36792] = i[71];
  assign o[36793] = i[71];
  assign o[36794] = i[71];
  assign o[36795] = i[71];
  assign o[36796] = i[71];
  assign o[36797] = i[71];
  assign o[36798] = i[71];
  assign o[36799] = i[71];
  assign o[36800] = i[71];
  assign o[36801] = i[71];
  assign o[36802] = i[71];
  assign o[36803] = i[71];
  assign o[36804] = i[71];
  assign o[36805] = i[71];
  assign o[36806] = i[71];
  assign o[36807] = i[71];
  assign o[36808] = i[71];
  assign o[36809] = i[71];
  assign o[36810] = i[71];
  assign o[36811] = i[71];
  assign o[36812] = i[71];
  assign o[36813] = i[71];
  assign o[36814] = i[71];
  assign o[36815] = i[71];
  assign o[36816] = i[71];
  assign o[36817] = i[71];
  assign o[36818] = i[71];
  assign o[36819] = i[71];
  assign o[36820] = i[71];
  assign o[36821] = i[71];
  assign o[36822] = i[71];
  assign o[36823] = i[71];
  assign o[36824] = i[71];
  assign o[36825] = i[71];
  assign o[36826] = i[71];
  assign o[36827] = i[71];
  assign o[36828] = i[71];
  assign o[36829] = i[71];
  assign o[36830] = i[71];
  assign o[36831] = i[71];
  assign o[36832] = i[71];
  assign o[36833] = i[71];
  assign o[36834] = i[71];
  assign o[36835] = i[71];
  assign o[36836] = i[71];
  assign o[36837] = i[71];
  assign o[36838] = i[71];
  assign o[36839] = i[71];
  assign o[36840] = i[71];
  assign o[36841] = i[71];
  assign o[36842] = i[71];
  assign o[36843] = i[71];
  assign o[36844] = i[71];
  assign o[36845] = i[71];
  assign o[36846] = i[71];
  assign o[36847] = i[71];
  assign o[36848] = i[71];
  assign o[36849] = i[71];
  assign o[36850] = i[71];
  assign o[36851] = i[71];
  assign o[36852] = i[71];
  assign o[36853] = i[71];
  assign o[36854] = i[71];
  assign o[36855] = i[71];
  assign o[36856] = i[71];
  assign o[36857] = i[71];
  assign o[36858] = i[71];
  assign o[36859] = i[71];
  assign o[36860] = i[71];
  assign o[36861] = i[71];
  assign o[36862] = i[71];
  assign o[36863] = i[71];
  assign o[35840] = i[70];
  assign o[35841] = i[70];
  assign o[35842] = i[70];
  assign o[35843] = i[70];
  assign o[35844] = i[70];
  assign o[35845] = i[70];
  assign o[35846] = i[70];
  assign o[35847] = i[70];
  assign o[35848] = i[70];
  assign o[35849] = i[70];
  assign o[35850] = i[70];
  assign o[35851] = i[70];
  assign o[35852] = i[70];
  assign o[35853] = i[70];
  assign o[35854] = i[70];
  assign o[35855] = i[70];
  assign o[35856] = i[70];
  assign o[35857] = i[70];
  assign o[35858] = i[70];
  assign o[35859] = i[70];
  assign o[35860] = i[70];
  assign o[35861] = i[70];
  assign o[35862] = i[70];
  assign o[35863] = i[70];
  assign o[35864] = i[70];
  assign o[35865] = i[70];
  assign o[35866] = i[70];
  assign o[35867] = i[70];
  assign o[35868] = i[70];
  assign o[35869] = i[70];
  assign o[35870] = i[70];
  assign o[35871] = i[70];
  assign o[35872] = i[70];
  assign o[35873] = i[70];
  assign o[35874] = i[70];
  assign o[35875] = i[70];
  assign o[35876] = i[70];
  assign o[35877] = i[70];
  assign o[35878] = i[70];
  assign o[35879] = i[70];
  assign o[35880] = i[70];
  assign o[35881] = i[70];
  assign o[35882] = i[70];
  assign o[35883] = i[70];
  assign o[35884] = i[70];
  assign o[35885] = i[70];
  assign o[35886] = i[70];
  assign o[35887] = i[70];
  assign o[35888] = i[70];
  assign o[35889] = i[70];
  assign o[35890] = i[70];
  assign o[35891] = i[70];
  assign o[35892] = i[70];
  assign o[35893] = i[70];
  assign o[35894] = i[70];
  assign o[35895] = i[70];
  assign o[35896] = i[70];
  assign o[35897] = i[70];
  assign o[35898] = i[70];
  assign o[35899] = i[70];
  assign o[35900] = i[70];
  assign o[35901] = i[70];
  assign o[35902] = i[70];
  assign o[35903] = i[70];
  assign o[35904] = i[70];
  assign o[35905] = i[70];
  assign o[35906] = i[70];
  assign o[35907] = i[70];
  assign o[35908] = i[70];
  assign o[35909] = i[70];
  assign o[35910] = i[70];
  assign o[35911] = i[70];
  assign o[35912] = i[70];
  assign o[35913] = i[70];
  assign o[35914] = i[70];
  assign o[35915] = i[70];
  assign o[35916] = i[70];
  assign o[35917] = i[70];
  assign o[35918] = i[70];
  assign o[35919] = i[70];
  assign o[35920] = i[70];
  assign o[35921] = i[70];
  assign o[35922] = i[70];
  assign o[35923] = i[70];
  assign o[35924] = i[70];
  assign o[35925] = i[70];
  assign o[35926] = i[70];
  assign o[35927] = i[70];
  assign o[35928] = i[70];
  assign o[35929] = i[70];
  assign o[35930] = i[70];
  assign o[35931] = i[70];
  assign o[35932] = i[70];
  assign o[35933] = i[70];
  assign o[35934] = i[70];
  assign o[35935] = i[70];
  assign o[35936] = i[70];
  assign o[35937] = i[70];
  assign o[35938] = i[70];
  assign o[35939] = i[70];
  assign o[35940] = i[70];
  assign o[35941] = i[70];
  assign o[35942] = i[70];
  assign o[35943] = i[70];
  assign o[35944] = i[70];
  assign o[35945] = i[70];
  assign o[35946] = i[70];
  assign o[35947] = i[70];
  assign o[35948] = i[70];
  assign o[35949] = i[70];
  assign o[35950] = i[70];
  assign o[35951] = i[70];
  assign o[35952] = i[70];
  assign o[35953] = i[70];
  assign o[35954] = i[70];
  assign o[35955] = i[70];
  assign o[35956] = i[70];
  assign o[35957] = i[70];
  assign o[35958] = i[70];
  assign o[35959] = i[70];
  assign o[35960] = i[70];
  assign o[35961] = i[70];
  assign o[35962] = i[70];
  assign o[35963] = i[70];
  assign o[35964] = i[70];
  assign o[35965] = i[70];
  assign o[35966] = i[70];
  assign o[35967] = i[70];
  assign o[35968] = i[70];
  assign o[35969] = i[70];
  assign o[35970] = i[70];
  assign o[35971] = i[70];
  assign o[35972] = i[70];
  assign o[35973] = i[70];
  assign o[35974] = i[70];
  assign o[35975] = i[70];
  assign o[35976] = i[70];
  assign o[35977] = i[70];
  assign o[35978] = i[70];
  assign o[35979] = i[70];
  assign o[35980] = i[70];
  assign o[35981] = i[70];
  assign o[35982] = i[70];
  assign o[35983] = i[70];
  assign o[35984] = i[70];
  assign o[35985] = i[70];
  assign o[35986] = i[70];
  assign o[35987] = i[70];
  assign o[35988] = i[70];
  assign o[35989] = i[70];
  assign o[35990] = i[70];
  assign o[35991] = i[70];
  assign o[35992] = i[70];
  assign o[35993] = i[70];
  assign o[35994] = i[70];
  assign o[35995] = i[70];
  assign o[35996] = i[70];
  assign o[35997] = i[70];
  assign o[35998] = i[70];
  assign o[35999] = i[70];
  assign o[36000] = i[70];
  assign o[36001] = i[70];
  assign o[36002] = i[70];
  assign o[36003] = i[70];
  assign o[36004] = i[70];
  assign o[36005] = i[70];
  assign o[36006] = i[70];
  assign o[36007] = i[70];
  assign o[36008] = i[70];
  assign o[36009] = i[70];
  assign o[36010] = i[70];
  assign o[36011] = i[70];
  assign o[36012] = i[70];
  assign o[36013] = i[70];
  assign o[36014] = i[70];
  assign o[36015] = i[70];
  assign o[36016] = i[70];
  assign o[36017] = i[70];
  assign o[36018] = i[70];
  assign o[36019] = i[70];
  assign o[36020] = i[70];
  assign o[36021] = i[70];
  assign o[36022] = i[70];
  assign o[36023] = i[70];
  assign o[36024] = i[70];
  assign o[36025] = i[70];
  assign o[36026] = i[70];
  assign o[36027] = i[70];
  assign o[36028] = i[70];
  assign o[36029] = i[70];
  assign o[36030] = i[70];
  assign o[36031] = i[70];
  assign o[36032] = i[70];
  assign o[36033] = i[70];
  assign o[36034] = i[70];
  assign o[36035] = i[70];
  assign o[36036] = i[70];
  assign o[36037] = i[70];
  assign o[36038] = i[70];
  assign o[36039] = i[70];
  assign o[36040] = i[70];
  assign o[36041] = i[70];
  assign o[36042] = i[70];
  assign o[36043] = i[70];
  assign o[36044] = i[70];
  assign o[36045] = i[70];
  assign o[36046] = i[70];
  assign o[36047] = i[70];
  assign o[36048] = i[70];
  assign o[36049] = i[70];
  assign o[36050] = i[70];
  assign o[36051] = i[70];
  assign o[36052] = i[70];
  assign o[36053] = i[70];
  assign o[36054] = i[70];
  assign o[36055] = i[70];
  assign o[36056] = i[70];
  assign o[36057] = i[70];
  assign o[36058] = i[70];
  assign o[36059] = i[70];
  assign o[36060] = i[70];
  assign o[36061] = i[70];
  assign o[36062] = i[70];
  assign o[36063] = i[70];
  assign o[36064] = i[70];
  assign o[36065] = i[70];
  assign o[36066] = i[70];
  assign o[36067] = i[70];
  assign o[36068] = i[70];
  assign o[36069] = i[70];
  assign o[36070] = i[70];
  assign o[36071] = i[70];
  assign o[36072] = i[70];
  assign o[36073] = i[70];
  assign o[36074] = i[70];
  assign o[36075] = i[70];
  assign o[36076] = i[70];
  assign o[36077] = i[70];
  assign o[36078] = i[70];
  assign o[36079] = i[70];
  assign o[36080] = i[70];
  assign o[36081] = i[70];
  assign o[36082] = i[70];
  assign o[36083] = i[70];
  assign o[36084] = i[70];
  assign o[36085] = i[70];
  assign o[36086] = i[70];
  assign o[36087] = i[70];
  assign o[36088] = i[70];
  assign o[36089] = i[70];
  assign o[36090] = i[70];
  assign o[36091] = i[70];
  assign o[36092] = i[70];
  assign o[36093] = i[70];
  assign o[36094] = i[70];
  assign o[36095] = i[70];
  assign o[36096] = i[70];
  assign o[36097] = i[70];
  assign o[36098] = i[70];
  assign o[36099] = i[70];
  assign o[36100] = i[70];
  assign o[36101] = i[70];
  assign o[36102] = i[70];
  assign o[36103] = i[70];
  assign o[36104] = i[70];
  assign o[36105] = i[70];
  assign o[36106] = i[70];
  assign o[36107] = i[70];
  assign o[36108] = i[70];
  assign o[36109] = i[70];
  assign o[36110] = i[70];
  assign o[36111] = i[70];
  assign o[36112] = i[70];
  assign o[36113] = i[70];
  assign o[36114] = i[70];
  assign o[36115] = i[70];
  assign o[36116] = i[70];
  assign o[36117] = i[70];
  assign o[36118] = i[70];
  assign o[36119] = i[70];
  assign o[36120] = i[70];
  assign o[36121] = i[70];
  assign o[36122] = i[70];
  assign o[36123] = i[70];
  assign o[36124] = i[70];
  assign o[36125] = i[70];
  assign o[36126] = i[70];
  assign o[36127] = i[70];
  assign o[36128] = i[70];
  assign o[36129] = i[70];
  assign o[36130] = i[70];
  assign o[36131] = i[70];
  assign o[36132] = i[70];
  assign o[36133] = i[70];
  assign o[36134] = i[70];
  assign o[36135] = i[70];
  assign o[36136] = i[70];
  assign o[36137] = i[70];
  assign o[36138] = i[70];
  assign o[36139] = i[70];
  assign o[36140] = i[70];
  assign o[36141] = i[70];
  assign o[36142] = i[70];
  assign o[36143] = i[70];
  assign o[36144] = i[70];
  assign o[36145] = i[70];
  assign o[36146] = i[70];
  assign o[36147] = i[70];
  assign o[36148] = i[70];
  assign o[36149] = i[70];
  assign o[36150] = i[70];
  assign o[36151] = i[70];
  assign o[36152] = i[70];
  assign o[36153] = i[70];
  assign o[36154] = i[70];
  assign o[36155] = i[70];
  assign o[36156] = i[70];
  assign o[36157] = i[70];
  assign o[36158] = i[70];
  assign o[36159] = i[70];
  assign o[36160] = i[70];
  assign o[36161] = i[70];
  assign o[36162] = i[70];
  assign o[36163] = i[70];
  assign o[36164] = i[70];
  assign o[36165] = i[70];
  assign o[36166] = i[70];
  assign o[36167] = i[70];
  assign o[36168] = i[70];
  assign o[36169] = i[70];
  assign o[36170] = i[70];
  assign o[36171] = i[70];
  assign o[36172] = i[70];
  assign o[36173] = i[70];
  assign o[36174] = i[70];
  assign o[36175] = i[70];
  assign o[36176] = i[70];
  assign o[36177] = i[70];
  assign o[36178] = i[70];
  assign o[36179] = i[70];
  assign o[36180] = i[70];
  assign o[36181] = i[70];
  assign o[36182] = i[70];
  assign o[36183] = i[70];
  assign o[36184] = i[70];
  assign o[36185] = i[70];
  assign o[36186] = i[70];
  assign o[36187] = i[70];
  assign o[36188] = i[70];
  assign o[36189] = i[70];
  assign o[36190] = i[70];
  assign o[36191] = i[70];
  assign o[36192] = i[70];
  assign o[36193] = i[70];
  assign o[36194] = i[70];
  assign o[36195] = i[70];
  assign o[36196] = i[70];
  assign o[36197] = i[70];
  assign o[36198] = i[70];
  assign o[36199] = i[70];
  assign o[36200] = i[70];
  assign o[36201] = i[70];
  assign o[36202] = i[70];
  assign o[36203] = i[70];
  assign o[36204] = i[70];
  assign o[36205] = i[70];
  assign o[36206] = i[70];
  assign o[36207] = i[70];
  assign o[36208] = i[70];
  assign o[36209] = i[70];
  assign o[36210] = i[70];
  assign o[36211] = i[70];
  assign o[36212] = i[70];
  assign o[36213] = i[70];
  assign o[36214] = i[70];
  assign o[36215] = i[70];
  assign o[36216] = i[70];
  assign o[36217] = i[70];
  assign o[36218] = i[70];
  assign o[36219] = i[70];
  assign o[36220] = i[70];
  assign o[36221] = i[70];
  assign o[36222] = i[70];
  assign o[36223] = i[70];
  assign o[36224] = i[70];
  assign o[36225] = i[70];
  assign o[36226] = i[70];
  assign o[36227] = i[70];
  assign o[36228] = i[70];
  assign o[36229] = i[70];
  assign o[36230] = i[70];
  assign o[36231] = i[70];
  assign o[36232] = i[70];
  assign o[36233] = i[70];
  assign o[36234] = i[70];
  assign o[36235] = i[70];
  assign o[36236] = i[70];
  assign o[36237] = i[70];
  assign o[36238] = i[70];
  assign o[36239] = i[70];
  assign o[36240] = i[70];
  assign o[36241] = i[70];
  assign o[36242] = i[70];
  assign o[36243] = i[70];
  assign o[36244] = i[70];
  assign o[36245] = i[70];
  assign o[36246] = i[70];
  assign o[36247] = i[70];
  assign o[36248] = i[70];
  assign o[36249] = i[70];
  assign o[36250] = i[70];
  assign o[36251] = i[70];
  assign o[36252] = i[70];
  assign o[36253] = i[70];
  assign o[36254] = i[70];
  assign o[36255] = i[70];
  assign o[36256] = i[70];
  assign o[36257] = i[70];
  assign o[36258] = i[70];
  assign o[36259] = i[70];
  assign o[36260] = i[70];
  assign o[36261] = i[70];
  assign o[36262] = i[70];
  assign o[36263] = i[70];
  assign o[36264] = i[70];
  assign o[36265] = i[70];
  assign o[36266] = i[70];
  assign o[36267] = i[70];
  assign o[36268] = i[70];
  assign o[36269] = i[70];
  assign o[36270] = i[70];
  assign o[36271] = i[70];
  assign o[36272] = i[70];
  assign o[36273] = i[70];
  assign o[36274] = i[70];
  assign o[36275] = i[70];
  assign o[36276] = i[70];
  assign o[36277] = i[70];
  assign o[36278] = i[70];
  assign o[36279] = i[70];
  assign o[36280] = i[70];
  assign o[36281] = i[70];
  assign o[36282] = i[70];
  assign o[36283] = i[70];
  assign o[36284] = i[70];
  assign o[36285] = i[70];
  assign o[36286] = i[70];
  assign o[36287] = i[70];
  assign o[36288] = i[70];
  assign o[36289] = i[70];
  assign o[36290] = i[70];
  assign o[36291] = i[70];
  assign o[36292] = i[70];
  assign o[36293] = i[70];
  assign o[36294] = i[70];
  assign o[36295] = i[70];
  assign o[36296] = i[70];
  assign o[36297] = i[70];
  assign o[36298] = i[70];
  assign o[36299] = i[70];
  assign o[36300] = i[70];
  assign o[36301] = i[70];
  assign o[36302] = i[70];
  assign o[36303] = i[70];
  assign o[36304] = i[70];
  assign o[36305] = i[70];
  assign o[36306] = i[70];
  assign o[36307] = i[70];
  assign o[36308] = i[70];
  assign o[36309] = i[70];
  assign o[36310] = i[70];
  assign o[36311] = i[70];
  assign o[36312] = i[70];
  assign o[36313] = i[70];
  assign o[36314] = i[70];
  assign o[36315] = i[70];
  assign o[36316] = i[70];
  assign o[36317] = i[70];
  assign o[36318] = i[70];
  assign o[36319] = i[70];
  assign o[36320] = i[70];
  assign o[36321] = i[70];
  assign o[36322] = i[70];
  assign o[36323] = i[70];
  assign o[36324] = i[70];
  assign o[36325] = i[70];
  assign o[36326] = i[70];
  assign o[36327] = i[70];
  assign o[36328] = i[70];
  assign o[36329] = i[70];
  assign o[36330] = i[70];
  assign o[36331] = i[70];
  assign o[36332] = i[70];
  assign o[36333] = i[70];
  assign o[36334] = i[70];
  assign o[36335] = i[70];
  assign o[36336] = i[70];
  assign o[36337] = i[70];
  assign o[36338] = i[70];
  assign o[36339] = i[70];
  assign o[36340] = i[70];
  assign o[36341] = i[70];
  assign o[36342] = i[70];
  assign o[36343] = i[70];
  assign o[36344] = i[70];
  assign o[36345] = i[70];
  assign o[36346] = i[70];
  assign o[36347] = i[70];
  assign o[36348] = i[70];
  assign o[36349] = i[70];
  assign o[36350] = i[70];
  assign o[36351] = i[70];
  assign o[35328] = i[69];
  assign o[35329] = i[69];
  assign o[35330] = i[69];
  assign o[35331] = i[69];
  assign o[35332] = i[69];
  assign o[35333] = i[69];
  assign o[35334] = i[69];
  assign o[35335] = i[69];
  assign o[35336] = i[69];
  assign o[35337] = i[69];
  assign o[35338] = i[69];
  assign o[35339] = i[69];
  assign o[35340] = i[69];
  assign o[35341] = i[69];
  assign o[35342] = i[69];
  assign o[35343] = i[69];
  assign o[35344] = i[69];
  assign o[35345] = i[69];
  assign o[35346] = i[69];
  assign o[35347] = i[69];
  assign o[35348] = i[69];
  assign o[35349] = i[69];
  assign o[35350] = i[69];
  assign o[35351] = i[69];
  assign o[35352] = i[69];
  assign o[35353] = i[69];
  assign o[35354] = i[69];
  assign o[35355] = i[69];
  assign o[35356] = i[69];
  assign o[35357] = i[69];
  assign o[35358] = i[69];
  assign o[35359] = i[69];
  assign o[35360] = i[69];
  assign o[35361] = i[69];
  assign o[35362] = i[69];
  assign o[35363] = i[69];
  assign o[35364] = i[69];
  assign o[35365] = i[69];
  assign o[35366] = i[69];
  assign o[35367] = i[69];
  assign o[35368] = i[69];
  assign o[35369] = i[69];
  assign o[35370] = i[69];
  assign o[35371] = i[69];
  assign o[35372] = i[69];
  assign o[35373] = i[69];
  assign o[35374] = i[69];
  assign o[35375] = i[69];
  assign o[35376] = i[69];
  assign o[35377] = i[69];
  assign o[35378] = i[69];
  assign o[35379] = i[69];
  assign o[35380] = i[69];
  assign o[35381] = i[69];
  assign o[35382] = i[69];
  assign o[35383] = i[69];
  assign o[35384] = i[69];
  assign o[35385] = i[69];
  assign o[35386] = i[69];
  assign o[35387] = i[69];
  assign o[35388] = i[69];
  assign o[35389] = i[69];
  assign o[35390] = i[69];
  assign o[35391] = i[69];
  assign o[35392] = i[69];
  assign o[35393] = i[69];
  assign o[35394] = i[69];
  assign o[35395] = i[69];
  assign o[35396] = i[69];
  assign o[35397] = i[69];
  assign o[35398] = i[69];
  assign o[35399] = i[69];
  assign o[35400] = i[69];
  assign o[35401] = i[69];
  assign o[35402] = i[69];
  assign o[35403] = i[69];
  assign o[35404] = i[69];
  assign o[35405] = i[69];
  assign o[35406] = i[69];
  assign o[35407] = i[69];
  assign o[35408] = i[69];
  assign o[35409] = i[69];
  assign o[35410] = i[69];
  assign o[35411] = i[69];
  assign o[35412] = i[69];
  assign o[35413] = i[69];
  assign o[35414] = i[69];
  assign o[35415] = i[69];
  assign o[35416] = i[69];
  assign o[35417] = i[69];
  assign o[35418] = i[69];
  assign o[35419] = i[69];
  assign o[35420] = i[69];
  assign o[35421] = i[69];
  assign o[35422] = i[69];
  assign o[35423] = i[69];
  assign o[35424] = i[69];
  assign o[35425] = i[69];
  assign o[35426] = i[69];
  assign o[35427] = i[69];
  assign o[35428] = i[69];
  assign o[35429] = i[69];
  assign o[35430] = i[69];
  assign o[35431] = i[69];
  assign o[35432] = i[69];
  assign o[35433] = i[69];
  assign o[35434] = i[69];
  assign o[35435] = i[69];
  assign o[35436] = i[69];
  assign o[35437] = i[69];
  assign o[35438] = i[69];
  assign o[35439] = i[69];
  assign o[35440] = i[69];
  assign o[35441] = i[69];
  assign o[35442] = i[69];
  assign o[35443] = i[69];
  assign o[35444] = i[69];
  assign o[35445] = i[69];
  assign o[35446] = i[69];
  assign o[35447] = i[69];
  assign o[35448] = i[69];
  assign o[35449] = i[69];
  assign o[35450] = i[69];
  assign o[35451] = i[69];
  assign o[35452] = i[69];
  assign o[35453] = i[69];
  assign o[35454] = i[69];
  assign o[35455] = i[69];
  assign o[35456] = i[69];
  assign o[35457] = i[69];
  assign o[35458] = i[69];
  assign o[35459] = i[69];
  assign o[35460] = i[69];
  assign o[35461] = i[69];
  assign o[35462] = i[69];
  assign o[35463] = i[69];
  assign o[35464] = i[69];
  assign o[35465] = i[69];
  assign o[35466] = i[69];
  assign o[35467] = i[69];
  assign o[35468] = i[69];
  assign o[35469] = i[69];
  assign o[35470] = i[69];
  assign o[35471] = i[69];
  assign o[35472] = i[69];
  assign o[35473] = i[69];
  assign o[35474] = i[69];
  assign o[35475] = i[69];
  assign o[35476] = i[69];
  assign o[35477] = i[69];
  assign o[35478] = i[69];
  assign o[35479] = i[69];
  assign o[35480] = i[69];
  assign o[35481] = i[69];
  assign o[35482] = i[69];
  assign o[35483] = i[69];
  assign o[35484] = i[69];
  assign o[35485] = i[69];
  assign o[35486] = i[69];
  assign o[35487] = i[69];
  assign o[35488] = i[69];
  assign o[35489] = i[69];
  assign o[35490] = i[69];
  assign o[35491] = i[69];
  assign o[35492] = i[69];
  assign o[35493] = i[69];
  assign o[35494] = i[69];
  assign o[35495] = i[69];
  assign o[35496] = i[69];
  assign o[35497] = i[69];
  assign o[35498] = i[69];
  assign o[35499] = i[69];
  assign o[35500] = i[69];
  assign o[35501] = i[69];
  assign o[35502] = i[69];
  assign o[35503] = i[69];
  assign o[35504] = i[69];
  assign o[35505] = i[69];
  assign o[35506] = i[69];
  assign o[35507] = i[69];
  assign o[35508] = i[69];
  assign o[35509] = i[69];
  assign o[35510] = i[69];
  assign o[35511] = i[69];
  assign o[35512] = i[69];
  assign o[35513] = i[69];
  assign o[35514] = i[69];
  assign o[35515] = i[69];
  assign o[35516] = i[69];
  assign o[35517] = i[69];
  assign o[35518] = i[69];
  assign o[35519] = i[69];
  assign o[35520] = i[69];
  assign o[35521] = i[69];
  assign o[35522] = i[69];
  assign o[35523] = i[69];
  assign o[35524] = i[69];
  assign o[35525] = i[69];
  assign o[35526] = i[69];
  assign o[35527] = i[69];
  assign o[35528] = i[69];
  assign o[35529] = i[69];
  assign o[35530] = i[69];
  assign o[35531] = i[69];
  assign o[35532] = i[69];
  assign o[35533] = i[69];
  assign o[35534] = i[69];
  assign o[35535] = i[69];
  assign o[35536] = i[69];
  assign o[35537] = i[69];
  assign o[35538] = i[69];
  assign o[35539] = i[69];
  assign o[35540] = i[69];
  assign o[35541] = i[69];
  assign o[35542] = i[69];
  assign o[35543] = i[69];
  assign o[35544] = i[69];
  assign o[35545] = i[69];
  assign o[35546] = i[69];
  assign o[35547] = i[69];
  assign o[35548] = i[69];
  assign o[35549] = i[69];
  assign o[35550] = i[69];
  assign o[35551] = i[69];
  assign o[35552] = i[69];
  assign o[35553] = i[69];
  assign o[35554] = i[69];
  assign o[35555] = i[69];
  assign o[35556] = i[69];
  assign o[35557] = i[69];
  assign o[35558] = i[69];
  assign o[35559] = i[69];
  assign o[35560] = i[69];
  assign o[35561] = i[69];
  assign o[35562] = i[69];
  assign o[35563] = i[69];
  assign o[35564] = i[69];
  assign o[35565] = i[69];
  assign o[35566] = i[69];
  assign o[35567] = i[69];
  assign o[35568] = i[69];
  assign o[35569] = i[69];
  assign o[35570] = i[69];
  assign o[35571] = i[69];
  assign o[35572] = i[69];
  assign o[35573] = i[69];
  assign o[35574] = i[69];
  assign o[35575] = i[69];
  assign o[35576] = i[69];
  assign o[35577] = i[69];
  assign o[35578] = i[69];
  assign o[35579] = i[69];
  assign o[35580] = i[69];
  assign o[35581] = i[69];
  assign o[35582] = i[69];
  assign o[35583] = i[69];
  assign o[35584] = i[69];
  assign o[35585] = i[69];
  assign o[35586] = i[69];
  assign o[35587] = i[69];
  assign o[35588] = i[69];
  assign o[35589] = i[69];
  assign o[35590] = i[69];
  assign o[35591] = i[69];
  assign o[35592] = i[69];
  assign o[35593] = i[69];
  assign o[35594] = i[69];
  assign o[35595] = i[69];
  assign o[35596] = i[69];
  assign o[35597] = i[69];
  assign o[35598] = i[69];
  assign o[35599] = i[69];
  assign o[35600] = i[69];
  assign o[35601] = i[69];
  assign o[35602] = i[69];
  assign o[35603] = i[69];
  assign o[35604] = i[69];
  assign o[35605] = i[69];
  assign o[35606] = i[69];
  assign o[35607] = i[69];
  assign o[35608] = i[69];
  assign o[35609] = i[69];
  assign o[35610] = i[69];
  assign o[35611] = i[69];
  assign o[35612] = i[69];
  assign o[35613] = i[69];
  assign o[35614] = i[69];
  assign o[35615] = i[69];
  assign o[35616] = i[69];
  assign o[35617] = i[69];
  assign o[35618] = i[69];
  assign o[35619] = i[69];
  assign o[35620] = i[69];
  assign o[35621] = i[69];
  assign o[35622] = i[69];
  assign o[35623] = i[69];
  assign o[35624] = i[69];
  assign o[35625] = i[69];
  assign o[35626] = i[69];
  assign o[35627] = i[69];
  assign o[35628] = i[69];
  assign o[35629] = i[69];
  assign o[35630] = i[69];
  assign o[35631] = i[69];
  assign o[35632] = i[69];
  assign o[35633] = i[69];
  assign o[35634] = i[69];
  assign o[35635] = i[69];
  assign o[35636] = i[69];
  assign o[35637] = i[69];
  assign o[35638] = i[69];
  assign o[35639] = i[69];
  assign o[35640] = i[69];
  assign o[35641] = i[69];
  assign o[35642] = i[69];
  assign o[35643] = i[69];
  assign o[35644] = i[69];
  assign o[35645] = i[69];
  assign o[35646] = i[69];
  assign o[35647] = i[69];
  assign o[35648] = i[69];
  assign o[35649] = i[69];
  assign o[35650] = i[69];
  assign o[35651] = i[69];
  assign o[35652] = i[69];
  assign o[35653] = i[69];
  assign o[35654] = i[69];
  assign o[35655] = i[69];
  assign o[35656] = i[69];
  assign o[35657] = i[69];
  assign o[35658] = i[69];
  assign o[35659] = i[69];
  assign o[35660] = i[69];
  assign o[35661] = i[69];
  assign o[35662] = i[69];
  assign o[35663] = i[69];
  assign o[35664] = i[69];
  assign o[35665] = i[69];
  assign o[35666] = i[69];
  assign o[35667] = i[69];
  assign o[35668] = i[69];
  assign o[35669] = i[69];
  assign o[35670] = i[69];
  assign o[35671] = i[69];
  assign o[35672] = i[69];
  assign o[35673] = i[69];
  assign o[35674] = i[69];
  assign o[35675] = i[69];
  assign o[35676] = i[69];
  assign o[35677] = i[69];
  assign o[35678] = i[69];
  assign o[35679] = i[69];
  assign o[35680] = i[69];
  assign o[35681] = i[69];
  assign o[35682] = i[69];
  assign o[35683] = i[69];
  assign o[35684] = i[69];
  assign o[35685] = i[69];
  assign o[35686] = i[69];
  assign o[35687] = i[69];
  assign o[35688] = i[69];
  assign o[35689] = i[69];
  assign o[35690] = i[69];
  assign o[35691] = i[69];
  assign o[35692] = i[69];
  assign o[35693] = i[69];
  assign o[35694] = i[69];
  assign o[35695] = i[69];
  assign o[35696] = i[69];
  assign o[35697] = i[69];
  assign o[35698] = i[69];
  assign o[35699] = i[69];
  assign o[35700] = i[69];
  assign o[35701] = i[69];
  assign o[35702] = i[69];
  assign o[35703] = i[69];
  assign o[35704] = i[69];
  assign o[35705] = i[69];
  assign o[35706] = i[69];
  assign o[35707] = i[69];
  assign o[35708] = i[69];
  assign o[35709] = i[69];
  assign o[35710] = i[69];
  assign o[35711] = i[69];
  assign o[35712] = i[69];
  assign o[35713] = i[69];
  assign o[35714] = i[69];
  assign o[35715] = i[69];
  assign o[35716] = i[69];
  assign o[35717] = i[69];
  assign o[35718] = i[69];
  assign o[35719] = i[69];
  assign o[35720] = i[69];
  assign o[35721] = i[69];
  assign o[35722] = i[69];
  assign o[35723] = i[69];
  assign o[35724] = i[69];
  assign o[35725] = i[69];
  assign o[35726] = i[69];
  assign o[35727] = i[69];
  assign o[35728] = i[69];
  assign o[35729] = i[69];
  assign o[35730] = i[69];
  assign o[35731] = i[69];
  assign o[35732] = i[69];
  assign o[35733] = i[69];
  assign o[35734] = i[69];
  assign o[35735] = i[69];
  assign o[35736] = i[69];
  assign o[35737] = i[69];
  assign o[35738] = i[69];
  assign o[35739] = i[69];
  assign o[35740] = i[69];
  assign o[35741] = i[69];
  assign o[35742] = i[69];
  assign o[35743] = i[69];
  assign o[35744] = i[69];
  assign o[35745] = i[69];
  assign o[35746] = i[69];
  assign o[35747] = i[69];
  assign o[35748] = i[69];
  assign o[35749] = i[69];
  assign o[35750] = i[69];
  assign o[35751] = i[69];
  assign o[35752] = i[69];
  assign o[35753] = i[69];
  assign o[35754] = i[69];
  assign o[35755] = i[69];
  assign o[35756] = i[69];
  assign o[35757] = i[69];
  assign o[35758] = i[69];
  assign o[35759] = i[69];
  assign o[35760] = i[69];
  assign o[35761] = i[69];
  assign o[35762] = i[69];
  assign o[35763] = i[69];
  assign o[35764] = i[69];
  assign o[35765] = i[69];
  assign o[35766] = i[69];
  assign o[35767] = i[69];
  assign o[35768] = i[69];
  assign o[35769] = i[69];
  assign o[35770] = i[69];
  assign o[35771] = i[69];
  assign o[35772] = i[69];
  assign o[35773] = i[69];
  assign o[35774] = i[69];
  assign o[35775] = i[69];
  assign o[35776] = i[69];
  assign o[35777] = i[69];
  assign o[35778] = i[69];
  assign o[35779] = i[69];
  assign o[35780] = i[69];
  assign o[35781] = i[69];
  assign o[35782] = i[69];
  assign o[35783] = i[69];
  assign o[35784] = i[69];
  assign o[35785] = i[69];
  assign o[35786] = i[69];
  assign o[35787] = i[69];
  assign o[35788] = i[69];
  assign o[35789] = i[69];
  assign o[35790] = i[69];
  assign o[35791] = i[69];
  assign o[35792] = i[69];
  assign o[35793] = i[69];
  assign o[35794] = i[69];
  assign o[35795] = i[69];
  assign o[35796] = i[69];
  assign o[35797] = i[69];
  assign o[35798] = i[69];
  assign o[35799] = i[69];
  assign o[35800] = i[69];
  assign o[35801] = i[69];
  assign o[35802] = i[69];
  assign o[35803] = i[69];
  assign o[35804] = i[69];
  assign o[35805] = i[69];
  assign o[35806] = i[69];
  assign o[35807] = i[69];
  assign o[35808] = i[69];
  assign o[35809] = i[69];
  assign o[35810] = i[69];
  assign o[35811] = i[69];
  assign o[35812] = i[69];
  assign o[35813] = i[69];
  assign o[35814] = i[69];
  assign o[35815] = i[69];
  assign o[35816] = i[69];
  assign o[35817] = i[69];
  assign o[35818] = i[69];
  assign o[35819] = i[69];
  assign o[35820] = i[69];
  assign o[35821] = i[69];
  assign o[35822] = i[69];
  assign o[35823] = i[69];
  assign o[35824] = i[69];
  assign o[35825] = i[69];
  assign o[35826] = i[69];
  assign o[35827] = i[69];
  assign o[35828] = i[69];
  assign o[35829] = i[69];
  assign o[35830] = i[69];
  assign o[35831] = i[69];
  assign o[35832] = i[69];
  assign o[35833] = i[69];
  assign o[35834] = i[69];
  assign o[35835] = i[69];
  assign o[35836] = i[69];
  assign o[35837] = i[69];
  assign o[35838] = i[69];
  assign o[35839] = i[69];
  assign o[34816] = i[68];
  assign o[34817] = i[68];
  assign o[34818] = i[68];
  assign o[34819] = i[68];
  assign o[34820] = i[68];
  assign o[34821] = i[68];
  assign o[34822] = i[68];
  assign o[34823] = i[68];
  assign o[34824] = i[68];
  assign o[34825] = i[68];
  assign o[34826] = i[68];
  assign o[34827] = i[68];
  assign o[34828] = i[68];
  assign o[34829] = i[68];
  assign o[34830] = i[68];
  assign o[34831] = i[68];
  assign o[34832] = i[68];
  assign o[34833] = i[68];
  assign o[34834] = i[68];
  assign o[34835] = i[68];
  assign o[34836] = i[68];
  assign o[34837] = i[68];
  assign o[34838] = i[68];
  assign o[34839] = i[68];
  assign o[34840] = i[68];
  assign o[34841] = i[68];
  assign o[34842] = i[68];
  assign o[34843] = i[68];
  assign o[34844] = i[68];
  assign o[34845] = i[68];
  assign o[34846] = i[68];
  assign o[34847] = i[68];
  assign o[34848] = i[68];
  assign o[34849] = i[68];
  assign o[34850] = i[68];
  assign o[34851] = i[68];
  assign o[34852] = i[68];
  assign o[34853] = i[68];
  assign o[34854] = i[68];
  assign o[34855] = i[68];
  assign o[34856] = i[68];
  assign o[34857] = i[68];
  assign o[34858] = i[68];
  assign o[34859] = i[68];
  assign o[34860] = i[68];
  assign o[34861] = i[68];
  assign o[34862] = i[68];
  assign o[34863] = i[68];
  assign o[34864] = i[68];
  assign o[34865] = i[68];
  assign o[34866] = i[68];
  assign o[34867] = i[68];
  assign o[34868] = i[68];
  assign o[34869] = i[68];
  assign o[34870] = i[68];
  assign o[34871] = i[68];
  assign o[34872] = i[68];
  assign o[34873] = i[68];
  assign o[34874] = i[68];
  assign o[34875] = i[68];
  assign o[34876] = i[68];
  assign o[34877] = i[68];
  assign o[34878] = i[68];
  assign o[34879] = i[68];
  assign o[34880] = i[68];
  assign o[34881] = i[68];
  assign o[34882] = i[68];
  assign o[34883] = i[68];
  assign o[34884] = i[68];
  assign o[34885] = i[68];
  assign o[34886] = i[68];
  assign o[34887] = i[68];
  assign o[34888] = i[68];
  assign o[34889] = i[68];
  assign o[34890] = i[68];
  assign o[34891] = i[68];
  assign o[34892] = i[68];
  assign o[34893] = i[68];
  assign o[34894] = i[68];
  assign o[34895] = i[68];
  assign o[34896] = i[68];
  assign o[34897] = i[68];
  assign o[34898] = i[68];
  assign o[34899] = i[68];
  assign o[34900] = i[68];
  assign o[34901] = i[68];
  assign o[34902] = i[68];
  assign o[34903] = i[68];
  assign o[34904] = i[68];
  assign o[34905] = i[68];
  assign o[34906] = i[68];
  assign o[34907] = i[68];
  assign o[34908] = i[68];
  assign o[34909] = i[68];
  assign o[34910] = i[68];
  assign o[34911] = i[68];
  assign o[34912] = i[68];
  assign o[34913] = i[68];
  assign o[34914] = i[68];
  assign o[34915] = i[68];
  assign o[34916] = i[68];
  assign o[34917] = i[68];
  assign o[34918] = i[68];
  assign o[34919] = i[68];
  assign o[34920] = i[68];
  assign o[34921] = i[68];
  assign o[34922] = i[68];
  assign o[34923] = i[68];
  assign o[34924] = i[68];
  assign o[34925] = i[68];
  assign o[34926] = i[68];
  assign o[34927] = i[68];
  assign o[34928] = i[68];
  assign o[34929] = i[68];
  assign o[34930] = i[68];
  assign o[34931] = i[68];
  assign o[34932] = i[68];
  assign o[34933] = i[68];
  assign o[34934] = i[68];
  assign o[34935] = i[68];
  assign o[34936] = i[68];
  assign o[34937] = i[68];
  assign o[34938] = i[68];
  assign o[34939] = i[68];
  assign o[34940] = i[68];
  assign o[34941] = i[68];
  assign o[34942] = i[68];
  assign o[34943] = i[68];
  assign o[34944] = i[68];
  assign o[34945] = i[68];
  assign o[34946] = i[68];
  assign o[34947] = i[68];
  assign o[34948] = i[68];
  assign o[34949] = i[68];
  assign o[34950] = i[68];
  assign o[34951] = i[68];
  assign o[34952] = i[68];
  assign o[34953] = i[68];
  assign o[34954] = i[68];
  assign o[34955] = i[68];
  assign o[34956] = i[68];
  assign o[34957] = i[68];
  assign o[34958] = i[68];
  assign o[34959] = i[68];
  assign o[34960] = i[68];
  assign o[34961] = i[68];
  assign o[34962] = i[68];
  assign o[34963] = i[68];
  assign o[34964] = i[68];
  assign o[34965] = i[68];
  assign o[34966] = i[68];
  assign o[34967] = i[68];
  assign o[34968] = i[68];
  assign o[34969] = i[68];
  assign o[34970] = i[68];
  assign o[34971] = i[68];
  assign o[34972] = i[68];
  assign o[34973] = i[68];
  assign o[34974] = i[68];
  assign o[34975] = i[68];
  assign o[34976] = i[68];
  assign o[34977] = i[68];
  assign o[34978] = i[68];
  assign o[34979] = i[68];
  assign o[34980] = i[68];
  assign o[34981] = i[68];
  assign o[34982] = i[68];
  assign o[34983] = i[68];
  assign o[34984] = i[68];
  assign o[34985] = i[68];
  assign o[34986] = i[68];
  assign o[34987] = i[68];
  assign o[34988] = i[68];
  assign o[34989] = i[68];
  assign o[34990] = i[68];
  assign o[34991] = i[68];
  assign o[34992] = i[68];
  assign o[34993] = i[68];
  assign o[34994] = i[68];
  assign o[34995] = i[68];
  assign o[34996] = i[68];
  assign o[34997] = i[68];
  assign o[34998] = i[68];
  assign o[34999] = i[68];
  assign o[35000] = i[68];
  assign o[35001] = i[68];
  assign o[35002] = i[68];
  assign o[35003] = i[68];
  assign o[35004] = i[68];
  assign o[35005] = i[68];
  assign o[35006] = i[68];
  assign o[35007] = i[68];
  assign o[35008] = i[68];
  assign o[35009] = i[68];
  assign o[35010] = i[68];
  assign o[35011] = i[68];
  assign o[35012] = i[68];
  assign o[35013] = i[68];
  assign o[35014] = i[68];
  assign o[35015] = i[68];
  assign o[35016] = i[68];
  assign o[35017] = i[68];
  assign o[35018] = i[68];
  assign o[35019] = i[68];
  assign o[35020] = i[68];
  assign o[35021] = i[68];
  assign o[35022] = i[68];
  assign o[35023] = i[68];
  assign o[35024] = i[68];
  assign o[35025] = i[68];
  assign o[35026] = i[68];
  assign o[35027] = i[68];
  assign o[35028] = i[68];
  assign o[35029] = i[68];
  assign o[35030] = i[68];
  assign o[35031] = i[68];
  assign o[35032] = i[68];
  assign o[35033] = i[68];
  assign o[35034] = i[68];
  assign o[35035] = i[68];
  assign o[35036] = i[68];
  assign o[35037] = i[68];
  assign o[35038] = i[68];
  assign o[35039] = i[68];
  assign o[35040] = i[68];
  assign o[35041] = i[68];
  assign o[35042] = i[68];
  assign o[35043] = i[68];
  assign o[35044] = i[68];
  assign o[35045] = i[68];
  assign o[35046] = i[68];
  assign o[35047] = i[68];
  assign o[35048] = i[68];
  assign o[35049] = i[68];
  assign o[35050] = i[68];
  assign o[35051] = i[68];
  assign o[35052] = i[68];
  assign o[35053] = i[68];
  assign o[35054] = i[68];
  assign o[35055] = i[68];
  assign o[35056] = i[68];
  assign o[35057] = i[68];
  assign o[35058] = i[68];
  assign o[35059] = i[68];
  assign o[35060] = i[68];
  assign o[35061] = i[68];
  assign o[35062] = i[68];
  assign o[35063] = i[68];
  assign o[35064] = i[68];
  assign o[35065] = i[68];
  assign o[35066] = i[68];
  assign o[35067] = i[68];
  assign o[35068] = i[68];
  assign o[35069] = i[68];
  assign o[35070] = i[68];
  assign o[35071] = i[68];
  assign o[35072] = i[68];
  assign o[35073] = i[68];
  assign o[35074] = i[68];
  assign o[35075] = i[68];
  assign o[35076] = i[68];
  assign o[35077] = i[68];
  assign o[35078] = i[68];
  assign o[35079] = i[68];
  assign o[35080] = i[68];
  assign o[35081] = i[68];
  assign o[35082] = i[68];
  assign o[35083] = i[68];
  assign o[35084] = i[68];
  assign o[35085] = i[68];
  assign o[35086] = i[68];
  assign o[35087] = i[68];
  assign o[35088] = i[68];
  assign o[35089] = i[68];
  assign o[35090] = i[68];
  assign o[35091] = i[68];
  assign o[35092] = i[68];
  assign o[35093] = i[68];
  assign o[35094] = i[68];
  assign o[35095] = i[68];
  assign o[35096] = i[68];
  assign o[35097] = i[68];
  assign o[35098] = i[68];
  assign o[35099] = i[68];
  assign o[35100] = i[68];
  assign o[35101] = i[68];
  assign o[35102] = i[68];
  assign o[35103] = i[68];
  assign o[35104] = i[68];
  assign o[35105] = i[68];
  assign o[35106] = i[68];
  assign o[35107] = i[68];
  assign o[35108] = i[68];
  assign o[35109] = i[68];
  assign o[35110] = i[68];
  assign o[35111] = i[68];
  assign o[35112] = i[68];
  assign o[35113] = i[68];
  assign o[35114] = i[68];
  assign o[35115] = i[68];
  assign o[35116] = i[68];
  assign o[35117] = i[68];
  assign o[35118] = i[68];
  assign o[35119] = i[68];
  assign o[35120] = i[68];
  assign o[35121] = i[68];
  assign o[35122] = i[68];
  assign o[35123] = i[68];
  assign o[35124] = i[68];
  assign o[35125] = i[68];
  assign o[35126] = i[68];
  assign o[35127] = i[68];
  assign o[35128] = i[68];
  assign o[35129] = i[68];
  assign o[35130] = i[68];
  assign o[35131] = i[68];
  assign o[35132] = i[68];
  assign o[35133] = i[68];
  assign o[35134] = i[68];
  assign o[35135] = i[68];
  assign o[35136] = i[68];
  assign o[35137] = i[68];
  assign o[35138] = i[68];
  assign o[35139] = i[68];
  assign o[35140] = i[68];
  assign o[35141] = i[68];
  assign o[35142] = i[68];
  assign o[35143] = i[68];
  assign o[35144] = i[68];
  assign o[35145] = i[68];
  assign o[35146] = i[68];
  assign o[35147] = i[68];
  assign o[35148] = i[68];
  assign o[35149] = i[68];
  assign o[35150] = i[68];
  assign o[35151] = i[68];
  assign o[35152] = i[68];
  assign o[35153] = i[68];
  assign o[35154] = i[68];
  assign o[35155] = i[68];
  assign o[35156] = i[68];
  assign o[35157] = i[68];
  assign o[35158] = i[68];
  assign o[35159] = i[68];
  assign o[35160] = i[68];
  assign o[35161] = i[68];
  assign o[35162] = i[68];
  assign o[35163] = i[68];
  assign o[35164] = i[68];
  assign o[35165] = i[68];
  assign o[35166] = i[68];
  assign o[35167] = i[68];
  assign o[35168] = i[68];
  assign o[35169] = i[68];
  assign o[35170] = i[68];
  assign o[35171] = i[68];
  assign o[35172] = i[68];
  assign o[35173] = i[68];
  assign o[35174] = i[68];
  assign o[35175] = i[68];
  assign o[35176] = i[68];
  assign o[35177] = i[68];
  assign o[35178] = i[68];
  assign o[35179] = i[68];
  assign o[35180] = i[68];
  assign o[35181] = i[68];
  assign o[35182] = i[68];
  assign o[35183] = i[68];
  assign o[35184] = i[68];
  assign o[35185] = i[68];
  assign o[35186] = i[68];
  assign o[35187] = i[68];
  assign o[35188] = i[68];
  assign o[35189] = i[68];
  assign o[35190] = i[68];
  assign o[35191] = i[68];
  assign o[35192] = i[68];
  assign o[35193] = i[68];
  assign o[35194] = i[68];
  assign o[35195] = i[68];
  assign o[35196] = i[68];
  assign o[35197] = i[68];
  assign o[35198] = i[68];
  assign o[35199] = i[68];
  assign o[35200] = i[68];
  assign o[35201] = i[68];
  assign o[35202] = i[68];
  assign o[35203] = i[68];
  assign o[35204] = i[68];
  assign o[35205] = i[68];
  assign o[35206] = i[68];
  assign o[35207] = i[68];
  assign o[35208] = i[68];
  assign o[35209] = i[68];
  assign o[35210] = i[68];
  assign o[35211] = i[68];
  assign o[35212] = i[68];
  assign o[35213] = i[68];
  assign o[35214] = i[68];
  assign o[35215] = i[68];
  assign o[35216] = i[68];
  assign o[35217] = i[68];
  assign o[35218] = i[68];
  assign o[35219] = i[68];
  assign o[35220] = i[68];
  assign o[35221] = i[68];
  assign o[35222] = i[68];
  assign o[35223] = i[68];
  assign o[35224] = i[68];
  assign o[35225] = i[68];
  assign o[35226] = i[68];
  assign o[35227] = i[68];
  assign o[35228] = i[68];
  assign o[35229] = i[68];
  assign o[35230] = i[68];
  assign o[35231] = i[68];
  assign o[35232] = i[68];
  assign o[35233] = i[68];
  assign o[35234] = i[68];
  assign o[35235] = i[68];
  assign o[35236] = i[68];
  assign o[35237] = i[68];
  assign o[35238] = i[68];
  assign o[35239] = i[68];
  assign o[35240] = i[68];
  assign o[35241] = i[68];
  assign o[35242] = i[68];
  assign o[35243] = i[68];
  assign o[35244] = i[68];
  assign o[35245] = i[68];
  assign o[35246] = i[68];
  assign o[35247] = i[68];
  assign o[35248] = i[68];
  assign o[35249] = i[68];
  assign o[35250] = i[68];
  assign o[35251] = i[68];
  assign o[35252] = i[68];
  assign o[35253] = i[68];
  assign o[35254] = i[68];
  assign o[35255] = i[68];
  assign o[35256] = i[68];
  assign o[35257] = i[68];
  assign o[35258] = i[68];
  assign o[35259] = i[68];
  assign o[35260] = i[68];
  assign o[35261] = i[68];
  assign o[35262] = i[68];
  assign o[35263] = i[68];
  assign o[35264] = i[68];
  assign o[35265] = i[68];
  assign o[35266] = i[68];
  assign o[35267] = i[68];
  assign o[35268] = i[68];
  assign o[35269] = i[68];
  assign o[35270] = i[68];
  assign o[35271] = i[68];
  assign o[35272] = i[68];
  assign o[35273] = i[68];
  assign o[35274] = i[68];
  assign o[35275] = i[68];
  assign o[35276] = i[68];
  assign o[35277] = i[68];
  assign o[35278] = i[68];
  assign o[35279] = i[68];
  assign o[35280] = i[68];
  assign o[35281] = i[68];
  assign o[35282] = i[68];
  assign o[35283] = i[68];
  assign o[35284] = i[68];
  assign o[35285] = i[68];
  assign o[35286] = i[68];
  assign o[35287] = i[68];
  assign o[35288] = i[68];
  assign o[35289] = i[68];
  assign o[35290] = i[68];
  assign o[35291] = i[68];
  assign o[35292] = i[68];
  assign o[35293] = i[68];
  assign o[35294] = i[68];
  assign o[35295] = i[68];
  assign o[35296] = i[68];
  assign o[35297] = i[68];
  assign o[35298] = i[68];
  assign o[35299] = i[68];
  assign o[35300] = i[68];
  assign o[35301] = i[68];
  assign o[35302] = i[68];
  assign o[35303] = i[68];
  assign o[35304] = i[68];
  assign o[35305] = i[68];
  assign o[35306] = i[68];
  assign o[35307] = i[68];
  assign o[35308] = i[68];
  assign o[35309] = i[68];
  assign o[35310] = i[68];
  assign o[35311] = i[68];
  assign o[35312] = i[68];
  assign o[35313] = i[68];
  assign o[35314] = i[68];
  assign o[35315] = i[68];
  assign o[35316] = i[68];
  assign o[35317] = i[68];
  assign o[35318] = i[68];
  assign o[35319] = i[68];
  assign o[35320] = i[68];
  assign o[35321] = i[68];
  assign o[35322] = i[68];
  assign o[35323] = i[68];
  assign o[35324] = i[68];
  assign o[35325] = i[68];
  assign o[35326] = i[68];
  assign o[35327] = i[68];
  assign o[34304] = i[67];
  assign o[34305] = i[67];
  assign o[34306] = i[67];
  assign o[34307] = i[67];
  assign o[34308] = i[67];
  assign o[34309] = i[67];
  assign o[34310] = i[67];
  assign o[34311] = i[67];
  assign o[34312] = i[67];
  assign o[34313] = i[67];
  assign o[34314] = i[67];
  assign o[34315] = i[67];
  assign o[34316] = i[67];
  assign o[34317] = i[67];
  assign o[34318] = i[67];
  assign o[34319] = i[67];
  assign o[34320] = i[67];
  assign o[34321] = i[67];
  assign o[34322] = i[67];
  assign o[34323] = i[67];
  assign o[34324] = i[67];
  assign o[34325] = i[67];
  assign o[34326] = i[67];
  assign o[34327] = i[67];
  assign o[34328] = i[67];
  assign o[34329] = i[67];
  assign o[34330] = i[67];
  assign o[34331] = i[67];
  assign o[34332] = i[67];
  assign o[34333] = i[67];
  assign o[34334] = i[67];
  assign o[34335] = i[67];
  assign o[34336] = i[67];
  assign o[34337] = i[67];
  assign o[34338] = i[67];
  assign o[34339] = i[67];
  assign o[34340] = i[67];
  assign o[34341] = i[67];
  assign o[34342] = i[67];
  assign o[34343] = i[67];
  assign o[34344] = i[67];
  assign o[34345] = i[67];
  assign o[34346] = i[67];
  assign o[34347] = i[67];
  assign o[34348] = i[67];
  assign o[34349] = i[67];
  assign o[34350] = i[67];
  assign o[34351] = i[67];
  assign o[34352] = i[67];
  assign o[34353] = i[67];
  assign o[34354] = i[67];
  assign o[34355] = i[67];
  assign o[34356] = i[67];
  assign o[34357] = i[67];
  assign o[34358] = i[67];
  assign o[34359] = i[67];
  assign o[34360] = i[67];
  assign o[34361] = i[67];
  assign o[34362] = i[67];
  assign o[34363] = i[67];
  assign o[34364] = i[67];
  assign o[34365] = i[67];
  assign o[34366] = i[67];
  assign o[34367] = i[67];
  assign o[34368] = i[67];
  assign o[34369] = i[67];
  assign o[34370] = i[67];
  assign o[34371] = i[67];
  assign o[34372] = i[67];
  assign o[34373] = i[67];
  assign o[34374] = i[67];
  assign o[34375] = i[67];
  assign o[34376] = i[67];
  assign o[34377] = i[67];
  assign o[34378] = i[67];
  assign o[34379] = i[67];
  assign o[34380] = i[67];
  assign o[34381] = i[67];
  assign o[34382] = i[67];
  assign o[34383] = i[67];
  assign o[34384] = i[67];
  assign o[34385] = i[67];
  assign o[34386] = i[67];
  assign o[34387] = i[67];
  assign o[34388] = i[67];
  assign o[34389] = i[67];
  assign o[34390] = i[67];
  assign o[34391] = i[67];
  assign o[34392] = i[67];
  assign o[34393] = i[67];
  assign o[34394] = i[67];
  assign o[34395] = i[67];
  assign o[34396] = i[67];
  assign o[34397] = i[67];
  assign o[34398] = i[67];
  assign o[34399] = i[67];
  assign o[34400] = i[67];
  assign o[34401] = i[67];
  assign o[34402] = i[67];
  assign o[34403] = i[67];
  assign o[34404] = i[67];
  assign o[34405] = i[67];
  assign o[34406] = i[67];
  assign o[34407] = i[67];
  assign o[34408] = i[67];
  assign o[34409] = i[67];
  assign o[34410] = i[67];
  assign o[34411] = i[67];
  assign o[34412] = i[67];
  assign o[34413] = i[67];
  assign o[34414] = i[67];
  assign o[34415] = i[67];
  assign o[34416] = i[67];
  assign o[34417] = i[67];
  assign o[34418] = i[67];
  assign o[34419] = i[67];
  assign o[34420] = i[67];
  assign o[34421] = i[67];
  assign o[34422] = i[67];
  assign o[34423] = i[67];
  assign o[34424] = i[67];
  assign o[34425] = i[67];
  assign o[34426] = i[67];
  assign o[34427] = i[67];
  assign o[34428] = i[67];
  assign o[34429] = i[67];
  assign o[34430] = i[67];
  assign o[34431] = i[67];
  assign o[34432] = i[67];
  assign o[34433] = i[67];
  assign o[34434] = i[67];
  assign o[34435] = i[67];
  assign o[34436] = i[67];
  assign o[34437] = i[67];
  assign o[34438] = i[67];
  assign o[34439] = i[67];
  assign o[34440] = i[67];
  assign o[34441] = i[67];
  assign o[34442] = i[67];
  assign o[34443] = i[67];
  assign o[34444] = i[67];
  assign o[34445] = i[67];
  assign o[34446] = i[67];
  assign o[34447] = i[67];
  assign o[34448] = i[67];
  assign o[34449] = i[67];
  assign o[34450] = i[67];
  assign o[34451] = i[67];
  assign o[34452] = i[67];
  assign o[34453] = i[67];
  assign o[34454] = i[67];
  assign o[34455] = i[67];
  assign o[34456] = i[67];
  assign o[34457] = i[67];
  assign o[34458] = i[67];
  assign o[34459] = i[67];
  assign o[34460] = i[67];
  assign o[34461] = i[67];
  assign o[34462] = i[67];
  assign o[34463] = i[67];
  assign o[34464] = i[67];
  assign o[34465] = i[67];
  assign o[34466] = i[67];
  assign o[34467] = i[67];
  assign o[34468] = i[67];
  assign o[34469] = i[67];
  assign o[34470] = i[67];
  assign o[34471] = i[67];
  assign o[34472] = i[67];
  assign o[34473] = i[67];
  assign o[34474] = i[67];
  assign o[34475] = i[67];
  assign o[34476] = i[67];
  assign o[34477] = i[67];
  assign o[34478] = i[67];
  assign o[34479] = i[67];
  assign o[34480] = i[67];
  assign o[34481] = i[67];
  assign o[34482] = i[67];
  assign o[34483] = i[67];
  assign o[34484] = i[67];
  assign o[34485] = i[67];
  assign o[34486] = i[67];
  assign o[34487] = i[67];
  assign o[34488] = i[67];
  assign o[34489] = i[67];
  assign o[34490] = i[67];
  assign o[34491] = i[67];
  assign o[34492] = i[67];
  assign o[34493] = i[67];
  assign o[34494] = i[67];
  assign o[34495] = i[67];
  assign o[34496] = i[67];
  assign o[34497] = i[67];
  assign o[34498] = i[67];
  assign o[34499] = i[67];
  assign o[34500] = i[67];
  assign o[34501] = i[67];
  assign o[34502] = i[67];
  assign o[34503] = i[67];
  assign o[34504] = i[67];
  assign o[34505] = i[67];
  assign o[34506] = i[67];
  assign o[34507] = i[67];
  assign o[34508] = i[67];
  assign o[34509] = i[67];
  assign o[34510] = i[67];
  assign o[34511] = i[67];
  assign o[34512] = i[67];
  assign o[34513] = i[67];
  assign o[34514] = i[67];
  assign o[34515] = i[67];
  assign o[34516] = i[67];
  assign o[34517] = i[67];
  assign o[34518] = i[67];
  assign o[34519] = i[67];
  assign o[34520] = i[67];
  assign o[34521] = i[67];
  assign o[34522] = i[67];
  assign o[34523] = i[67];
  assign o[34524] = i[67];
  assign o[34525] = i[67];
  assign o[34526] = i[67];
  assign o[34527] = i[67];
  assign o[34528] = i[67];
  assign o[34529] = i[67];
  assign o[34530] = i[67];
  assign o[34531] = i[67];
  assign o[34532] = i[67];
  assign o[34533] = i[67];
  assign o[34534] = i[67];
  assign o[34535] = i[67];
  assign o[34536] = i[67];
  assign o[34537] = i[67];
  assign o[34538] = i[67];
  assign o[34539] = i[67];
  assign o[34540] = i[67];
  assign o[34541] = i[67];
  assign o[34542] = i[67];
  assign o[34543] = i[67];
  assign o[34544] = i[67];
  assign o[34545] = i[67];
  assign o[34546] = i[67];
  assign o[34547] = i[67];
  assign o[34548] = i[67];
  assign o[34549] = i[67];
  assign o[34550] = i[67];
  assign o[34551] = i[67];
  assign o[34552] = i[67];
  assign o[34553] = i[67];
  assign o[34554] = i[67];
  assign o[34555] = i[67];
  assign o[34556] = i[67];
  assign o[34557] = i[67];
  assign o[34558] = i[67];
  assign o[34559] = i[67];
  assign o[34560] = i[67];
  assign o[34561] = i[67];
  assign o[34562] = i[67];
  assign o[34563] = i[67];
  assign o[34564] = i[67];
  assign o[34565] = i[67];
  assign o[34566] = i[67];
  assign o[34567] = i[67];
  assign o[34568] = i[67];
  assign o[34569] = i[67];
  assign o[34570] = i[67];
  assign o[34571] = i[67];
  assign o[34572] = i[67];
  assign o[34573] = i[67];
  assign o[34574] = i[67];
  assign o[34575] = i[67];
  assign o[34576] = i[67];
  assign o[34577] = i[67];
  assign o[34578] = i[67];
  assign o[34579] = i[67];
  assign o[34580] = i[67];
  assign o[34581] = i[67];
  assign o[34582] = i[67];
  assign o[34583] = i[67];
  assign o[34584] = i[67];
  assign o[34585] = i[67];
  assign o[34586] = i[67];
  assign o[34587] = i[67];
  assign o[34588] = i[67];
  assign o[34589] = i[67];
  assign o[34590] = i[67];
  assign o[34591] = i[67];
  assign o[34592] = i[67];
  assign o[34593] = i[67];
  assign o[34594] = i[67];
  assign o[34595] = i[67];
  assign o[34596] = i[67];
  assign o[34597] = i[67];
  assign o[34598] = i[67];
  assign o[34599] = i[67];
  assign o[34600] = i[67];
  assign o[34601] = i[67];
  assign o[34602] = i[67];
  assign o[34603] = i[67];
  assign o[34604] = i[67];
  assign o[34605] = i[67];
  assign o[34606] = i[67];
  assign o[34607] = i[67];
  assign o[34608] = i[67];
  assign o[34609] = i[67];
  assign o[34610] = i[67];
  assign o[34611] = i[67];
  assign o[34612] = i[67];
  assign o[34613] = i[67];
  assign o[34614] = i[67];
  assign o[34615] = i[67];
  assign o[34616] = i[67];
  assign o[34617] = i[67];
  assign o[34618] = i[67];
  assign o[34619] = i[67];
  assign o[34620] = i[67];
  assign o[34621] = i[67];
  assign o[34622] = i[67];
  assign o[34623] = i[67];
  assign o[34624] = i[67];
  assign o[34625] = i[67];
  assign o[34626] = i[67];
  assign o[34627] = i[67];
  assign o[34628] = i[67];
  assign o[34629] = i[67];
  assign o[34630] = i[67];
  assign o[34631] = i[67];
  assign o[34632] = i[67];
  assign o[34633] = i[67];
  assign o[34634] = i[67];
  assign o[34635] = i[67];
  assign o[34636] = i[67];
  assign o[34637] = i[67];
  assign o[34638] = i[67];
  assign o[34639] = i[67];
  assign o[34640] = i[67];
  assign o[34641] = i[67];
  assign o[34642] = i[67];
  assign o[34643] = i[67];
  assign o[34644] = i[67];
  assign o[34645] = i[67];
  assign o[34646] = i[67];
  assign o[34647] = i[67];
  assign o[34648] = i[67];
  assign o[34649] = i[67];
  assign o[34650] = i[67];
  assign o[34651] = i[67];
  assign o[34652] = i[67];
  assign o[34653] = i[67];
  assign o[34654] = i[67];
  assign o[34655] = i[67];
  assign o[34656] = i[67];
  assign o[34657] = i[67];
  assign o[34658] = i[67];
  assign o[34659] = i[67];
  assign o[34660] = i[67];
  assign o[34661] = i[67];
  assign o[34662] = i[67];
  assign o[34663] = i[67];
  assign o[34664] = i[67];
  assign o[34665] = i[67];
  assign o[34666] = i[67];
  assign o[34667] = i[67];
  assign o[34668] = i[67];
  assign o[34669] = i[67];
  assign o[34670] = i[67];
  assign o[34671] = i[67];
  assign o[34672] = i[67];
  assign o[34673] = i[67];
  assign o[34674] = i[67];
  assign o[34675] = i[67];
  assign o[34676] = i[67];
  assign o[34677] = i[67];
  assign o[34678] = i[67];
  assign o[34679] = i[67];
  assign o[34680] = i[67];
  assign o[34681] = i[67];
  assign o[34682] = i[67];
  assign o[34683] = i[67];
  assign o[34684] = i[67];
  assign o[34685] = i[67];
  assign o[34686] = i[67];
  assign o[34687] = i[67];
  assign o[34688] = i[67];
  assign o[34689] = i[67];
  assign o[34690] = i[67];
  assign o[34691] = i[67];
  assign o[34692] = i[67];
  assign o[34693] = i[67];
  assign o[34694] = i[67];
  assign o[34695] = i[67];
  assign o[34696] = i[67];
  assign o[34697] = i[67];
  assign o[34698] = i[67];
  assign o[34699] = i[67];
  assign o[34700] = i[67];
  assign o[34701] = i[67];
  assign o[34702] = i[67];
  assign o[34703] = i[67];
  assign o[34704] = i[67];
  assign o[34705] = i[67];
  assign o[34706] = i[67];
  assign o[34707] = i[67];
  assign o[34708] = i[67];
  assign o[34709] = i[67];
  assign o[34710] = i[67];
  assign o[34711] = i[67];
  assign o[34712] = i[67];
  assign o[34713] = i[67];
  assign o[34714] = i[67];
  assign o[34715] = i[67];
  assign o[34716] = i[67];
  assign o[34717] = i[67];
  assign o[34718] = i[67];
  assign o[34719] = i[67];
  assign o[34720] = i[67];
  assign o[34721] = i[67];
  assign o[34722] = i[67];
  assign o[34723] = i[67];
  assign o[34724] = i[67];
  assign o[34725] = i[67];
  assign o[34726] = i[67];
  assign o[34727] = i[67];
  assign o[34728] = i[67];
  assign o[34729] = i[67];
  assign o[34730] = i[67];
  assign o[34731] = i[67];
  assign o[34732] = i[67];
  assign o[34733] = i[67];
  assign o[34734] = i[67];
  assign o[34735] = i[67];
  assign o[34736] = i[67];
  assign o[34737] = i[67];
  assign o[34738] = i[67];
  assign o[34739] = i[67];
  assign o[34740] = i[67];
  assign o[34741] = i[67];
  assign o[34742] = i[67];
  assign o[34743] = i[67];
  assign o[34744] = i[67];
  assign o[34745] = i[67];
  assign o[34746] = i[67];
  assign o[34747] = i[67];
  assign o[34748] = i[67];
  assign o[34749] = i[67];
  assign o[34750] = i[67];
  assign o[34751] = i[67];
  assign o[34752] = i[67];
  assign o[34753] = i[67];
  assign o[34754] = i[67];
  assign o[34755] = i[67];
  assign o[34756] = i[67];
  assign o[34757] = i[67];
  assign o[34758] = i[67];
  assign o[34759] = i[67];
  assign o[34760] = i[67];
  assign o[34761] = i[67];
  assign o[34762] = i[67];
  assign o[34763] = i[67];
  assign o[34764] = i[67];
  assign o[34765] = i[67];
  assign o[34766] = i[67];
  assign o[34767] = i[67];
  assign o[34768] = i[67];
  assign o[34769] = i[67];
  assign o[34770] = i[67];
  assign o[34771] = i[67];
  assign o[34772] = i[67];
  assign o[34773] = i[67];
  assign o[34774] = i[67];
  assign o[34775] = i[67];
  assign o[34776] = i[67];
  assign o[34777] = i[67];
  assign o[34778] = i[67];
  assign o[34779] = i[67];
  assign o[34780] = i[67];
  assign o[34781] = i[67];
  assign o[34782] = i[67];
  assign o[34783] = i[67];
  assign o[34784] = i[67];
  assign o[34785] = i[67];
  assign o[34786] = i[67];
  assign o[34787] = i[67];
  assign o[34788] = i[67];
  assign o[34789] = i[67];
  assign o[34790] = i[67];
  assign o[34791] = i[67];
  assign o[34792] = i[67];
  assign o[34793] = i[67];
  assign o[34794] = i[67];
  assign o[34795] = i[67];
  assign o[34796] = i[67];
  assign o[34797] = i[67];
  assign o[34798] = i[67];
  assign o[34799] = i[67];
  assign o[34800] = i[67];
  assign o[34801] = i[67];
  assign o[34802] = i[67];
  assign o[34803] = i[67];
  assign o[34804] = i[67];
  assign o[34805] = i[67];
  assign o[34806] = i[67];
  assign o[34807] = i[67];
  assign o[34808] = i[67];
  assign o[34809] = i[67];
  assign o[34810] = i[67];
  assign o[34811] = i[67];
  assign o[34812] = i[67];
  assign o[34813] = i[67];
  assign o[34814] = i[67];
  assign o[34815] = i[67];
  assign o[33792] = i[66];
  assign o[33793] = i[66];
  assign o[33794] = i[66];
  assign o[33795] = i[66];
  assign o[33796] = i[66];
  assign o[33797] = i[66];
  assign o[33798] = i[66];
  assign o[33799] = i[66];
  assign o[33800] = i[66];
  assign o[33801] = i[66];
  assign o[33802] = i[66];
  assign o[33803] = i[66];
  assign o[33804] = i[66];
  assign o[33805] = i[66];
  assign o[33806] = i[66];
  assign o[33807] = i[66];
  assign o[33808] = i[66];
  assign o[33809] = i[66];
  assign o[33810] = i[66];
  assign o[33811] = i[66];
  assign o[33812] = i[66];
  assign o[33813] = i[66];
  assign o[33814] = i[66];
  assign o[33815] = i[66];
  assign o[33816] = i[66];
  assign o[33817] = i[66];
  assign o[33818] = i[66];
  assign o[33819] = i[66];
  assign o[33820] = i[66];
  assign o[33821] = i[66];
  assign o[33822] = i[66];
  assign o[33823] = i[66];
  assign o[33824] = i[66];
  assign o[33825] = i[66];
  assign o[33826] = i[66];
  assign o[33827] = i[66];
  assign o[33828] = i[66];
  assign o[33829] = i[66];
  assign o[33830] = i[66];
  assign o[33831] = i[66];
  assign o[33832] = i[66];
  assign o[33833] = i[66];
  assign o[33834] = i[66];
  assign o[33835] = i[66];
  assign o[33836] = i[66];
  assign o[33837] = i[66];
  assign o[33838] = i[66];
  assign o[33839] = i[66];
  assign o[33840] = i[66];
  assign o[33841] = i[66];
  assign o[33842] = i[66];
  assign o[33843] = i[66];
  assign o[33844] = i[66];
  assign o[33845] = i[66];
  assign o[33846] = i[66];
  assign o[33847] = i[66];
  assign o[33848] = i[66];
  assign o[33849] = i[66];
  assign o[33850] = i[66];
  assign o[33851] = i[66];
  assign o[33852] = i[66];
  assign o[33853] = i[66];
  assign o[33854] = i[66];
  assign o[33855] = i[66];
  assign o[33856] = i[66];
  assign o[33857] = i[66];
  assign o[33858] = i[66];
  assign o[33859] = i[66];
  assign o[33860] = i[66];
  assign o[33861] = i[66];
  assign o[33862] = i[66];
  assign o[33863] = i[66];
  assign o[33864] = i[66];
  assign o[33865] = i[66];
  assign o[33866] = i[66];
  assign o[33867] = i[66];
  assign o[33868] = i[66];
  assign o[33869] = i[66];
  assign o[33870] = i[66];
  assign o[33871] = i[66];
  assign o[33872] = i[66];
  assign o[33873] = i[66];
  assign o[33874] = i[66];
  assign o[33875] = i[66];
  assign o[33876] = i[66];
  assign o[33877] = i[66];
  assign o[33878] = i[66];
  assign o[33879] = i[66];
  assign o[33880] = i[66];
  assign o[33881] = i[66];
  assign o[33882] = i[66];
  assign o[33883] = i[66];
  assign o[33884] = i[66];
  assign o[33885] = i[66];
  assign o[33886] = i[66];
  assign o[33887] = i[66];
  assign o[33888] = i[66];
  assign o[33889] = i[66];
  assign o[33890] = i[66];
  assign o[33891] = i[66];
  assign o[33892] = i[66];
  assign o[33893] = i[66];
  assign o[33894] = i[66];
  assign o[33895] = i[66];
  assign o[33896] = i[66];
  assign o[33897] = i[66];
  assign o[33898] = i[66];
  assign o[33899] = i[66];
  assign o[33900] = i[66];
  assign o[33901] = i[66];
  assign o[33902] = i[66];
  assign o[33903] = i[66];
  assign o[33904] = i[66];
  assign o[33905] = i[66];
  assign o[33906] = i[66];
  assign o[33907] = i[66];
  assign o[33908] = i[66];
  assign o[33909] = i[66];
  assign o[33910] = i[66];
  assign o[33911] = i[66];
  assign o[33912] = i[66];
  assign o[33913] = i[66];
  assign o[33914] = i[66];
  assign o[33915] = i[66];
  assign o[33916] = i[66];
  assign o[33917] = i[66];
  assign o[33918] = i[66];
  assign o[33919] = i[66];
  assign o[33920] = i[66];
  assign o[33921] = i[66];
  assign o[33922] = i[66];
  assign o[33923] = i[66];
  assign o[33924] = i[66];
  assign o[33925] = i[66];
  assign o[33926] = i[66];
  assign o[33927] = i[66];
  assign o[33928] = i[66];
  assign o[33929] = i[66];
  assign o[33930] = i[66];
  assign o[33931] = i[66];
  assign o[33932] = i[66];
  assign o[33933] = i[66];
  assign o[33934] = i[66];
  assign o[33935] = i[66];
  assign o[33936] = i[66];
  assign o[33937] = i[66];
  assign o[33938] = i[66];
  assign o[33939] = i[66];
  assign o[33940] = i[66];
  assign o[33941] = i[66];
  assign o[33942] = i[66];
  assign o[33943] = i[66];
  assign o[33944] = i[66];
  assign o[33945] = i[66];
  assign o[33946] = i[66];
  assign o[33947] = i[66];
  assign o[33948] = i[66];
  assign o[33949] = i[66];
  assign o[33950] = i[66];
  assign o[33951] = i[66];
  assign o[33952] = i[66];
  assign o[33953] = i[66];
  assign o[33954] = i[66];
  assign o[33955] = i[66];
  assign o[33956] = i[66];
  assign o[33957] = i[66];
  assign o[33958] = i[66];
  assign o[33959] = i[66];
  assign o[33960] = i[66];
  assign o[33961] = i[66];
  assign o[33962] = i[66];
  assign o[33963] = i[66];
  assign o[33964] = i[66];
  assign o[33965] = i[66];
  assign o[33966] = i[66];
  assign o[33967] = i[66];
  assign o[33968] = i[66];
  assign o[33969] = i[66];
  assign o[33970] = i[66];
  assign o[33971] = i[66];
  assign o[33972] = i[66];
  assign o[33973] = i[66];
  assign o[33974] = i[66];
  assign o[33975] = i[66];
  assign o[33976] = i[66];
  assign o[33977] = i[66];
  assign o[33978] = i[66];
  assign o[33979] = i[66];
  assign o[33980] = i[66];
  assign o[33981] = i[66];
  assign o[33982] = i[66];
  assign o[33983] = i[66];
  assign o[33984] = i[66];
  assign o[33985] = i[66];
  assign o[33986] = i[66];
  assign o[33987] = i[66];
  assign o[33988] = i[66];
  assign o[33989] = i[66];
  assign o[33990] = i[66];
  assign o[33991] = i[66];
  assign o[33992] = i[66];
  assign o[33993] = i[66];
  assign o[33994] = i[66];
  assign o[33995] = i[66];
  assign o[33996] = i[66];
  assign o[33997] = i[66];
  assign o[33998] = i[66];
  assign o[33999] = i[66];
  assign o[34000] = i[66];
  assign o[34001] = i[66];
  assign o[34002] = i[66];
  assign o[34003] = i[66];
  assign o[34004] = i[66];
  assign o[34005] = i[66];
  assign o[34006] = i[66];
  assign o[34007] = i[66];
  assign o[34008] = i[66];
  assign o[34009] = i[66];
  assign o[34010] = i[66];
  assign o[34011] = i[66];
  assign o[34012] = i[66];
  assign o[34013] = i[66];
  assign o[34014] = i[66];
  assign o[34015] = i[66];
  assign o[34016] = i[66];
  assign o[34017] = i[66];
  assign o[34018] = i[66];
  assign o[34019] = i[66];
  assign o[34020] = i[66];
  assign o[34021] = i[66];
  assign o[34022] = i[66];
  assign o[34023] = i[66];
  assign o[34024] = i[66];
  assign o[34025] = i[66];
  assign o[34026] = i[66];
  assign o[34027] = i[66];
  assign o[34028] = i[66];
  assign o[34029] = i[66];
  assign o[34030] = i[66];
  assign o[34031] = i[66];
  assign o[34032] = i[66];
  assign o[34033] = i[66];
  assign o[34034] = i[66];
  assign o[34035] = i[66];
  assign o[34036] = i[66];
  assign o[34037] = i[66];
  assign o[34038] = i[66];
  assign o[34039] = i[66];
  assign o[34040] = i[66];
  assign o[34041] = i[66];
  assign o[34042] = i[66];
  assign o[34043] = i[66];
  assign o[34044] = i[66];
  assign o[34045] = i[66];
  assign o[34046] = i[66];
  assign o[34047] = i[66];
  assign o[34048] = i[66];
  assign o[34049] = i[66];
  assign o[34050] = i[66];
  assign o[34051] = i[66];
  assign o[34052] = i[66];
  assign o[34053] = i[66];
  assign o[34054] = i[66];
  assign o[34055] = i[66];
  assign o[34056] = i[66];
  assign o[34057] = i[66];
  assign o[34058] = i[66];
  assign o[34059] = i[66];
  assign o[34060] = i[66];
  assign o[34061] = i[66];
  assign o[34062] = i[66];
  assign o[34063] = i[66];
  assign o[34064] = i[66];
  assign o[34065] = i[66];
  assign o[34066] = i[66];
  assign o[34067] = i[66];
  assign o[34068] = i[66];
  assign o[34069] = i[66];
  assign o[34070] = i[66];
  assign o[34071] = i[66];
  assign o[34072] = i[66];
  assign o[34073] = i[66];
  assign o[34074] = i[66];
  assign o[34075] = i[66];
  assign o[34076] = i[66];
  assign o[34077] = i[66];
  assign o[34078] = i[66];
  assign o[34079] = i[66];
  assign o[34080] = i[66];
  assign o[34081] = i[66];
  assign o[34082] = i[66];
  assign o[34083] = i[66];
  assign o[34084] = i[66];
  assign o[34085] = i[66];
  assign o[34086] = i[66];
  assign o[34087] = i[66];
  assign o[34088] = i[66];
  assign o[34089] = i[66];
  assign o[34090] = i[66];
  assign o[34091] = i[66];
  assign o[34092] = i[66];
  assign o[34093] = i[66];
  assign o[34094] = i[66];
  assign o[34095] = i[66];
  assign o[34096] = i[66];
  assign o[34097] = i[66];
  assign o[34098] = i[66];
  assign o[34099] = i[66];
  assign o[34100] = i[66];
  assign o[34101] = i[66];
  assign o[34102] = i[66];
  assign o[34103] = i[66];
  assign o[34104] = i[66];
  assign o[34105] = i[66];
  assign o[34106] = i[66];
  assign o[34107] = i[66];
  assign o[34108] = i[66];
  assign o[34109] = i[66];
  assign o[34110] = i[66];
  assign o[34111] = i[66];
  assign o[34112] = i[66];
  assign o[34113] = i[66];
  assign o[34114] = i[66];
  assign o[34115] = i[66];
  assign o[34116] = i[66];
  assign o[34117] = i[66];
  assign o[34118] = i[66];
  assign o[34119] = i[66];
  assign o[34120] = i[66];
  assign o[34121] = i[66];
  assign o[34122] = i[66];
  assign o[34123] = i[66];
  assign o[34124] = i[66];
  assign o[34125] = i[66];
  assign o[34126] = i[66];
  assign o[34127] = i[66];
  assign o[34128] = i[66];
  assign o[34129] = i[66];
  assign o[34130] = i[66];
  assign o[34131] = i[66];
  assign o[34132] = i[66];
  assign o[34133] = i[66];
  assign o[34134] = i[66];
  assign o[34135] = i[66];
  assign o[34136] = i[66];
  assign o[34137] = i[66];
  assign o[34138] = i[66];
  assign o[34139] = i[66];
  assign o[34140] = i[66];
  assign o[34141] = i[66];
  assign o[34142] = i[66];
  assign o[34143] = i[66];
  assign o[34144] = i[66];
  assign o[34145] = i[66];
  assign o[34146] = i[66];
  assign o[34147] = i[66];
  assign o[34148] = i[66];
  assign o[34149] = i[66];
  assign o[34150] = i[66];
  assign o[34151] = i[66];
  assign o[34152] = i[66];
  assign o[34153] = i[66];
  assign o[34154] = i[66];
  assign o[34155] = i[66];
  assign o[34156] = i[66];
  assign o[34157] = i[66];
  assign o[34158] = i[66];
  assign o[34159] = i[66];
  assign o[34160] = i[66];
  assign o[34161] = i[66];
  assign o[34162] = i[66];
  assign o[34163] = i[66];
  assign o[34164] = i[66];
  assign o[34165] = i[66];
  assign o[34166] = i[66];
  assign o[34167] = i[66];
  assign o[34168] = i[66];
  assign o[34169] = i[66];
  assign o[34170] = i[66];
  assign o[34171] = i[66];
  assign o[34172] = i[66];
  assign o[34173] = i[66];
  assign o[34174] = i[66];
  assign o[34175] = i[66];
  assign o[34176] = i[66];
  assign o[34177] = i[66];
  assign o[34178] = i[66];
  assign o[34179] = i[66];
  assign o[34180] = i[66];
  assign o[34181] = i[66];
  assign o[34182] = i[66];
  assign o[34183] = i[66];
  assign o[34184] = i[66];
  assign o[34185] = i[66];
  assign o[34186] = i[66];
  assign o[34187] = i[66];
  assign o[34188] = i[66];
  assign o[34189] = i[66];
  assign o[34190] = i[66];
  assign o[34191] = i[66];
  assign o[34192] = i[66];
  assign o[34193] = i[66];
  assign o[34194] = i[66];
  assign o[34195] = i[66];
  assign o[34196] = i[66];
  assign o[34197] = i[66];
  assign o[34198] = i[66];
  assign o[34199] = i[66];
  assign o[34200] = i[66];
  assign o[34201] = i[66];
  assign o[34202] = i[66];
  assign o[34203] = i[66];
  assign o[34204] = i[66];
  assign o[34205] = i[66];
  assign o[34206] = i[66];
  assign o[34207] = i[66];
  assign o[34208] = i[66];
  assign o[34209] = i[66];
  assign o[34210] = i[66];
  assign o[34211] = i[66];
  assign o[34212] = i[66];
  assign o[34213] = i[66];
  assign o[34214] = i[66];
  assign o[34215] = i[66];
  assign o[34216] = i[66];
  assign o[34217] = i[66];
  assign o[34218] = i[66];
  assign o[34219] = i[66];
  assign o[34220] = i[66];
  assign o[34221] = i[66];
  assign o[34222] = i[66];
  assign o[34223] = i[66];
  assign o[34224] = i[66];
  assign o[34225] = i[66];
  assign o[34226] = i[66];
  assign o[34227] = i[66];
  assign o[34228] = i[66];
  assign o[34229] = i[66];
  assign o[34230] = i[66];
  assign o[34231] = i[66];
  assign o[34232] = i[66];
  assign o[34233] = i[66];
  assign o[34234] = i[66];
  assign o[34235] = i[66];
  assign o[34236] = i[66];
  assign o[34237] = i[66];
  assign o[34238] = i[66];
  assign o[34239] = i[66];
  assign o[34240] = i[66];
  assign o[34241] = i[66];
  assign o[34242] = i[66];
  assign o[34243] = i[66];
  assign o[34244] = i[66];
  assign o[34245] = i[66];
  assign o[34246] = i[66];
  assign o[34247] = i[66];
  assign o[34248] = i[66];
  assign o[34249] = i[66];
  assign o[34250] = i[66];
  assign o[34251] = i[66];
  assign o[34252] = i[66];
  assign o[34253] = i[66];
  assign o[34254] = i[66];
  assign o[34255] = i[66];
  assign o[34256] = i[66];
  assign o[34257] = i[66];
  assign o[34258] = i[66];
  assign o[34259] = i[66];
  assign o[34260] = i[66];
  assign o[34261] = i[66];
  assign o[34262] = i[66];
  assign o[34263] = i[66];
  assign o[34264] = i[66];
  assign o[34265] = i[66];
  assign o[34266] = i[66];
  assign o[34267] = i[66];
  assign o[34268] = i[66];
  assign o[34269] = i[66];
  assign o[34270] = i[66];
  assign o[34271] = i[66];
  assign o[34272] = i[66];
  assign o[34273] = i[66];
  assign o[34274] = i[66];
  assign o[34275] = i[66];
  assign o[34276] = i[66];
  assign o[34277] = i[66];
  assign o[34278] = i[66];
  assign o[34279] = i[66];
  assign o[34280] = i[66];
  assign o[34281] = i[66];
  assign o[34282] = i[66];
  assign o[34283] = i[66];
  assign o[34284] = i[66];
  assign o[34285] = i[66];
  assign o[34286] = i[66];
  assign o[34287] = i[66];
  assign o[34288] = i[66];
  assign o[34289] = i[66];
  assign o[34290] = i[66];
  assign o[34291] = i[66];
  assign o[34292] = i[66];
  assign o[34293] = i[66];
  assign o[34294] = i[66];
  assign o[34295] = i[66];
  assign o[34296] = i[66];
  assign o[34297] = i[66];
  assign o[34298] = i[66];
  assign o[34299] = i[66];
  assign o[34300] = i[66];
  assign o[34301] = i[66];
  assign o[34302] = i[66];
  assign o[34303] = i[66];
  assign o[33280] = i[65];
  assign o[33281] = i[65];
  assign o[33282] = i[65];
  assign o[33283] = i[65];
  assign o[33284] = i[65];
  assign o[33285] = i[65];
  assign o[33286] = i[65];
  assign o[33287] = i[65];
  assign o[33288] = i[65];
  assign o[33289] = i[65];
  assign o[33290] = i[65];
  assign o[33291] = i[65];
  assign o[33292] = i[65];
  assign o[33293] = i[65];
  assign o[33294] = i[65];
  assign o[33295] = i[65];
  assign o[33296] = i[65];
  assign o[33297] = i[65];
  assign o[33298] = i[65];
  assign o[33299] = i[65];
  assign o[33300] = i[65];
  assign o[33301] = i[65];
  assign o[33302] = i[65];
  assign o[33303] = i[65];
  assign o[33304] = i[65];
  assign o[33305] = i[65];
  assign o[33306] = i[65];
  assign o[33307] = i[65];
  assign o[33308] = i[65];
  assign o[33309] = i[65];
  assign o[33310] = i[65];
  assign o[33311] = i[65];
  assign o[33312] = i[65];
  assign o[33313] = i[65];
  assign o[33314] = i[65];
  assign o[33315] = i[65];
  assign o[33316] = i[65];
  assign o[33317] = i[65];
  assign o[33318] = i[65];
  assign o[33319] = i[65];
  assign o[33320] = i[65];
  assign o[33321] = i[65];
  assign o[33322] = i[65];
  assign o[33323] = i[65];
  assign o[33324] = i[65];
  assign o[33325] = i[65];
  assign o[33326] = i[65];
  assign o[33327] = i[65];
  assign o[33328] = i[65];
  assign o[33329] = i[65];
  assign o[33330] = i[65];
  assign o[33331] = i[65];
  assign o[33332] = i[65];
  assign o[33333] = i[65];
  assign o[33334] = i[65];
  assign o[33335] = i[65];
  assign o[33336] = i[65];
  assign o[33337] = i[65];
  assign o[33338] = i[65];
  assign o[33339] = i[65];
  assign o[33340] = i[65];
  assign o[33341] = i[65];
  assign o[33342] = i[65];
  assign o[33343] = i[65];
  assign o[33344] = i[65];
  assign o[33345] = i[65];
  assign o[33346] = i[65];
  assign o[33347] = i[65];
  assign o[33348] = i[65];
  assign o[33349] = i[65];
  assign o[33350] = i[65];
  assign o[33351] = i[65];
  assign o[33352] = i[65];
  assign o[33353] = i[65];
  assign o[33354] = i[65];
  assign o[33355] = i[65];
  assign o[33356] = i[65];
  assign o[33357] = i[65];
  assign o[33358] = i[65];
  assign o[33359] = i[65];
  assign o[33360] = i[65];
  assign o[33361] = i[65];
  assign o[33362] = i[65];
  assign o[33363] = i[65];
  assign o[33364] = i[65];
  assign o[33365] = i[65];
  assign o[33366] = i[65];
  assign o[33367] = i[65];
  assign o[33368] = i[65];
  assign o[33369] = i[65];
  assign o[33370] = i[65];
  assign o[33371] = i[65];
  assign o[33372] = i[65];
  assign o[33373] = i[65];
  assign o[33374] = i[65];
  assign o[33375] = i[65];
  assign o[33376] = i[65];
  assign o[33377] = i[65];
  assign o[33378] = i[65];
  assign o[33379] = i[65];
  assign o[33380] = i[65];
  assign o[33381] = i[65];
  assign o[33382] = i[65];
  assign o[33383] = i[65];
  assign o[33384] = i[65];
  assign o[33385] = i[65];
  assign o[33386] = i[65];
  assign o[33387] = i[65];
  assign o[33388] = i[65];
  assign o[33389] = i[65];
  assign o[33390] = i[65];
  assign o[33391] = i[65];
  assign o[33392] = i[65];
  assign o[33393] = i[65];
  assign o[33394] = i[65];
  assign o[33395] = i[65];
  assign o[33396] = i[65];
  assign o[33397] = i[65];
  assign o[33398] = i[65];
  assign o[33399] = i[65];
  assign o[33400] = i[65];
  assign o[33401] = i[65];
  assign o[33402] = i[65];
  assign o[33403] = i[65];
  assign o[33404] = i[65];
  assign o[33405] = i[65];
  assign o[33406] = i[65];
  assign o[33407] = i[65];
  assign o[33408] = i[65];
  assign o[33409] = i[65];
  assign o[33410] = i[65];
  assign o[33411] = i[65];
  assign o[33412] = i[65];
  assign o[33413] = i[65];
  assign o[33414] = i[65];
  assign o[33415] = i[65];
  assign o[33416] = i[65];
  assign o[33417] = i[65];
  assign o[33418] = i[65];
  assign o[33419] = i[65];
  assign o[33420] = i[65];
  assign o[33421] = i[65];
  assign o[33422] = i[65];
  assign o[33423] = i[65];
  assign o[33424] = i[65];
  assign o[33425] = i[65];
  assign o[33426] = i[65];
  assign o[33427] = i[65];
  assign o[33428] = i[65];
  assign o[33429] = i[65];
  assign o[33430] = i[65];
  assign o[33431] = i[65];
  assign o[33432] = i[65];
  assign o[33433] = i[65];
  assign o[33434] = i[65];
  assign o[33435] = i[65];
  assign o[33436] = i[65];
  assign o[33437] = i[65];
  assign o[33438] = i[65];
  assign o[33439] = i[65];
  assign o[33440] = i[65];
  assign o[33441] = i[65];
  assign o[33442] = i[65];
  assign o[33443] = i[65];
  assign o[33444] = i[65];
  assign o[33445] = i[65];
  assign o[33446] = i[65];
  assign o[33447] = i[65];
  assign o[33448] = i[65];
  assign o[33449] = i[65];
  assign o[33450] = i[65];
  assign o[33451] = i[65];
  assign o[33452] = i[65];
  assign o[33453] = i[65];
  assign o[33454] = i[65];
  assign o[33455] = i[65];
  assign o[33456] = i[65];
  assign o[33457] = i[65];
  assign o[33458] = i[65];
  assign o[33459] = i[65];
  assign o[33460] = i[65];
  assign o[33461] = i[65];
  assign o[33462] = i[65];
  assign o[33463] = i[65];
  assign o[33464] = i[65];
  assign o[33465] = i[65];
  assign o[33466] = i[65];
  assign o[33467] = i[65];
  assign o[33468] = i[65];
  assign o[33469] = i[65];
  assign o[33470] = i[65];
  assign o[33471] = i[65];
  assign o[33472] = i[65];
  assign o[33473] = i[65];
  assign o[33474] = i[65];
  assign o[33475] = i[65];
  assign o[33476] = i[65];
  assign o[33477] = i[65];
  assign o[33478] = i[65];
  assign o[33479] = i[65];
  assign o[33480] = i[65];
  assign o[33481] = i[65];
  assign o[33482] = i[65];
  assign o[33483] = i[65];
  assign o[33484] = i[65];
  assign o[33485] = i[65];
  assign o[33486] = i[65];
  assign o[33487] = i[65];
  assign o[33488] = i[65];
  assign o[33489] = i[65];
  assign o[33490] = i[65];
  assign o[33491] = i[65];
  assign o[33492] = i[65];
  assign o[33493] = i[65];
  assign o[33494] = i[65];
  assign o[33495] = i[65];
  assign o[33496] = i[65];
  assign o[33497] = i[65];
  assign o[33498] = i[65];
  assign o[33499] = i[65];
  assign o[33500] = i[65];
  assign o[33501] = i[65];
  assign o[33502] = i[65];
  assign o[33503] = i[65];
  assign o[33504] = i[65];
  assign o[33505] = i[65];
  assign o[33506] = i[65];
  assign o[33507] = i[65];
  assign o[33508] = i[65];
  assign o[33509] = i[65];
  assign o[33510] = i[65];
  assign o[33511] = i[65];
  assign o[33512] = i[65];
  assign o[33513] = i[65];
  assign o[33514] = i[65];
  assign o[33515] = i[65];
  assign o[33516] = i[65];
  assign o[33517] = i[65];
  assign o[33518] = i[65];
  assign o[33519] = i[65];
  assign o[33520] = i[65];
  assign o[33521] = i[65];
  assign o[33522] = i[65];
  assign o[33523] = i[65];
  assign o[33524] = i[65];
  assign o[33525] = i[65];
  assign o[33526] = i[65];
  assign o[33527] = i[65];
  assign o[33528] = i[65];
  assign o[33529] = i[65];
  assign o[33530] = i[65];
  assign o[33531] = i[65];
  assign o[33532] = i[65];
  assign o[33533] = i[65];
  assign o[33534] = i[65];
  assign o[33535] = i[65];
  assign o[33536] = i[65];
  assign o[33537] = i[65];
  assign o[33538] = i[65];
  assign o[33539] = i[65];
  assign o[33540] = i[65];
  assign o[33541] = i[65];
  assign o[33542] = i[65];
  assign o[33543] = i[65];
  assign o[33544] = i[65];
  assign o[33545] = i[65];
  assign o[33546] = i[65];
  assign o[33547] = i[65];
  assign o[33548] = i[65];
  assign o[33549] = i[65];
  assign o[33550] = i[65];
  assign o[33551] = i[65];
  assign o[33552] = i[65];
  assign o[33553] = i[65];
  assign o[33554] = i[65];
  assign o[33555] = i[65];
  assign o[33556] = i[65];
  assign o[33557] = i[65];
  assign o[33558] = i[65];
  assign o[33559] = i[65];
  assign o[33560] = i[65];
  assign o[33561] = i[65];
  assign o[33562] = i[65];
  assign o[33563] = i[65];
  assign o[33564] = i[65];
  assign o[33565] = i[65];
  assign o[33566] = i[65];
  assign o[33567] = i[65];
  assign o[33568] = i[65];
  assign o[33569] = i[65];
  assign o[33570] = i[65];
  assign o[33571] = i[65];
  assign o[33572] = i[65];
  assign o[33573] = i[65];
  assign o[33574] = i[65];
  assign o[33575] = i[65];
  assign o[33576] = i[65];
  assign o[33577] = i[65];
  assign o[33578] = i[65];
  assign o[33579] = i[65];
  assign o[33580] = i[65];
  assign o[33581] = i[65];
  assign o[33582] = i[65];
  assign o[33583] = i[65];
  assign o[33584] = i[65];
  assign o[33585] = i[65];
  assign o[33586] = i[65];
  assign o[33587] = i[65];
  assign o[33588] = i[65];
  assign o[33589] = i[65];
  assign o[33590] = i[65];
  assign o[33591] = i[65];
  assign o[33592] = i[65];
  assign o[33593] = i[65];
  assign o[33594] = i[65];
  assign o[33595] = i[65];
  assign o[33596] = i[65];
  assign o[33597] = i[65];
  assign o[33598] = i[65];
  assign o[33599] = i[65];
  assign o[33600] = i[65];
  assign o[33601] = i[65];
  assign o[33602] = i[65];
  assign o[33603] = i[65];
  assign o[33604] = i[65];
  assign o[33605] = i[65];
  assign o[33606] = i[65];
  assign o[33607] = i[65];
  assign o[33608] = i[65];
  assign o[33609] = i[65];
  assign o[33610] = i[65];
  assign o[33611] = i[65];
  assign o[33612] = i[65];
  assign o[33613] = i[65];
  assign o[33614] = i[65];
  assign o[33615] = i[65];
  assign o[33616] = i[65];
  assign o[33617] = i[65];
  assign o[33618] = i[65];
  assign o[33619] = i[65];
  assign o[33620] = i[65];
  assign o[33621] = i[65];
  assign o[33622] = i[65];
  assign o[33623] = i[65];
  assign o[33624] = i[65];
  assign o[33625] = i[65];
  assign o[33626] = i[65];
  assign o[33627] = i[65];
  assign o[33628] = i[65];
  assign o[33629] = i[65];
  assign o[33630] = i[65];
  assign o[33631] = i[65];
  assign o[33632] = i[65];
  assign o[33633] = i[65];
  assign o[33634] = i[65];
  assign o[33635] = i[65];
  assign o[33636] = i[65];
  assign o[33637] = i[65];
  assign o[33638] = i[65];
  assign o[33639] = i[65];
  assign o[33640] = i[65];
  assign o[33641] = i[65];
  assign o[33642] = i[65];
  assign o[33643] = i[65];
  assign o[33644] = i[65];
  assign o[33645] = i[65];
  assign o[33646] = i[65];
  assign o[33647] = i[65];
  assign o[33648] = i[65];
  assign o[33649] = i[65];
  assign o[33650] = i[65];
  assign o[33651] = i[65];
  assign o[33652] = i[65];
  assign o[33653] = i[65];
  assign o[33654] = i[65];
  assign o[33655] = i[65];
  assign o[33656] = i[65];
  assign o[33657] = i[65];
  assign o[33658] = i[65];
  assign o[33659] = i[65];
  assign o[33660] = i[65];
  assign o[33661] = i[65];
  assign o[33662] = i[65];
  assign o[33663] = i[65];
  assign o[33664] = i[65];
  assign o[33665] = i[65];
  assign o[33666] = i[65];
  assign o[33667] = i[65];
  assign o[33668] = i[65];
  assign o[33669] = i[65];
  assign o[33670] = i[65];
  assign o[33671] = i[65];
  assign o[33672] = i[65];
  assign o[33673] = i[65];
  assign o[33674] = i[65];
  assign o[33675] = i[65];
  assign o[33676] = i[65];
  assign o[33677] = i[65];
  assign o[33678] = i[65];
  assign o[33679] = i[65];
  assign o[33680] = i[65];
  assign o[33681] = i[65];
  assign o[33682] = i[65];
  assign o[33683] = i[65];
  assign o[33684] = i[65];
  assign o[33685] = i[65];
  assign o[33686] = i[65];
  assign o[33687] = i[65];
  assign o[33688] = i[65];
  assign o[33689] = i[65];
  assign o[33690] = i[65];
  assign o[33691] = i[65];
  assign o[33692] = i[65];
  assign o[33693] = i[65];
  assign o[33694] = i[65];
  assign o[33695] = i[65];
  assign o[33696] = i[65];
  assign o[33697] = i[65];
  assign o[33698] = i[65];
  assign o[33699] = i[65];
  assign o[33700] = i[65];
  assign o[33701] = i[65];
  assign o[33702] = i[65];
  assign o[33703] = i[65];
  assign o[33704] = i[65];
  assign o[33705] = i[65];
  assign o[33706] = i[65];
  assign o[33707] = i[65];
  assign o[33708] = i[65];
  assign o[33709] = i[65];
  assign o[33710] = i[65];
  assign o[33711] = i[65];
  assign o[33712] = i[65];
  assign o[33713] = i[65];
  assign o[33714] = i[65];
  assign o[33715] = i[65];
  assign o[33716] = i[65];
  assign o[33717] = i[65];
  assign o[33718] = i[65];
  assign o[33719] = i[65];
  assign o[33720] = i[65];
  assign o[33721] = i[65];
  assign o[33722] = i[65];
  assign o[33723] = i[65];
  assign o[33724] = i[65];
  assign o[33725] = i[65];
  assign o[33726] = i[65];
  assign o[33727] = i[65];
  assign o[33728] = i[65];
  assign o[33729] = i[65];
  assign o[33730] = i[65];
  assign o[33731] = i[65];
  assign o[33732] = i[65];
  assign o[33733] = i[65];
  assign o[33734] = i[65];
  assign o[33735] = i[65];
  assign o[33736] = i[65];
  assign o[33737] = i[65];
  assign o[33738] = i[65];
  assign o[33739] = i[65];
  assign o[33740] = i[65];
  assign o[33741] = i[65];
  assign o[33742] = i[65];
  assign o[33743] = i[65];
  assign o[33744] = i[65];
  assign o[33745] = i[65];
  assign o[33746] = i[65];
  assign o[33747] = i[65];
  assign o[33748] = i[65];
  assign o[33749] = i[65];
  assign o[33750] = i[65];
  assign o[33751] = i[65];
  assign o[33752] = i[65];
  assign o[33753] = i[65];
  assign o[33754] = i[65];
  assign o[33755] = i[65];
  assign o[33756] = i[65];
  assign o[33757] = i[65];
  assign o[33758] = i[65];
  assign o[33759] = i[65];
  assign o[33760] = i[65];
  assign o[33761] = i[65];
  assign o[33762] = i[65];
  assign o[33763] = i[65];
  assign o[33764] = i[65];
  assign o[33765] = i[65];
  assign o[33766] = i[65];
  assign o[33767] = i[65];
  assign o[33768] = i[65];
  assign o[33769] = i[65];
  assign o[33770] = i[65];
  assign o[33771] = i[65];
  assign o[33772] = i[65];
  assign o[33773] = i[65];
  assign o[33774] = i[65];
  assign o[33775] = i[65];
  assign o[33776] = i[65];
  assign o[33777] = i[65];
  assign o[33778] = i[65];
  assign o[33779] = i[65];
  assign o[33780] = i[65];
  assign o[33781] = i[65];
  assign o[33782] = i[65];
  assign o[33783] = i[65];
  assign o[33784] = i[65];
  assign o[33785] = i[65];
  assign o[33786] = i[65];
  assign o[33787] = i[65];
  assign o[33788] = i[65];
  assign o[33789] = i[65];
  assign o[33790] = i[65];
  assign o[33791] = i[65];
  assign o[32768] = i[64];
  assign o[32769] = i[64];
  assign o[32770] = i[64];
  assign o[32771] = i[64];
  assign o[32772] = i[64];
  assign o[32773] = i[64];
  assign o[32774] = i[64];
  assign o[32775] = i[64];
  assign o[32776] = i[64];
  assign o[32777] = i[64];
  assign o[32778] = i[64];
  assign o[32779] = i[64];
  assign o[32780] = i[64];
  assign o[32781] = i[64];
  assign o[32782] = i[64];
  assign o[32783] = i[64];
  assign o[32784] = i[64];
  assign o[32785] = i[64];
  assign o[32786] = i[64];
  assign o[32787] = i[64];
  assign o[32788] = i[64];
  assign o[32789] = i[64];
  assign o[32790] = i[64];
  assign o[32791] = i[64];
  assign o[32792] = i[64];
  assign o[32793] = i[64];
  assign o[32794] = i[64];
  assign o[32795] = i[64];
  assign o[32796] = i[64];
  assign o[32797] = i[64];
  assign o[32798] = i[64];
  assign o[32799] = i[64];
  assign o[32800] = i[64];
  assign o[32801] = i[64];
  assign o[32802] = i[64];
  assign o[32803] = i[64];
  assign o[32804] = i[64];
  assign o[32805] = i[64];
  assign o[32806] = i[64];
  assign o[32807] = i[64];
  assign o[32808] = i[64];
  assign o[32809] = i[64];
  assign o[32810] = i[64];
  assign o[32811] = i[64];
  assign o[32812] = i[64];
  assign o[32813] = i[64];
  assign o[32814] = i[64];
  assign o[32815] = i[64];
  assign o[32816] = i[64];
  assign o[32817] = i[64];
  assign o[32818] = i[64];
  assign o[32819] = i[64];
  assign o[32820] = i[64];
  assign o[32821] = i[64];
  assign o[32822] = i[64];
  assign o[32823] = i[64];
  assign o[32824] = i[64];
  assign o[32825] = i[64];
  assign o[32826] = i[64];
  assign o[32827] = i[64];
  assign o[32828] = i[64];
  assign o[32829] = i[64];
  assign o[32830] = i[64];
  assign o[32831] = i[64];
  assign o[32832] = i[64];
  assign o[32833] = i[64];
  assign o[32834] = i[64];
  assign o[32835] = i[64];
  assign o[32836] = i[64];
  assign o[32837] = i[64];
  assign o[32838] = i[64];
  assign o[32839] = i[64];
  assign o[32840] = i[64];
  assign o[32841] = i[64];
  assign o[32842] = i[64];
  assign o[32843] = i[64];
  assign o[32844] = i[64];
  assign o[32845] = i[64];
  assign o[32846] = i[64];
  assign o[32847] = i[64];
  assign o[32848] = i[64];
  assign o[32849] = i[64];
  assign o[32850] = i[64];
  assign o[32851] = i[64];
  assign o[32852] = i[64];
  assign o[32853] = i[64];
  assign o[32854] = i[64];
  assign o[32855] = i[64];
  assign o[32856] = i[64];
  assign o[32857] = i[64];
  assign o[32858] = i[64];
  assign o[32859] = i[64];
  assign o[32860] = i[64];
  assign o[32861] = i[64];
  assign o[32862] = i[64];
  assign o[32863] = i[64];
  assign o[32864] = i[64];
  assign o[32865] = i[64];
  assign o[32866] = i[64];
  assign o[32867] = i[64];
  assign o[32868] = i[64];
  assign o[32869] = i[64];
  assign o[32870] = i[64];
  assign o[32871] = i[64];
  assign o[32872] = i[64];
  assign o[32873] = i[64];
  assign o[32874] = i[64];
  assign o[32875] = i[64];
  assign o[32876] = i[64];
  assign o[32877] = i[64];
  assign o[32878] = i[64];
  assign o[32879] = i[64];
  assign o[32880] = i[64];
  assign o[32881] = i[64];
  assign o[32882] = i[64];
  assign o[32883] = i[64];
  assign o[32884] = i[64];
  assign o[32885] = i[64];
  assign o[32886] = i[64];
  assign o[32887] = i[64];
  assign o[32888] = i[64];
  assign o[32889] = i[64];
  assign o[32890] = i[64];
  assign o[32891] = i[64];
  assign o[32892] = i[64];
  assign o[32893] = i[64];
  assign o[32894] = i[64];
  assign o[32895] = i[64];
  assign o[32896] = i[64];
  assign o[32897] = i[64];
  assign o[32898] = i[64];
  assign o[32899] = i[64];
  assign o[32900] = i[64];
  assign o[32901] = i[64];
  assign o[32902] = i[64];
  assign o[32903] = i[64];
  assign o[32904] = i[64];
  assign o[32905] = i[64];
  assign o[32906] = i[64];
  assign o[32907] = i[64];
  assign o[32908] = i[64];
  assign o[32909] = i[64];
  assign o[32910] = i[64];
  assign o[32911] = i[64];
  assign o[32912] = i[64];
  assign o[32913] = i[64];
  assign o[32914] = i[64];
  assign o[32915] = i[64];
  assign o[32916] = i[64];
  assign o[32917] = i[64];
  assign o[32918] = i[64];
  assign o[32919] = i[64];
  assign o[32920] = i[64];
  assign o[32921] = i[64];
  assign o[32922] = i[64];
  assign o[32923] = i[64];
  assign o[32924] = i[64];
  assign o[32925] = i[64];
  assign o[32926] = i[64];
  assign o[32927] = i[64];
  assign o[32928] = i[64];
  assign o[32929] = i[64];
  assign o[32930] = i[64];
  assign o[32931] = i[64];
  assign o[32932] = i[64];
  assign o[32933] = i[64];
  assign o[32934] = i[64];
  assign o[32935] = i[64];
  assign o[32936] = i[64];
  assign o[32937] = i[64];
  assign o[32938] = i[64];
  assign o[32939] = i[64];
  assign o[32940] = i[64];
  assign o[32941] = i[64];
  assign o[32942] = i[64];
  assign o[32943] = i[64];
  assign o[32944] = i[64];
  assign o[32945] = i[64];
  assign o[32946] = i[64];
  assign o[32947] = i[64];
  assign o[32948] = i[64];
  assign o[32949] = i[64];
  assign o[32950] = i[64];
  assign o[32951] = i[64];
  assign o[32952] = i[64];
  assign o[32953] = i[64];
  assign o[32954] = i[64];
  assign o[32955] = i[64];
  assign o[32956] = i[64];
  assign o[32957] = i[64];
  assign o[32958] = i[64];
  assign o[32959] = i[64];
  assign o[32960] = i[64];
  assign o[32961] = i[64];
  assign o[32962] = i[64];
  assign o[32963] = i[64];
  assign o[32964] = i[64];
  assign o[32965] = i[64];
  assign o[32966] = i[64];
  assign o[32967] = i[64];
  assign o[32968] = i[64];
  assign o[32969] = i[64];
  assign o[32970] = i[64];
  assign o[32971] = i[64];
  assign o[32972] = i[64];
  assign o[32973] = i[64];
  assign o[32974] = i[64];
  assign o[32975] = i[64];
  assign o[32976] = i[64];
  assign o[32977] = i[64];
  assign o[32978] = i[64];
  assign o[32979] = i[64];
  assign o[32980] = i[64];
  assign o[32981] = i[64];
  assign o[32982] = i[64];
  assign o[32983] = i[64];
  assign o[32984] = i[64];
  assign o[32985] = i[64];
  assign o[32986] = i[64];
  assign o[32987] = i[64];
  assign o[32988] = i[64];
  assign o[32989] = i[64];
  assign o[32990] = i[64];
  assign o[32991] = i[64];
  assign o[32992] = i[64];
  assign o[32993] = i[64];
  assign o[32994] = i[64];
  assign o[32995] = i[64];
  assign o[32996] = i[64];
  assign o[32997] = i[64];
  assign o[32998] = i[64];
  assign o[32999] = i[64];
  assign o[33000] = i[64];
  assign o[33001] = i[64];
  assign o[33002] = i[64];
  assign o[33003] = i[64];
  assign o[33004] = i[64];
  assign o[33005] = i[64];
  assign o[33006] = i[64];
  assign o[33007] = i[64];
  assign o[33008] = i[64];
  assign o[33009] = i[64];
  assign o[33010] = i[64];
  assign o[33011] = i[64];
  assign o[33012] = i[64];
  assign o[33013] = i[64];
  assign o[33014] = i[64];
  assign o[33015] = i[64];
  assign o[33016] = i[64];
  assign o[33017] = i[64];
  assign o[33018] = i[64];
  assign o[33019] = i[64];
  assign o[33020] = i[64];
  assign o[33021] = i[64];
  assign o[33022] = i[64];
  assign o[33023] = i[64];
  assign o[33024] = i[64];
  assign o[33025] = i[64];
  assign o[33026] = i[64];
  assign o[33027] = i[64];
  assign o[33028] = i[64];
  assign o[33029] = i[64];
  assign o[33030] = i[64];
  assign o[33031] = i[64];
  assign o[33032] = i[64];
  assign o[33033] = i[64];
  assign o[33034] = i[64];
  assign o[33035] = i[64];
  assign o[33036] = i[64];
  assign o[33037] = i[64];
  assign o[33038] = i[64];
  assign o[33039] = i[64];
  assign o[33040] = i[64];
  assign o[33041] = i[64];
  assign o[33042] = i[64];
  assign o[33043] = i[64];
  assign o[33044] = i[64];
  assign o[33045] = i[64];
  assign o[33046] = i[64];
  assign o[33047] = i[64];
  assign o[33048] = i[64];
  assign o[33049] = i[64];
  assign o[33050] = i[64];
  assign o[33051] = i[64];
  assign o[33052] = i[64];
  assign o[33053] = i[64];
  assign o[33054] = i[64];
  assign o[33055] = i[64];
  assign o[33056] = i[64];
  assign o[33057] = i[64];
  assign o[33058] = i[64];
  assign o[33059] = i[64];
  assign o[33060] = i[64];
  assign o[33061] = i[64];
  assign o[33062] = i[64];
  assign o[33063] = i[64];
  assign o[33064] = i[64];
  assign o[33065] = i[64];
  assign o[33066] = i[64];
  assign o[33067] = i[64];
  assign o[33068] = i[64];
  assign o[33069] = i[64];
  assign o[33070] = i[64];
  assign o[33071] = i[64];
  assign o[33072] = i[64];
  assign o[33073] = i[64];
  assign o[33074] = i[64];
  assign o[33075] = i[64];
  assign o[33076] = i[64];
  assign o[33077] = i[64];
  assign o[33078] = i[64];
  assign o[33079] = i[64];
  assign o[33080] = i[64];
  assign o[33081] = i[64];
  assign o[33082] = i[64];
  assign o[33083] = i[64];
  assign o[33084] = i[64];
  assign o[33085] = i[64];
  assign o[33086] = i[64];
  assign o[33087] = i[64];
  assign o[33088] = i[64];
  assign o[33089] = i[64];
  assign o[33090] = i[64];
  assign o[33091] = i[64];
  assign o[33092] = i[64];
  assign o[33093] = i[64];
  assign o[33094] = i[64];
  assign o[33095] = i[64];
  assign o[33096] = i[64];
  assign o[33097] = i[64];
  assign o[33098] = i[64];
  assign o[33099] = i[64];
  assign o[33100] = i[64];
  assign o[33101] = i[64];
  assign o[33102] = i[64];
  assign o[33103] = i[64];
  assign o[33104] = i[64];
  assign o[33105] = i[64];
  assign o[33106] = i[64];
  assign o[33107] = i[64];
  assign o[33108] = i[64];
  assign o[33109] = i[64];
  assign o[33110] = i[64];
  assign o[33111] = i[64];
  assign o[33112] = i[64];
  assign o[33113] = i[64];
  assign o[33114] = i[64];
  assign o[33115] = i[64];
  assign o[33116] = i[64];
  assign o[33117] = i[64];
  assign o[33118] = i[64];
  assign o[33119] = i[64];
  assign o[33120] = i[64];
  assign o[33121] = i[64];
  assign o[33122] = i[64];
  assign o[33123] = i[64];
  assign o[33124] = i[64];
  assign o[33125] = i[64];
  assign o[33126] = i[64];
  assign o[33127] = i[64];
  assign o[33128] = i[64];
  assign o[33129] = i[64];
  assign o[33130] = i[64];
  assign o[33131] = i[64];
  assign o[33132] = i[64];
  assign o[33133] = i[64];
  assign o[33134] = i[64];
  assign o[33135] = i[64];
  assign o[33136] = i[64];
  assign o[33137] = i[64];
  assign o[33138] = i[64];
  assign o[33139] = i[64];
  assign o[33140] = i[64];
  assign o[33141] = i[64];
  assign o[33142] = i[64];
  assign o[33143] = i[64];
  assign o[33144] = i[64];
  assign o[33145] = i[64];
  assign o[33146] = i[64];
  assign o[33147] = i[64];
  assign o[33148] = i[64];
  assign o[33149] = i[64];
  assign o[33150] = i[64];
  assign o[33151] = i[64];
  assign o[33152] = i[64];
  assign o[33153] = i[64];
  assign o[33154] = i[64];
  assign o[33155] = i[64];
  assign o[33156] = i[64];
  assign o[33157] = i[64];
  assign o[33158] = i[64];
  assign o[33159] = i[64];
  assign o[33160] = i[64];
  assign o[33161] = i[64];
  assign o[33162] = i[64];
  assign o[33163] = i[64];
  assign o[33164] = i[64];
  assign o[33165] = i[64];
  assign o[33166] = i[64];
  assign o[33167] = i[64];
  assign o[33168] = i[64];
  assign o[33169] = i[64];
  assign o[33170] = i[64];
  assign o[33171] = i[64];
  assign o[33172] = i[64];
  assign o[33173] = i[64];
  assign o[33174] = i[64];
  assign o[33175] = i[64];
  assign o[33176] = i[64];
  assign o[33177] = i[64];
  assign o[33178] = i[64];
  assign o[33179] = i[64];
  assign o[33180] = i[64];
  assign o[33181] = i[64];
  assign o[33182] = i[64];
  assign o[33183] = i[64];
  assign o[33184] = i[64];
  assign o[33185] = i[64];
  assign o[33186] = i[64];
  assign o[33187] = i[64];
  assign o[33188] = i[64];
  assign o[33189] = i[64];
  assign o[33190] = i[64];
  assign o[33191] = i[64];
  assign o[33192] = i[64];
  assign o[33193] = i[64];
  assign o[33194] = i[64];
  assign o[33195] = i[64];
  assign o[33196] = i[64];
  assign o[33197] = i[64];
  assign o[33198] = i[64];
  assign o[33199] = i[64];
  assign o[33200] = i[64];
  assign o[33201] = i[64];
  assign o[33202] = i[64];
  assign o[33203] = i[64];
  assign o[33204] = i[64];
  assign o[33205] = i[64];
  assign o[33206] = i[64];
  assign o[33207] = i[64];
  assign o[33208] = i[64];
  assign o[33209] = i[64];
  assign o[33210] = i[64];
  assign o[33211] = i[64];
  assign o[33212] = i[64];
  assign o[33213] = i[64];
  assign o[33214] = i[64];
  assign o[33215] = i[64];
  assign o[33216] = i[64];
  assign o[33217] = i[64];
  assign o[33218] = i[64];
  assign o[33219] = i[64];
  assign o[33220] = i[64];
  assign o[33221] = i[64];
  assign o[33222] = i[64];
  assign o[33223] = i[64];
  assign o[33224] = i[64];
  assign o[33225] = i[64];
  assign o[33226] = i[64];
  assign o[33227] = i[64];
  assign o[33228] = i[64];
  assign o[33229] = i[64];
  assign o[33230] = i[64];
  assign o[33231] = i[64];
  assign o[33232] = i[64];
  assign o[33233] = i[64];
  assign o[33234] = i[64];
  assign o[33235] = i[64];
  assign o[33236] = i[64];
  assign o[33237] = i[64];
  assign o[33238] = i[64];
  assign o[33239] = i[64];
  assign o[33240] = i[64];
  assign o[33241] = i[64];
  assign o[33242] = i[64];
  assign o[33243] = i[64];
  assign o[33244] = i[64];
  assign o[33245] = i[64];
  assign o[33246] = i[64];
  assign o[33247] = i[64];
  assign o[33248] = i[64];
  assign o[33249] = i[64];
  assign o[33250] = i[64];
  assign o[33251] = i[64];
  assign o[33252] = i[64];
  assign o[33253] = i[64];
  assign o[33254] = i[64];
  assign o[33255] = i[64];
  assign o[33256] = i[64];
  assign o[33257] = i[64];
  assign o[33258] = i[64];
  assign o[33259] = i[64];
  assign o[33260] = i[64];
  assign o[33261] = i[64];
  assign o[33262] = i[64];
  assign o[33263] = i[64];
  assign o[33264] = i[64];
  assign o[33265] = i[64];
  assign o[33266] = i[64];
  assign o[33267] = i[64];
  assign o[33268] = i[64];
  assign o[33269] = i[64];
  assign o[33270] = i[64];
  assign o[33271] = i[64];
  assign o[33272] = i[64];
  assign o[33273] = i[64];
  assign o[33274] = i[64];
  assign o[33275] = i[64];
  assign o[33276] = i[64];
  assign o[33277] = i[64];
  assign o[33278] = i[64];
  assign o[33279] = i[64];
  assign o[32256] = i[63];
  assign o[32257] = i[63];
  assign o[32258] = i[63];
  assign o[32259] = i[63];
  assign o[32260] = i[63];
  assign o[32261] = i[63];
  assign o[32262] = i[63];
  assign o[32263] = i[63];
  assign o[32264] = i[63];
  assign o[32265] = i[63];
  assign o[32266] = i[63];
  assign o[32267] = i[63];
  assign o[32268] = i[63];
  assign o[32269] = i[63];
  assign o[32270] = i[63];
  assign o[32271] = i[63];
  assign o[32272] = i[63];
  assign o[32273] = i[63];
  assign o[32274] = i[63];
  assign o[32275] = i[63];
  assign o[32276] = i[63];
  assign o[32277] = i[63];
  assign o[32278] = i[63];
  assign o[32279] = i[63];
  assign o[32280] = i[63];
  assign o[32281] = i[63];
  assign o[32282] = i[63];
  assign o[32283] = i[63];
  assign o[32284] = i[63];
  assign o[32285] = i[63];
  assign o[32286] = i[63];
  assign o[32287] = i[63];
  assign o[32288] = i[63];
  assign o[32289] = i[63];
  assign o[32290] = i[63];
  assign o[32291] = i[63];
  assign o[32292] = i[63];
  assign o[32293] = i[63];
  assign o[32294] = i[63];
  assign o[32295] = i[63];
  assign o[32296] = i[63];
  assign o[32297] = i[63];
  assign o[32298] = i[63];
  assign o[32299] = i[63];
  assign o[32300] = i[63];
  assign o[32301] = i[63];
  assign o[32302] = i[63];
  assign o[32303] = i[63];
  assign o[32304] = i[63];
  assign o[32305] = i[63];
  assign o[32306] = i[63];
  assign o[32307] = i[63];
  assign o[32308] = i[63];
  assign o[32309] = i[63];
  assign o[32310] = i[63];
  assign o[32311] = i[63];
  assign o[32312] = i[63];
  assign o[32313] = i[63];
  assign o[32314] = i[63];
  assign o[32315] = i[63];
  assign o[32316] = i[63];
  assign o[32317] = i[63];
  assign o[32318] = i[63];
  assign o[32319] = i[63];
  assign o[32320] = i[63];
  assign o[32321] = i[63];
  assign o[32322] = i[63];
  assign o[32323] = i[63];
  assign o[32324] = i[63];
  assign o[32325] = i[63];
  assign o[32326] = i[63];
  assign o[32327] = i[63];
  assign o[32328] = i[63];
  assign o[32329] = i[63];
  assign o[32330] = i[63];
  assign o[32331] = i[63];
  assign o[32332] = i[63];
  assign o[32333] = i[63];
  assign o[32334] = i[63];
  assign o[32335] = i[63];
  assign o[32336] = i[63];
  assign o[32337] = i[63];
  assign o[32338] = i[63];
  assign o[32339] = i[63];
  assign o[32340] = i[63];
  assign o[32341] = i[63];
  assign o[32342] = i[63];
  assign o[32343] = i[63];
  assign o[32344] = i[63];
  assign o[32345] = i[63];
  assign o[32346] = i[63];
  assign o[32347] = i[63];
  assign o[32348] = i[63];
  assign o[32349] = i[63];
  assign o[32350] = i[63];
  assign o[32351] = i[63];
  assign o[32352] = i[63];
  assign o[32353] = i[63];
  assign o[32354] = i[63];
  assign o[32355] = i[63];
  assign o[32356] = i[63];
  assign o[32357] = i[63];
  assign o[32358] = i[63];
  assign o[32359] = i[63];
  assign o[32360] = i[63];
  assign o[32361] = i[63];
  assign o[32362] = i[63];
  assign o[32363] = i[63];
  assign o[32364] = i[63];
  assign o[32365] = i[63];
  assign o[32366] = i[63];
  assign o[32367] = i[63];
  assign o[32368] = i[63];
  assign o[32369] = i[63];
  assign o[32370] = i[63];
  assign o[32371] = i[63];
  assign o[32372] = i[63];
  assign o[32373] = i[63];
  assign o[32374] = i[63];
  assign o[32375] = i[63];
  assign o[32376] = i[63];
  assign o[32377] = i[63];
  assign o[32378] = i[63];
  assign o[32379] = i[63];
  assign o[32380] = i[63];
  assign o[32381] = i[63];
  assign o[32382] = i[63];
  assign o[32383] = i[63];
  assign o[32384] = i[63];
  assign o[32385] = i[63];
  assign o[32386] = i[63];
  assign o[32387] = i[63];
  assign o[32388] = i[63];
  assign o[32389] = i[63];
  assign o[32390] = i[63];
  assign o[32391] = i[63];
  assign o[32392] = i[63];
  assign o[32393] = i[63];
  assign o[32394] = i[63];
  assign o[32395] = i[63];
  assign o[32396] = i[63];
  assign o[32397] = i[63];
  assign o[32398] = i[63];
  assign o[32399] = i[63];
  assign o[32400] = i[63];
  assign o[32401] = i[63];
  assign o[32402] = i[63];
  assign o[32403] = i[63];
  assign o[32404] = i[63];
  assign o[32405] = i[63];
  assign o[32406] = i[63];
  assign o[32407] = i[63];
  assign o[32408] = i[63];
  assign o[32409] = i[63];
  assign o[32410] = i[63];
  assign o[32411] = i[63];
  assign o[32412] = i[63];
  assign o[32413] = i[63];
  assign o[32414] = i[63];
  assign o[32415] = i[63];
  assign o[32416] = i[63];
  assign o[32417] = i[63];
  assign o[32418] = i[63];
  assign o[32419] = i[63];
  assign o[32420] = i[63];
  assign o[32421] = i[63];
  assign o[32422] = i[63];
  assign o[32423] = i[63];
  assign o[32424] = i[63];
  assign o[32425] = i[63];
  assign o[32426] = i[63];
  assign o[32427] = i[63];
  assign o[32428] = i[63];
  assign o[32429] = i[63];
  assign o[32430] = i[63];
  assign o[32431] = i[63];
  assign o[32432] = i[63];
  assign o[32433] = i[63];
  assign o[32434] = i[63];
  assign o[32435] = i[63];
  assign o[32436] = i[63];
  assign o[32437] = i[63];
  assign o[32438] = i[63];
  assign o[32439] = i[63];
  assign o[32440] = i[63];
  assign o[32441] = i[63];
  assign o[32442] = i[63];
  assign o[32443] = i[63];
  assign o[32444] = i[63];
  assign o[32445] = i[63];
  assign o[32446] = i[63];
  assign o[32447] = i[63];
  assign o[32448] = i[63];
  assign o[32449] = i[63];
  assign o[32450] = i[63];
  assign o[32451] = i[63];
  assign o[32452] = i[63];
  assign o[32453] = i[63];
  assign o[32454] = i[63];
  assign o[32455] = i[63];
  assign o[32456] = i[63];
  assign o[32457] = i[63];
  assign o[32458] = i[63];
  assign o[32459] = i[63];
  assign o[32460] = i[63];
  assign o[32461] = i[63];
  assign o[32462] = i[63];
  assign o[32463] = i[63];
  assign o[32464] = i[63];
  assign o[32465] = i[63];
  assign o[32466] = i[63];
  assign o[32467] = i[63];
  assign o[32468] = i[63];
  assign o[32469] = i[63];
  assign o[32470] = i[63];
  assign o[32471] = i[63];
  assign o[32472] = i[63];
  assign o[32473] = i[63];
  assign o[32474] = i[63];
  assign o[32475] = i[63];
  assign o[32476] = i[63];
  assign o[32477] = i[63];
  assign o[32478] = i[63];
  assign o[32479] = i[63];
  assign o[32480] = i[63];
  assign o[32481] = i[63];
  assign o[32482] = i[63];
  assign o[32483] = i[63];
  assign o[32484] = i[63];
  assign o[32485] = i[63];
  assign o[32486] = i[63];
  assign o[32487] = i[63];
  assign o[32488] = i[63];
  assign o[32489] = i[63];
  assign o[32490] = i[63];
  assign o[32491] = i[63];
  assign o[32492] = i[63];
  assign o[32493] = i[63];
  assign o[32494] = i[63];
  assign o[32495] = i[63];
  assign o[32496] = i[63];
  assign o[32497] = i[63];
  assign o[32498] = i[63];
  assign o[32499] = i[63];
  assign o[32500] = i[63];
  assign o[32501] = i[63];
  assign o[32502] = i[63];
  assign o[32503] = i[63];
  assign o[32504] = i[63];
  assign o[32505] = i[63];
  assign o[32506] = i[63];
  assign o[32507] = i[63];
  assign o[32508] = i[63];
  assign o[32509] = i[63];
  assign o[32510] = i[63];
  assign o[32511] = i[63];
  assign o[32512] = i[63];
  assign o[32513] = i[63];
  assign o[32514] = i[63];
  assign o[32515] = i[63];
  assign o[32516] = i[63];
  assign o[32517] = i[63];
  assign o[32518] = i[63];
  assign o[32519] = i[63];
  assign o[32520] = i[63];
  assign o[32521] = i[63];
  assign o[32522] = i[63];
  assign o[32523] = i[63];
  assign o[32524] = i[63];
  assign o[32525] = i[63];
  assign o[32526] = i[63];
  assign o[32527] = i[63];
  assign o[32528] = i[63];
  assign o[32529] = i[63];
  assign o[32530] = i[63];
  assign o[32531] = i[63];
  assign o[32532] = i[63];
  assign o[32533] = i[63];
  assign o[32534] = i[63];
  assign o[32535] = i[63];
  assign o[32536] = i[63];
  assign o[32537] = i[63];
  assign o[32538] = i[63];
  assign o[32539] = i[63];
  assign o[32540] = i[63];
  assign o[32541] = i[63];
  assign o[32542] = i[63];
  assign o[32543] = i[63];
  assign o[32544] = i[63];
  assign o[32545] = i[63];
  assign o[32546] = i[63];
  assign o[32547] = i[63];
  assign o[32548] = i[63];
  assign o[32549] = i[63];
  assign o[32550] = i[63];
  assign o[32551] = i[63];
  assign o[32552] = i[63];
  assign o[32553] = i[63];
  assign o[32554] = i[63];
  assign o[32555] = i[63];
  assign o[32556] = i[63];
  assign o[32557] = i[63];
  assign o[32558] = i[63];
  assign o[32559] = i[63];
  assign o[32560] = i[63];
  assign o[32561] = i[63];
  assign o[32562] = i[63];
  assign o[32563] = i[63];
  assign o[32564] = i[63];
  assign o[32565] = i[63];
  assign o[32566] = i[63];
  assign o[32567] = i[63];
  assign o[32568] = i[63];
  assign o[32569] = i[63];
  assign o[32570] = i[63];
  assign o[32571] = i[63];
  assign o[32572] = i[63];
  assign o[32573] = i[63];
  assign o[32574] = i[63];
  assign o[32575] = i[63];
  assign o[32576] = i[63];
  assign o[32577] = i[63];
  assign o[32578] = i[63];
  assign o[32579] = i[63];
  assign o[32580] = i[63];
  assign o[32581] = i[63];
  assign o[32582] = i[63];
  assign o[32583] = i[63];
  assign o[32584] = i[63];
  assign o[32585] = i[63];
  assign o[32586] = i[63];
  assign o[32587] = i[63];
  assign o[32588] = i[63];
  assign o[32589] = i[63];
  assign o[32590] = i[63];
  assign o[32591] = i[63];
  assign o[32592] = i[63];
  assign o[32593] = i[63];
  assign o[32594] = i[63];
  assign o[32595] = i[63];
  assign o[32596] = i[63];
  assign o[32597] = i[63];
  assign o[32598] = i[63];
  assign o[32599] = i[63];
  assign o[32600] = i[63];
  assign o[32601] = i[63];
  assign o[32602] = i[63];
  assign o[32603] = i[63];
  assign o[32604] = i[63];
  assign o[32605] = i[63];
  assign o[32606] = i[63];
  assign o[32607] = i[63];
  assign o[32608] = i[63];
  assign o[32609] = i[63];
  assign o[32610] = i[63];
  assign o[32611] = i[63];
  assign o[32612] = i[63];
  assign o[32613] = i[63];
  assign o[32614] = i[63];
  assign o[32615] = i[63];
  assign o[32616] = i[63];
  assign o[32617] = i[63];
  assign o[32618] = i[63];
  assign o[32619] = i[63];
  assign o[32620] = i[63];
  assign o[32621] = i[63];
  assign o[32622] = i[63];
  assign o[32623] = i[63];
  assign o[32624] = i[63];
  assign o[32625] = i[63];
  assign o[32626] = i[63];
  assign o[32627] = i[63];
  assign o[32628] = i[63];
  assign o[32629] = i[63];
  assign o[32630] = i[63];
  assign o[32631] = i[63];
  assign o[32632] = i[63];
  assign o[32633] = i[63];
  assign o[32634] = i[63];
  assign o[32635] = i[63];
  assign o[32636] = i[63];
  assign o[32637] = i[63];
  assign o[32638] = i[63];
  assign o[32639] = i[63];
  assign o[32640] = i[63];
  assign o[32641] = i[63];
  assign o[32642] = i[63];
  assign o[32643] = i[63];
  assign o[32644] = i[63];
  assign o[32645] = i[63];
  assign o[32646] = i[63];
  assign o[32647] = i[63];
  assign o[32648] = i[63];
  assign o[32649] = i[63];
  assign o[32650] = i[63];
  assign o[32651] = i[63];
  assign o[32652] = i[63];
  assign o[32653] = i[63];
  assign o[32654] = i[63];
  assign o[32655] = i[63];
  assign o[32656] = i[63];
  assign o[32657] = i[63];
  assign o[32658] = i[63];
  assign o[32659] = i[63];
  assign o[32660] = i[63];
  assign o[32661] = i[63];
  assign o[32662] = i[63];
  assign o[32663] = i[63];
  assign o[32664] = i[63];
  assign o[32665] = i[63];
  assign o[32666] = i[63];
  assign o[32667] = i[63];
  assign o[32668] = i[63];
  assign o[32669] = i[63];
  assign o[32670] = i[63];
  assign o[32671] = i[63];
  assign o[32672] = i[63];
  assign o[32673] = i[63];
  assign o[32674] = i[63];
  assign o[32675] = i[63];
  assign o[32676] = i[63];
  assign o[32677] = i[63];
  assign o[32678] = i[63];
  assign o[32679] = i[63];
  assign o[32680] = i[63];
  assign o[32681] = i[63];
  assign o[32682] = i[63];
  assign o[32683] = i[63];
  assign o[32684] = i[63];
  assign o[32685] = i[63];
  assign o[32686] = i[63];
  assign o[32687] = i[63];
  assign o[32688] = i[63];
  assign o[32689] = i[63];
  assign o[32690] = i[63];
  assign o[32691] = i[63];
  assign o[32692] = i[63];
  assign o[32693] = i[63];
  assign o[32694] = i[63];
  assign o[32695] = i[63];
  assign o[32696] = i[63];
  assign o[32697] = i[63];
  assign o[32698] = i[63];
  assign o[32699] = i[63];
  assign o[32700] = i[63];
  assign o[32701] = i[63];
  assign o[32702] = i[63];
  assign o[32703] = i[63];
  assign o[32704] = i[63];
  assign o[32705] = i[63];
  assign o[32706] = i[63];
  assign o[32707] = i[63];
  assign o[32708] = i[63];
  assign o[32709] = i[63];
  assign o[32710] = i[63];
  assign o[32711] = i[63];
  assign o[32712] = i[63];
  assign o[32713] = i[63];
  assign o[32714] = i[63];
  assign o[32715] = i[63];
  assign o[32716] = i[63];
  assign o[32717] = i[63];
  assign o[32718] = i[63];
  assign o[32719] = i[63];
  assign o[32720] = i[63];
  assign o[32721] = i[63];
  assign o[32722] = i[63];
  assign o[32723] = i[63];
  assign o[32724] = i[63];
  assign o[32725] = i[63];
  assign o[32726] = i[63];
  assign o[32727] = i[63];
  assign o[32728] = i[63];
  assign o[32729] = i[63];
  assign o[32730] = i[63];
  assign o[32731] = i[63];
  assign o[32732] = i[63];
  assign o[32733] = i[63];
  assign o[32734] = i[63];
  assign o[32735] = i[63];
  assign o[32736] = i[63];
  assign o[32737] = i[63];
  assign o[32738] = i[63];
  assign o[32739] = i[63];
  assign o[32740] = i[63];
  assign o[32741] = i[63];
  assign o[32742] = i[63];
  assign o[32743] = i[63];
  assign o[32744] = i[63];
  assign o[32745] = i[63];
  assign o[32746] = i[63];
  assign o[32747] = i[63];
  assign o[32748] = i[63];
  assign o[32749] = i[63];
  assign o[32750] = i[63];
  assign o[32751] = i[63];
  assign o[32752] = i[63];
  assign o[32753] = i[63];
  assign o[32754] = i[63];
  assign o[32755] = i[63];
  assign o[32756] = i[63];
  assign o[32757] = i[63];
  assign o[32758] = i[63];
  assign o[32759] = i[63];
  assign o[32760] = i[63];
  assign o[32761] = i[63];
  assign o[32762] = i[63];
  assign o[32763] = i[63];
  assign o[32764] = i[63];
  assign o[32765] = i[63];
  assign o[32766] = i[63];
  assign o[32767] = i[63];
  assign o[31744] = i[62];
  assign o[31745] = i[62];
  assign o[31746] = i[62];
  assign o[31747] = i[62];
  assign o[31748] = i[62];
  assign o[31749] = i[62];
  assign o[31750] = i[62];
  assign o[31751] = i[62];
  assign o[31752] = i[62];
  assign o[31753] = i[62];
  assign o[31754] = i[62];
  assign o[31755] = i[62];
  assign o[31756] = i[62];
  assign o[31757] = i[62];
  assign o[31758] = i[62];
  assign o[31759] = i[62];
  assign o[31760] = i[62];
  assign o[31761] = i[62];
  assign o[31762] = i[62];
  assign o[31763] = i[62];
  assign o[31764] = i[62];
  assign o[31765] = i[62];
  assign o[31766] = i[62];
  assign o[31767] = i[62];
  assign o[31768] = i[62];
  assign o[31769] = i[62];
  assign o[31770] = i[62];
  assign o[31771] = i[62];
  assign o[31772] = i[62];
  assign o[31773] = i[62];
  assign o[31774] = i[62];
  assign o[31775] = i[62];
  assign o[31776] = i[62];
  assign o[31777] = i[62];
  assign o[31778] = i[62];
  assign o[31779] = i[62];
  assign o[31780] = i[62];
  assign o[31781] = i[62];
  assign o[31782] = i[62];
  assign o[31783] = i[62];
  assign o[31784] = i[62];
  assign o[31785] = i[62];
  assign o[31786] = i[62];
  assign o[31787] = i[62];
  assign o[31788] = i[62];
  assign o[31789] = i[62];
  assign o[31790] = i[62];
  assign o[31791] = i[62];
  assign o[31792] = i[62];
  assign o[31793] = i[62];
  assign o[31794] = i[62];
  assign o[31795] = i[62];
  assign o[31796] = i[62];
  assign o[31797] = i[62];
  assign o[31798] = i[62];
  assign o[31799] = i[62];
  assign o[31800] = i[62];
  assign o[31801] = i[62];
  assign o[31802] = i[62];
  assign o[31803] = i[62];
  assign o[31804] = i[62];
  assign o[31805] = i[62];
  assign o[31806] = i[62];
  assign o[31807] = i[62];
  assign o[31808] = i[62];
  assign o[31809] = i[62];
  assign o[31810] = i[62];
  assign o[31811] = i[62];
  assign o[31812] = i[62];
  assign o[31813] = i[62];
  assign o[31814] = i[62];
  assign o[31815] = i[62];
  assign o[31816] = i[62];
  assign o[31817] = i[62];
  assign o[31818] = i[62];
  assign o[31819] = i[62];
  assign o[31820] = i[62];
  assign o[31821] = i[62];
  assign o[31822] = i[62];
  assign o[31823] = i[62];
  assign o[31824] = i[62];
  assign o[31825] = i[62];
  assign o[31826] = i[62];
  assign o[31827] = i[62];
  assign o[31828] = i[62];
  assign o[31829] = i[62];
  assign o[31830] = i[62];
  assign o[31831] = i[62];
  assign o[31832] = i[62];
  assign o[31833] = i[62];
  assign o[31834] = i[62];
  assign o[31835] = i[62];
  assign o[31836] = i[62];
  assign o[31837] = i[62];
  assign o[31838] = i[62];
  assign o[31839] = i[62];
  assign o[31840] = i[62];
  assign o[31841] = i[62];
  assign o[31842] = i[62];
  assign o[31843] = i[62];
  assign o[31844] = i[62];
  assign o[31845] = i[62];
  assign o[31846] = i[62];
  assign o[31847] = i[62];
  assign o[31848] = i[62];
  assign o[31849] = i[62];
  assign o[31850] = i[62];
  assign o[31851] = i[62];
  assign o[31852] = i[62];
  assign o[31853] = i[62];
  assign o[31854] = i[62];
  assign o[31855] = i[62];
  assign o[31856] = i[62];
  assign o[31857] = i[62];
  assign o[31858] = i[62];
  assign o[31859] = i[62];
  assign o[31860] = i[62];
  assign o[31861] = i[62];
  assign o[31862] = i[62];
  assign o[31863] = i[62];
  assign o[31864] = i[62];
  assign o[31865] = i[62];
  assign o[31866] = i[62];
  assign o[31867] = i[62];
  assign o[31868] = i[62];
  assign o[31869] = i[62];
  assign o[31870] = i[62];
  assign o[31871] = i[62];
  assign o[31872] = i[62];
  assign o[31873] = i[62];
  assign o[31874] = i[62];
  assign o[31875] = i[62];
  assign o[31876] = i[62];
  assign o[31877] = i[62];
  assign o[31878] = i[62];
  assign o[31879] = i[62];
  assign o[31880] = i[62];
  assign o[31881] = i[62];
  assign o[31882] = i[62];
  assign o[31883] = i[62];
  assign o[31884] = i[62];
  assign o[31885] = i[62];
  assign o[31886] = i[62];
  assign o[31887] = i[62];
  assign o[31888] = i[62];
  assign o[31889] = i[62];
  assign o[31890] = i[62];
  assign o[31891] = i[62];
  assign o[31892] = i[62];
  assign o[31893] = i[62];
  assign o[31894] = i[62];
  assign o[31895] = i[62];
  assign o[31896] = i[62];
  assign o[31897] = i[62];
  assign o[31898] = i[62];
  assign o[31899] = i[62];
  assign o[31900] = i[62];
  assign o[31901] = i[62];
  assign o[31902] = i[62];
  assign o[31903] = i[62];
  assign o[31904] = i[62];
  assign o[31905] = i[62];
  assign o[31906] = i[62];
  assign o[31907] = i[62];
  assign o[31908] = i[62];
  assign o[31909] = i[62];
  assign o[31910] = i[62];
  assign o[31911] = i[62];
  assign o[31912] = i[62];
  assign o[31913] = i[62];
  assign o[31914] = i[62];
  assign o[31915] = i[62];
  assign o[31916] = i[62];
  assign o[31917] = i[62];
  assign o[31918] = i[62];
  assign o[31919] = i[62];
  assign o[31920] = i[62];
  assign o[31921] = i[62];
  assign o[31922] = i[62];
  assign o[31923] = i[62];
  assign o[31924] = i[62];
  assign o[31925] = i[62];
  assign o[31926] = i[62];
  assign o[31927] = i[62];
  assign o[31928] = i[62];
  assign o[31929] = i[62];
  assign o[31930] = i[62];
  assign o[31931] = i[62];
  assign o[31932] = i[62];
  assign o[31933] = i[62];
  assign o[31934] = i[62];
  assign o[31935] = i[62];
  assign o[31936] = i[62];
  assign o[31937] = i[62];
  assign o[31938] = i[62];
  assign o[31939] = i[62];
  assign o[31940] = i[62];
  assign o[31941] = i[62];
  assign o[31942] = i[62];
  assign o[31943] = i[62];
  assign o[31944] = i[62];
  assign o[31945] = i[62];
  assign o[31946] = i[62];
  assign o[31947] = i[62];
  assign o[31948] = i[62];
  assign o[31949] = i[62];
  assign o[31950] = i[62];
  assign o[31951] = i[62];
  assign o[31952] = i[62];
  assign o[31953] = i[62];
  assign o[31954] = i[62];
  assign o[31955] = i[62];
  assign o[31956] = i[62];
  assign o[31957] = i[62];
  assign o[31958] = i[62];
  assign o[31959] = i[62];
  assign o[31960] = i[62];
  assign o[31961] = i[62];
  assign o[31962] = i[62];
  assign o[31963] = i[62];
  assign o[31964] = i[62];
  assign o[31965] = i[62];
  assign o[31966] = i[62];
  assign o[31967] = i[62];
  assign o[31968] = i[62];
  assign o[31969] = i[62];
  assign o[31970] = i[62];
  assign o[31971] = i[62];
  assign o[31972] = i[62];
  assign o[31973] = i[62];
  assign o[31974] = i[62];
  assign o[31975] = i[62];
  assign o[31976] = i[62];
  assign o[31977] = i[62];
  assign o[31978] = i[62];
  assign o[31979] = i[62];
  assign o[31980] = i[62];
  assign o[31981] = i[62];
  assign o[31982] = i[62];
  assign o[31983] = i[62];
  assign o[31984] = i[62];
  assign o[31985] = i[62];
  assign o[31986] = i[62];
  assign o[31987] = i[62];
  assign o[31988] = i[62];
  assign o[31989] = i[62];
  assign o[31990] = i[62];
  assign o[31991] = i[62];
  assign o[31992] = i[62];
  assign o[31993] = i[62];
  assign o[31994] = i[62];
  assign o[31995] = i[62];
  assign o[31996] = i[62];
  assign o[31997] = i[62];
  assign o[31998] = i[62];
  assign o[31999] = i[62];
  assign o[32000] = i[62];
  assign o[32001] = i[62];
  assign o[32002] = i[62];
  assign o[32003] = i[62];
  assign o[32004] = i[62];
  assign o[32005] = i[62];
  assign o[32006] = i[62];
  assign o[32007] = i[62];
  assign o[32008] = i[62];
  assign o[32009] = i[62];
  assign o[32010] = i[62];
  assign o[32011] = i[62];
  assign o[32012] = i[62];
  assign o[32013] = i[62];
  assign o[32014] = i[62];
  assign o[32015] = i[62];
  assign o[32016] = i[62];
  assign o[32017] = i[62];
  assign o[32018] = i[62];
  assign o[32019] = i[62];
  assign o[32020] = i[62];
  assign o[32021] = i[62];
  assign o[32022] = i[62];
  assign o[32023] = i[62];
  assign o[32024] = i[62];
  assign o[32025] = i[62];
  assign o[32026] = i[62];
  assign o[32027] = i[62];
  assign o[32028] = i[62];
  assign o[32029] = i[62];
  assign o[32030] = i[62];
  assign o[32031] = i[62];
  assign o[32032] = i[62];
  assign o[32033] = i[62];
  assign o[32034] = i[62];
  assign o[32035] = i[62];
  assign o[32036] = i[62];
  assign o[32037] = i[62];
  assign o[32038] = i[62];
  assign o[32039] = i[62];
  assign o[32040] = i[62];
  assign o[32041] = i[62];
  assign o[32042] = i[62];
  assign o[32043] = i[62];
  assign o[32044] = i[62];
  assign o[32045] = i[62];
  assign o[32046] = i[62];
  assign o[32047] = i[62];
  assign o[32048] = i[62];
  assign o[32049] = i[62];
  assign o[32050] = i[62];
  assign o[32051] = i[62];
  assign o[32052] = i[62];
  assign o[32053] = i[62];
  assign o[32054] = i[62];
  assign o[32055] = i[62];
  assign o[32056] = i[62];
  assign o[32057] = i[62];
  assign o[32058] = i[62];
  assign o[32059] = i[62];
  assign o[32060] = i[62];
  assign o[32061] = i[62];
  assign o[32062] = i[62];
  assign o[32063] = i[62];
  assign o[32064] = i[62];
  assign o[32065] = i[62];
  assign o[32066] = i[62];
  assign o[32067] = i[62];
  assign o[32068] = i[62];
  assign o[32069] = i[62];
  assign o[32070] = i[62];
  assign o[32071] = i[62];
  assign o[32072] = i[62];
  assign o[32073] = i[62];
  assign o[32074] = i[62];
  assign o[32075] = i[62];
  assign o[32076] = i[62];
  assign o[32077] = i[62];
  assign o[32078] = i[62];
  assign o[32079] = i[62];
  assign o[32080] = i[62];
  assign o[32081] = i[62];
  assign o[32082] = i[62];
  assign o[32083] = i[62];
  assign o[32084] = i[62];
  assign o[32085] = i[62];
  assign o[32086] = i[62];
  assign o[32087] = i[62];
  assign o[32088] = i[62];
  assign o[32089] = i[62];
  assign o[32090] = i[62];
  assign o[32091] = i[62];
  assign o[32092] = i[62];
  assign o[32093] = i[62];
  assign o[32094] = i[62];
  assign o[32095] = i[62];
  assign o[32096] = i[62];
  assign o[32097] = i[62];
  assign o[32098] = i[62];
  assign o[32099] = i[62];
  assign o[32100] = i[62];
  assign o[32101] = i[62];
  assign o[32102] = i[62];
  assign o[32103] = i[62];
  assign o[32104] = i[62];
  assign o[32105] = i[62];
  assign o[32106] = i[62];
  assign o[32107] = i[62];
  assign o[32108] = i[62];
  assign o[32109] = i[62];
  assign o[32110] = i[62];
  assign o[32111] = i[62];
  assign o[32112] = i[62];
  assign o[32113] = i[62];
  assign o[32114] = i[62];
  assign o[32115] = i[62];
  assign o[32116] = i[62];
  assign o[32117] = i[62];
  assign o[32118] = i[62];
  assign o[32119] = i[62];
  assign o[32120] = i[62];
  assign o[32121] = i[62];
  assign o[32122] = i[62];
  assign o[32123] = i[62];
  assign o[32124] = i[62];
  assign o[32125] = i[62];
  assign o[32126] = i[62];
  assign o[32127] = i[62];
  assign o[32128] = i[62];
  assign o[32129] = i[62];
  assign o[32130] = i[62];
  assign o[32131] = i[62];
  assign o[32132] = i[62];
  assign o[32133] = i[62];
  assign o[32134] = i[62];
  assign o[32135] = i[62];
  assign o[32136] = i[62];
  assign o[32137] = i[62];
  assign o[32138] = i[62];
  assign o[32139] = i[62];
  assign o[32140] = i[62];
  assign o[32141] = i[62];
  assign o[32142] = i[62];
  assign o[32143] = i[62];
  assign o[32144] = i[62];
  assign o[32145] = i[62];
  assign o[32146] = i[62];
  assign o[32147] = i[62];
  assign o[32148] = i[62];
  assign o[32149] = i[62];
  assign o[32150] = i[62];
  assign o[32151] = i[62];
  assign o[32152] = i[62];
  assign o[32153] = i[62];
  assign o[32154] = i[62];
  assign o[32155] = i[62];
  assign o[32156] = i[62];
  assign o[32157] = i[62];
  assign o[32158] = i[62];
  assign o[32159] = i[62];
  assign o[32160] = i[62];
  assign o[32161] = i[62];
  assign o[32162] = i[62];
  assign o[32163] = i[62];
  assign o[32164] = i[62];
  assign o[32165] = i[62];
  assign o[32166] = i[62];
  assign o[32167] = i[62];
  assign o[32168] = i[62];
  assign o[32169] = i[62];
  assign o[32170] = i[62];
  assign o[32171] = i[62];
  assign o[32172] = i[62];
  assign o[32173] = i[62];
  assign o[32174] = i[62];
  assign o[32175] = i[62];
  assign o[32176] = i[62];
  assign o[32177] = i[62];
  assign o[32178] = i[62];
  assign o[32179] = i[62];
  assign o[32180] = i[62];
  assign o[32181] = i[62];
  assign o[32182] = i[62];
  assign o[32183] = i[62];
  assign o[32184] = i[62];
  assign o[32185] = i[62];
  assign o[32186] = i[62];
  assign o[32187] = i[62];
  assign o[32188] = i[62];
  assign o[32189] = i[62];
  assign o[32190] = i[62];
  assign o[32191] = i[62];
  assign o[32192] = i[62];
  assign o[32193] = i[62];
  assign o[32194] = i[62];
  assign o[32195] = i[62];
  assign o[32196] = i[62];
  assign o[32197] = i[62];
  assign o[32198] = i[62];
  assign o[32199] = i[62];
  assign o[32200] = i[62];
  assign o[32201] = i[62];
  assign o[32202] = i[62];
  assign o[32203] = i[62];
  assign o[32204] = i[62];
  assign o[32205] = i[62];
  assign o[32206] = i[62];
  assign o[32207] = i[62];
  assign o[32208] = i[62];
  assign o[32209] = i[62];
  assign o[32210] = i[62];
  assign o[32211] = i[62];
  assign o[32212] = i[62];
  assign o[32213] = i[62];
  assign o[32214] = i[62];
  assign o[32215] = i[62];
  assign o[32216] = i[62];
  assign o[32217] = i[62];
  assign o[32218] = i[62];
  assign o[32219] = i[62];
  assign o[32220] = i[62];
  assign o[32221] = i[62];
  assign o[32222] = i[62];
  assign o[32223] = i[62];
  assign o[32224] = i[62];
  assign o[32225] = i[62];
  assign o[32226] = i[62];
  assign o[32227] = i[62];
  assign o[32228] = i[62];
  assign o[32229] = i[62];
  assign o[32230] = i[62];
  assign o[32231] = i[62];
  assign o[32232] = i[62];
  assign o[32233] = i[62];
  assign o[32234] = i[62];
  assign o[32235] = i[62];
  assign o[32236] = i[62];
  assign o[32237] = i[62];
  assign o[32238] = i[62];
  assign o[32239] = i[62];
  assign o[32240] = i[62];
  assign o[32241] = i[62];
  assign o[32242] = i[62];
  assign o[32243] = i[62];
  assign o[32244] = i[62];
  assign o[32245] = i[62];
  assign o[32246] = i[62];
  assign o[32247] = i[62];
  assign o[32248] = i[62];
  assign o[32249] = i[62];
  assign o[32250] = i[62];
  assign o[32251] = i[62];
  assign o[32252] = i[62];
  assign o[32253] = i[62];
  assign o[32254] = i[62];
  assign o[32255] = i[62];
  assign o[31232] = i[61];
  assign o[31233] = i[61];
  assign o[31234] = i[61];
  assign o[31235] = i[61];
  assign o[31236] = i[61];
  assign o[31237] = i[61];
  assign o[31238] = i[61];
  assign o[31239] = i[61];
  assign o[31240] = i[61];
  assign o[31241] = i[61];
  assign o[31242] = i[61];
  assign o[31243] = i[61];
  assign o[31244] = i[61];
  assign o[31245] = i[61];
  assign o[31246] = i[61];
  assign o[31247] = i[61];
  assign o[31248] = i[61];
  assign o[31249] = i[61];
  assign o[31250] = i[61];
  assign o[31251] = i[61];
  assign o[31252] = i[61];
  assign o[31253] = i[61];
  assign o[31254] = i[61];
  assign o[31255] = i[61];
  assign o[31256] = i[61];
  assign o[31257] = i[61];
  assign o[31258] = i[61];
  assign o[31259] = i[61];
  assign o[31260] = i[61];
  assign o[31261] = i[61];
  assign o[31262] = i[61];
  assign o[31263] = i[61];
  assign o[31264] = i[61];
  assign o[31265] = i[61];
  assign o[31266] = i[61];
  assign o[31267] = i[61];
  assign o[31268] = i[61];
  assign o[31269] = i[61];
  assign o[31270] = i[61];
  assign o[31271] = i[61];
  assign o[31272] = i[61];
  assign o[31273] = i[61];
  assign o[31274] = i[61];
  assign o[31275] = i[61];
  assign o[31276] = i[61];
  assign o[31277] = i[61];
  assign o[31278] = i[61];
  assign o[31279] = i[61];
  assign o[31280] = i[61];
  assign o[31281] = i[61];
  assign o[31282] = i[61];
  assign o[31283] = i[61];
  assign o[31284] = i[61];
  assign o[31285] = i[61];
  assign o[31286] = i[61];
  assign o[31287] = i[61];
  assign o[31288] = i[61];
  assign o[31289] = i[61];
  assign o[31290] = i[61];
  assign o[31291] = i[61];
  assign o[31292] = i[61];
  assign o[31293] = i[61];
  assign o[31294] = i[61];
  assign o[31295] = i[61];
  assign o[31296] = i[61];
  assign o[31297] = i[61];
  assign o[31298] = i[61];
  assign o[31299] = i[61];
  assign o[31300] = i[61];
  assign o[31301] = i[61];
  assign o[31302] = i[61];
  assign o[31303] = i[61];
  assign o[31304] = i[61];
  assign o[31305] = i[61];
  assign o[31306] = i[61];
  assign o[31307] = i[61];
  assign o[31308] = i[61];
  assign o[31309] = i[61];
  assign o[31310] = i[61];
  assign o[31311] = i[61];
  assign o[31312] = i[61];
  assign o[31313] = i[61];
  assign o[31314] = i[61];
  assign o[31315] = i[61];
  assign o[31316] = i[61];
  assign o[31317] = i[61];
  assign o[31318] = i[61];
  assign o[31319] = i[61];
  assign o[31320] = i[61];
  assign o[31321] = i[61];
  assign o[31322] = i[61];
  assign o[31323] = i[61];
  assign o[31324] = i[61];
  assign o[31325] = i[61];
  assign o[31326] = i[61];
  assign o[31327] = i[61];
  assign o[31328] = i[61];
  assign o[31329] = i[61];
  assign o[31330] = i[61];
  assign o[31331] = i[61];
  assign o[31332] = i[61];
  assign o[31333] = i[61];
  assign o[31334] = i[61];
  assign o[31335] = i[61];
  assign o[31336] = i[61];
  assign o[31337] = i[61];
  assign o[31338] = i[61];
  assign o[31339] = i[61];
  assign o[31340] = i[61];
  assign o[31341] = i[61];
  assign o[31342] = i[61];
  assign o[31343] = i[61];
  assign o[31344] = i[61];
  assign o[31345] = i[61];
  assign o[31346] = i[61];
  assign o[31347] = i[61];
  assign o[31348] = i[61];
  assign o[31349] = i[61];
  assign o[31350] = i[61];
  assign o[31351] = i[61];
  assign o[31352] = i[61];
  assign o[31353] = i[61];
  assign o[31354] = i[61];
  assign o[31355] = i[61];
  assign o[31356] = i[61];
  assign o[31357] = i[61];
  assign o[31358] = i[61];
  assign o[31359] = i[61];
  assign o[31360] = i[61];
  assign o[31361] = i[61];
  assign o[31362] = i[61];
  assign o[31363] = i[61];
  assign o[31364] = i[61];
  assign o[31365] = i[61];
  assign o[31366] = i[61];
  assign o[31367] = i[61];
  assign o[31368] = i[61];
  assign o[31369] = i[61];
  assign o[31370] = i[61];
  assign o[31371] = i[61];
  assign o[31372] = i[61];
  assign o[31373] = i[61];
  assign o[31374] = i[61];
  assign o[31375] = i[61];
  assign o[31376] = i[61];
  assign o[31377] = i[61];
  assign o[31378] = i[61];
  assign o[31379] = i[61];
  assign o[31380] = i[61];
  assign o[31381] = i[61];
  assign o[31382] = i[61];
  assign o[31383] = i[61];
  assign o[31384] = i[61];
  assign o[31385] = i[61];
  assign o[31386] = i[61];
  assign o[31387] = i[61];
  assign o[31388] = i[61];
  assign o[31389] = i[61];
  assign o[31390] = i[61];
  assign o[31391] = i[61];
  assign o[31392] = i[61];
  assign o[31393] = i[61];
  assign o[31394] = i[61];
  assign o[31395] = i[61];
  assign o[31396] = i[61];
  assign o[31397] = i[61];
  assign o[31398] = i[61];
  assign o[31399] = i[61];
  assign o[31400] = i[61];
  assign o[31401] = i[61];
  assign o[31402] = i[61];
  assign o[31403] = i[61];
  assign o[31404] = i[61];
  assign o[31405] = i[61];
  assign o[31406] = i[61];
  assign o[31407] = i[61];
  assign o[31408] = i[61];
  assign o[31409] = i[61];
  assign o[31410] = i[61];
  assign o[31411] = i[61];
  assign o[31412] = i[61];
  assign o[31413] = i[61];
  assign o[31414] = i[61];
  assign o[31415] = i[61];
  assign o[31416] = i[61];
  assign o[31417] = i[61];
  assign o[31418] = i[61];
  assign o[31419] = i[61];
  assign o[31420] = i[61];
  assign o[31421] = i[61];
  assign o[31422] = i[61];
  assign o[31423] = i[61];
  assign o[31424] = i[61];
  assign o[31425] = i[61];
  assign o[31426] = i[61];
  assign o[31427] = i[61];
  assign o[31428] = i[61];
  assign o[31429] = i[61];
  assign o[31430] = i[61];
  assign o[31431] = i[61];
  assign o[31432] = i[61];
  assign o[31433] = i[61];
  assign o[31434] = i[61];
  assign o[31435] = i[61];
  assign o[31436] = i[61];
  assign o[31437] = i[61];
  assign o[31438] = i[61];
  assign o[31439] = i[61];
  assign o[31440] = i[61];
  assign o[31441] = i[61];
  assign o[31442] = i[61];
  assign o[31443] = i[61];
  assign o[31444] = i[61];
  assign o[31445] = i[61];
  assign o[31446] = i[61];
  assign o[31447] = i[61];
  assign o[31448] = i[61];
  assign o[31449] = i[61];
  assign o[31450] = i[61];
  assign o[31451] = i[61];
  assign o[31452] = i[61];
  assign o[31453] = i[61];
  assign o[31454] = i[61];
  assign o[31455] = i[61];
  assign o[31456] = i[61];
  assign o[31457] = i[61];
  assign o[31458] = i[61];
  assign o[31459] = i[61];
  assign o[31460] = i[61];
  assign o[31461] = i[61];
  assign o[31462] = i[61];
  assign o[31463] = i[61];
  assign o[31464] = i[61];
  assign o[31465] = i[61];
  assign o[31466] = i[61];
  assign o[31467] = i[61];
  assign o[31468] = i[61];
  assign o[31469] = i[61];
  assign o[31470] = i[61];
  assign o[31471] = i[61];
  assign o[31472] = i[61];
  assign o[31473] = i[61];
  assign o[31474] = i[61];
  assign o[31475] = i[61];
  assign o[31476] = i[61];
  assign o[31477] = i[61];
  assign o[31478] = i[61];
  assign o[31479] = i[61];
  assign o[31480] = i[61];
  assign o[31481] = i[61];
  assign o[31482] = i[61];
  assign o[31483] = i[61];
  assign o[31484] = i[61];
  assign o[31485] = i[61];
  assign o[31486] = i[61];
  assign o[31487] = i[61];
  assign o[31488] = i[61];
  assign o[31489] = i[61];
  assign o[31490] = i[61];
  assign o[31491] = i[61];
  assign o[31492] = i[61];
  assign o[31493] = i[61];
  assign o[31494] = i[61];
  assign o[31495] = i[61];
  assign o[31496] = i[61];
  assign o[31497] = i[61];
  assign o[31498] = i[61];
  assign o[31499] = i[61];
  assign o[31500] = i[61];
  assign o[31501] = i[61];
  assign o[31502] = i[61];
  assign o[31503] = i[61];
  assign o[31504] = i[61];
  assign o[31505] = i[61];
  assign o[31506] = i[61];
  assign o[31507] = i[61];
  assign o[31508] = i[61];
  assign o[31509] = i[61];
  assign o[31510] = i[61];
  assign o[31511] = i[61];
  assign o[31512] = i[61];
  assign o[31513] = i[61];
  assign o[31514] = i[61];
  assign o[31515] = i[61];
  assign o[31516] = i[61];
  assign o[31517] = i[61];
  assign o[31518] = i[61];
  assign o[31519] = i[61];
  assign o[31520] = i[61];
  assign o[31521] = i[61];
  assign o[31522] = i[61];
  assign o[31523] = i[61];
  assign o[31524] = i[61];
  assign o[31525] = i[61];
  assign o[31526] = i[61];
  assign o[31527] = i[61];
  assign o[31528] = i[61];
  assign o[31529] = i[61];
  assign o[31530] = i[61];
  assign o[31531] = i[61];
  assign o[31532] = i[61];
  assign o[31533] = i[61];
  assign o[31534] = i[61];
  assign o[31535] = i[61];
  assign o[31536] = i[61];
  assign o[31537] = i[61];
  assign o[31538] = i[61];
  assign o[31539] = i[61];
  assign o[31540] = i[61];
  assign o[31541] = i[61];
  assign o[31542] = i[61];
  assign o[31543] = i[61];
  assign o[31544] = i[61];
  assign o[31545] = i[61];
  assign o[31546] = i[61];
  assign o[31547] = i[61];
  assign o[31548] = i[61];
  assign o[31549] = i[61];
  assign o[31550] = i[61];
  assign o[31551] = i[61];
  assign o[31552] = i[61];
  assign o[31553] = i[61];
  assign o[31554] = i[61];
  assign o[31555] = i[61];
  assign o[31556] = i[61];
  assign o[31557] = i[61];
  assign o[31558] = i[61];
  assign o[31559] = i[61];
  assign o[31560] = i[61];
  assign o[31561] = i[61];
  assign o[31562] = i[61];
  assign o[31563] = i[61];
  assign o[31564] = i[61];
  assign o[31565] = i[61];
  assign o[31566] = i[61];
  assign o[31567] = i[61];
  assign o[31568] = i[61];
  assign o[31569] = i[61];
  assign o[31570] = i[61];
  assign o[31571] = i[61];
  assign o[31572] = i[61];
  assign o[31573] = i[61];
  assign o[31574] = i[61];
  assign o[31575] = i[61];
  assign o[31576] = i[61];
  assign o[31577] = i[61];
  assign o[31578] = i[61];
  assign o[31579] = i[61];
  assign o[31580] = i[61];
  assign o[31581] = i[61];
  assign o[31582] = i[61];
  assign o[31583] = i[61];
  assign o[31584] = i[61];
  assign o[31585] = i[61];
  assign o[31586] = i[61];
  assign o[31587] = i[61];
  assign o[31588] = i[61];
  assign o[31589] = i[61];
  assign o[31590] = i[61];
  assign o[31591] = i[61];
  assign o[31592] = i[61];
  assign o[31593] = i[61];
  assign o[31594] = i[61];
  assign o[31595] = i[61];
  assign o[31596] = i[61];
  assign o[31597] = i[61];
  assign o[31598] = i[61];
  assign o[31599] = i[61];
  assign o[31600] = i[61];
  assign o[31601] = i[61];
  assign o[31602] = i[61];
  assign o[31603] = i[61];
  assign o[31604] = i[61];
  assign o[31605] = i[61];
  assign o[31606] = i[61];
  assign o[31607] = i[61];
  assign o[31608] = i[61];
  assign o[31609] = i[61];
  assign o[31610] = i[61];
  assign o[31611] = i[61];
  assign o[31612] = i[61];
  assign o[31613] = i[61];
  assign o[31614] = i[61];
  assign o[31615] = i[61];
  assign o[31616] = i[61];
  assign o[31617] = i[61];
  assign o[31618] = i[61];
  assign o[31619] = i[61];
  assign o[31620] = i[61];
  assign o[31621] = i[61];
  assign o[31622] = i[61];
  assign o[31623] = i[61];
  assign o[31624] = i[61];
  assign o[31625] = i[61];
  assign o[31626] = i[61];
  assign o[31627] = i[61];
  assign o[31628] = i[61];
  assign o[31629] = i[61];
  assign o[31630] = i[61];
  assign o[31631] = i[61];
  assign o[31632] = i[61];
  assign o[31633] = i[61];
  assign o[31634] = i[61];
  assign o[31635] = i[61];
  assign o[31636] = i[61];
  assign o[31637] = i[61];
  assign o[31638] = i[61];
  assign o[31639] = i[61];
  assign o[31640] = i[61];
  assign o[31641] = i[61];
  assign o[31642] = i[61];
  assign o[31643] = i[61];
  assign o[31644] = i[61];
  assign o[31645] = i[61];
  assign o[31646] = i[61];
  assign o[31647] = i[61];
  assign o[31648] = i[61];
  assign o[31649] = i[61];
  assign o[31650] = i[61];
  assign o[31651] = i[61];
  assign o[31652] = i[61];
  assign o[31653] = i[61];
  assign o[31654] = i[61];
  assign o[31655] = i[61];
  assign o[31656] = i[61];
  assign o[31657] = i[61];
  assign o[31658] = i[61];
  assign o[31659] = i[61];
  assign o[31660] = i[61];
  assign o[31661] = i[61];
  assign o[31662] = i[61];
  assign o[31663] = i[61];
  assign o[31664] = i[61];
  assign o[31665] = i[61];
  assign o[31666] = i[61];
  assign o[31667] = i[61];
  assign o[31668] = i[61];
  assign o[31669] = i[61];
  assign o[31670] = i[61];
  assign o[31671] = i[61];
  assign o[31672] = i[61];
  assign o[31673] = i[61];
  assign o[31674] = i[61];
  assign o[31675] = i[61];
  assign o[31676] = i[61];
  assign o[31677] = i[61];
  assign o[31678] = i[61];
  assign o[31679] = i[61];
  assign o[31680] = i[61];
  assign o[31681] = i[61];
  assign o[31682] = i[61];
  assign o[31683] = i[61];
  assign o[31684] = i[61];
  assign o[31685] = i[61];
  assign o[31686] = i[61];
  assign o[31687] = i[61];
  assign o[31688] = i[61];
  assign o[31689] = i[61];
  assign o[31690] = i[61];
  assign o[31691] = i[61];
  assign o[31692] = i[61];
  assign o[31693] = i[61];
  assign o[31694] = i[61];
  assign o[31695] = i[61];
  assign o[31696] = i[61];
  assign o[31697] = i[61];
  assign o[31698] = i[61];
  assign o[31699] = i[61];
  assign o[31700] = i[61];
  assign o[31701] = i[61];
  assign o[31702] = i[61];
  assign o[31703] = i[61];
  assign o[31704] = i[61];
  assign o[31705] = i[61];
  assign o[31706] = i[61];
  assign o[31707] = i[61];
  assign o[31708] = i[61];
  assign o[31709] = i[61];
  assign o[31710] = i[61];
  assign o[31711] = i[61];
  assign o[31712] = i[61];
  assign o[31713] = i[61];
  assign o[31714] = i[61];
  assign o[31715] = i[61];
  assign o[31716] = i[61];
  assign o[31717] = i[61];
  assign o[31718] = i[61];
  assign o[31719] = i[61];
  assign o[31720] = i[61];
  assign o[31721] = i[61];
  assign o[31722] = i[61];
  assign o[31723] = i[61];
  assign o[31724] = i[61];
  assign o[31725] = i[61];
  assign o[31726] = i[61];
  assign o[31727] = i[61];
  assign o[31728] = i[61];
  assign o[31729] = i[61];
  assign o[31730] = i[61];
  assign o[31731] = i[61];
  assign o[31732] = i[61];
  assign o[31733] = i[61];
  assign o[31734] = i[61];
  assign o[31735] = i[61];
  assign o[31736] = i[61];
  assign o[31737] = i[61];
  assign o[31738] = i[61];
  assign o[31739] = i[61];
  assign o[31740] = i[61];
  assign o[31741] = i[61];
  assign o[31742] = i[61];
  assign o[31743] = i[61];
  assign o[30720] = i[60];
  assign o[30721] = i[60];
  assign o[30722] = i[60];
  assign o[30723] = i[60];
  assign o[30724] = i[60];
  assign o[30725] = i[60];
  assign o[30726] = i[60];
  assign o[30727] = i[60];
  assign o[30728] = i[60];
  assign o[30729] = i[60];
  assign o[30730] = i[60];
  assign o[30731] = i[60];
  assign o[30732] = i[60];
  assign o[30733] = i[60];
  assign o[30734] = i[60];
  assign o[30735] = i[60];
  assign o[30736] = i[60];
  assign o[30737] = i[60];
  assign o[30738] = i[60];
  assign o[30739] = i[60];
  assign o[30740] = i[60];
  assign o[30741] = i[60];
  assign o[30742] = i[60];
  assign o[30743] = i[60];
  assign o[30744] = i[60];
  assign o[30745] = i[60];
  assign o[30746] = i[60];
  assign o[30747] = i[60];
  assign o[30748] = i[60];
  assign o[30749] = i[60];
  assign o[30750] = i[60];
  assign o[30751] = i[60];
  assign o[30752] = i[60];
  assign o[30753] = i[60];
  assign o[30754] = i[60];
  assign o[30755] = i[60];
  assign o[30756] = i[60];
  assign o[30757] = i[60];
  assign o[30758] = i[60];
  assign o[30759] = i[60];
  assign o[30760] = i[60];
  assign o[30761] = i[60];
  assign o[30762] = i[60];
  assign o[30763] = i[60];
  assign o[30764] = i[60];
  assign o[30765] = i[60];
  assign o[30766] = i[60];
  assign o[30767] = i[60];
  assign o[30768] = i[60];
  assign o[30769] = i[60];
  assign o[30770] = i[60];
  assign o[30771] = i[60];
  assign o[30772] = i[60];
  assign o[30773] = i[60];
  assign o[30774] = i[60];
  assign o[30775] = i[60];
  assign o[30776] = i[60];
  assign o[30777] = i[60];
  assign o[30778] = i[60];
  assign o[30779] = i[60];
  assign o[30780] = i[60];
  assign o[30781] = i[60];
  assign o[30782] = i[60];
  assign o[30783] = i[60];
  assign o[30784] = i[60];
  assign o[30785] = i[60];
  assign o[30786] = i[60];
  assign o[30787] = i[60];
  assign o[30788] = i[60];
  assign o[30789] = i[60];
  assign o[30790] = i[60];
  assign o[30791] = i[60];
  assign o[30792] = i[60];
  assign o[30793] = i[60];
  assign o[30794] = i[60];
  assign o[30795] = i[60];
  assign o[30796] = i[60];
  assign o[30797] = i[60];
  assign o[30798] = i[60];
  assign o[30799] = i[60];
  assign o[30800] = i[60];
  assign o[30801] = i[60];
  assign o[30802] = i[60];
  assign o[30803] = i[60];
  assign o[30804] = i[60];
  assign o[30805] = i[60];
  assign o[30806] = i[60];
  assign o[30807] = i[60];
  assign o[30808] = i[60];
  assign o[30809] = i[60];
  assign o[30810] = i[60];
  assign o[30811] = i[60];
  assign o[30812] = i[60];
  assign o[30813] = i[60];
  assign o[30814] = i[60];
  assign o[30815] = i[60];
  assign o[30816] = i[60];
  assign o[30817] = i[60];
  assign o[30818] = i[60];
  assign o[30819] = i[60];
  assign o[30820] = i[60];
  assign o[30821] = i[60];
  assign o[30822] = i[60];
  assign o[30823] = i[60];
  assign o[30824] = i[60];
  assign o[30825] = i[60];
  assign o[30826] = i[60];
  assign o[30827] = i[60];
  assign o[30828] = i[60];
  assign o[30829] = i[60];
  assign o[30830] = i[60];
  assign o[30831] = i[60];
  assign o[30832] = i[60];
  assign o[30833] = i[60];
  assign o[30834] = i[60];
  assign o[30835] = i[60];
  assign o[30836] = i[60];
  assign o[30837] = i[60];
  assign o[30838] = i[60];
  assign o[30839] = i[60];
  assign o[30840] = i[60];
  assign o[30841] = i[60];
  assign o[30842] = i[60];
  assign o[30843] = i[60];
  assign o[30844] = i[60];
  assign o[30845] = i[60];
  assign o[30846] = i[60];
  assign o[30847] = i[60];
  assign o[30848] = i[60];
  assign o[30849] = i[60];
  assign o[30850] = i[60];
  assign o[30851] = i[60];
  assign o[30852] = i[60];
  assign o[30853] = i[60];
  assign o[30854] = i[60];
  assign o[30855] = i[60];
  assign o[30856] = i[60];
  assign o[30857] = i[60];
  assign o[30858] = i[60];
  assign o[30859] = i[60];
  assign o[30860] = i[60];
  assign o[30861] = i[60];
  assign o[30862] = i[60];
  assign o[30863] = i[60];
  assign o[30864] = i[60];
  assign o[30865] = i[60];
  assign o[30866] = i[60];
  assign o[30867] = i[60];
  assign o[30868] = i[60];
  assign o[30869] = i[60];
  assign o[30870] = i[60];
  assign o[30871] = i[60];
  assign o[30872] = i[60];
  assign o[30873] = i[60];
  assign o[30874] = i[60];
  assign o[30875] = i[60];
  assign o[30876] = i[60];
  assign o[30877] = i[60];
  assign o[30878] = i[60];
  assign o[30879] = i[60];
  assign o[30880] = i[60];
  assign o[30881] = i[60];
  assign o[30882] = i[60];
  assign o[30883] = i[60];
  assign o[30884] = i[60];
  assign o[30885] = i[60];
  assign o[30886] = i[60];
  assign o[30887] = i[60];
  assign o[30888] = i[60];
  assign o[30889] = i[60];
  assign o[30890] = i[60];
  assign o[30891] = i[60];
  assign o[30892] = i[60];
  assign o[30893] = i[60];
  assign o[30894] = i[60];
  assign o[30895] = i[60];
  assign o[30896] = i[60];
  assign o[30897] = i[60];
  assign o[30898] = i[60];
  assign o[30899] = i[60];
  assign o[30900] = i[60];
  assign o[30901] = i[60];
  assign o[30902] = i[60];
  assign o[30903] = i[60];
  assign o[30904] = i[60];
  assign o[30905] = i[60];
  assign o[30906] = i[60];
  assign o[30907] = i[60];
  assign o[30908] = i[60];
  assign o[30909] = i[60];
  assign o[30910] = i[60];
  assign o[30911] = i[60];
  assign o[30912] = i[60];
  assign o[30913] = i[60];
  assign o[30914] = i[60];
  assign o[30915] = i[60];
  assign o[30916] = i[60];
  assign o[30917] = i[60];
  assign o[30918] = i[60];
  assign o[30919] = i[60];
  assign o[30920] = i[60];
  assign o[30921] = i[60];
  assign o[30922] = i[60];
  assign o[30923] = i[60];
  assign o[30924] = i[60];
  assign o[30925] = i[60];
  assign o[30926] = i[60];
  assign o[30927] = i[60];
  assign o[30928] = i[60];
  assign o[30929] = i[60];
  assign o[30930] = i[60];
  assign o[30931] = i[60];
  assign o[30932] = i[60];
  assign o[30933] = i[60];
  assign o[30934] = i[60];
  assign o[30935] = i[60];
  assign o[30936] = i[60];
  assign o[30937] = i[60];
  assign o[30938] = i[60];
  assign o[30939] = i[60];
  assign o[30940] = i[60];
  assign o[30941] = i[60];
  assign o[30942] = i[60];
  assign o[30943] = i[60];
  assign o[30944] = i[60];
  assign o[30945] = i[60];
  assign o[30946] = i[60];
  assign o[30947] = i[60];
  assign o[30948] = i[60];
  assign o[30949] = i[60];
  assign o[30950] = i[60];
  assign o[30951] = i[60];
  assign o[30952] = i[60];
  assign o[30953] = i[60];
  assign o[30954] = i[60];
  assign o[30955] = i[60];
  assign o[30956] = i[60];
  assign o[30957] = i[60];
  assign o[30958] = i[60];
  assign o[30959] = i[60];
  assign o[30960] = i[60];
  assign o[30961] = i[60];
  assign o[30962] = i[60];
  assign o[30963] = i[60];
  assign o[30964] = i[60];
  assign o[30965] = i[60];
  assign o[30966] = i[60];
  assign o[30967] = i[60];
  assign o[30968] = i[60];
  assign o[30969] = i[60];
  assign o[30970] = i[60];
  assign o[30971] = i[60];
  assign o[30972] = i[60];
  assign o[30973] = i[60];
  assign o[30974] = i[60];
  assign o[30975] = i[60];
  assign o[30976] = i[60];
  assign o[30977] = i[60];
  assign o[30978] = i[60];
  assign o[30979] = i[60];
  assign o[30980] = i[60];
  assign o[30981] = i[60];
  assign o[30982] = i[60];
  assign o[30983] = i[60];
  assign o[30984] = i[60];
  assign o[30985] = i[60];
  assign o[30986] = i[60];
  assign o[30987] = i[60];
  assign o[30988] = i[60];
  assign o[30989] = i[60];
  assign o[30990] = i[60];
  assign o[30991] = i[60];
  assign o[30992] = i[60];
  assign o[30993] = i[60];
  assign o[30994] = i[60];
  assign o[30995] = i[60];
  assign o[30996] = i[60];
  assign o[30997] = i[60];
  assign o[30998] = i[60];
  assign o[30999] = i[60];
  assign o[31000] = i[60];
  assign o[31001] = i[60];
  assign o[31002] = i[60];
  assign o[31003] = i[60];
  assign o[31004] = i[60];
  assign o[31005] = i[60];
  assign o[31006] = i[60];
  assign o[31007] = i[60];
  assign o[31008] = i[60];
  assign o[31009] = i[60];
  assign o[31010] = i[60];
  assign o[31011] = i[60];
  assign o[31012] = i[60];
  assign o[31013] = i[60];
  assign o[31014] = i[60];
  assign o[31015] = i[60];
  assign o[31016] = i[60];
  assign o[31017] = i[60];
  assign o[31018] = i[60];
  assign o[31019] = i[60];
  assign o[31020] = i[60];
  assign o[31021] = i[60];
  assign o[31022] = i[60];
  assign o[31023] = i[60];
  assign o[31024] = i[60];
  assign o[31025] = i[60];
  assign o[31026] = i[60];
  assign o[31027] = i[60];
  assign o[31028] = i[60];
  assign o[31029] = i[60];
  assign o[31030] = i[60];
  assign o[31031] = i[60];
  assign o[31032] = i[60];
  assign o[31033] = i[60];
  assign o[31034] = i[60];
  assign o[31035] = i[60];
  assign o[31036] = i[60];
  assign o[31037] = i[60];
  assign o[31038] = i[60];
  assign o[31039] = i[60];
  assign o[31040] = i[60];
  assign o[31041] = i[60];
  assign o[31042] = i[60];
  assign o[31043] = i[60];
  assign o[31044] = i[60];
  assign o[31045] = i[60];
  assign o[31046] = i[60];
  assign o[31047] = i[60];
  assign o[31048] = i[60];
  assign o[31049] = i[60];
  assign o[31050] = i[60];
  assign o[31051] = i[60];
  assign o[31052] = i[60];
  assign o[31053] = i[60];
  assign o[31054] = i[60];
  assign o[31055] = i[60];
  assign o[31056] = i[60];
  assign o[31057] = i[60];
  assign o[31058] = i[60];
  assign o[31059] = i[60];
  assign o[31060] = i[60];
  assign o[31061] = i[60];
  assign o[31062] = i[60];
  assign o[31063] = i[60];
  assign o[31064] = i[60];
  assign o[31065] = i[60];
  assign o[31066] = i[60];
  assign o[31067] = i[60];
  assign o[31068] = i[60];
  assign o[31069] = i[60];
  assign o[31070] = i[60];
  assign o[31071] = i[60];
  assign o[31072] = i[60];
  assign o[31073] = i[60];
  assign o[31074] = i[60];
  assign o[31075] = i[60];
  assign o[31076] = i[60];
  assign o[31077] = i[60];
  assign o[31078] = i[60];
  assign o[31079] = i[60];
  assign o[31080] = i[60];
  assign o[31081] = i[60];
  assign o[31082] = i[60];
  assign o[31083] = i[60];
  assign o[31084] = i[60];
  assign o[31085] = i[60];
  assign o[31086] = i[60];
  assign o[31087] = i[60];
  assign o[31088] = i[60];
  assign o[31089] = i[60];
  assign o[31090] = i[60];
  assign o[31091] = i[60];
  assign o[31092] = i[60];
  assign o[31093] = i[60];
  assign o[31094] = i[60];
  assign o[31095] = i[60];
  assign o[31096] = i[60];
  assign o[31097] = i[60];
  assign o[31098] = i[60];
  assign o[31099] = i[60];
  assign o[31100] = i[60];
  assign o[31101] = i[60];
  assign o[31102] = i[60];
  assign o[31103] = i[60];
  assign o[31104] = i[60];
  assign o[31105] = i[60];
  assign o[31106] = i[60];
  assign o[31107] = i[60];
  assign o[31108] = i[60];
  assign o[31109] = i[60];
  assign o[31110] = i[60];
  assign o[31111] = i[60];
  assign o[31112] = i[60];
  assign o[31113] = i[60];
  assign o[31114] = i[60];
  assign o[31115] = i[60];
  assign o[31116] = i[60];
  assign o[31117] = i[60];
  assign o[31118] = i[60];
  assign o[31119] = i[60];
  assign o[31120] = i[60];
  assign o[31121] = i[60];
  assign o[31122] = i[60];
  assign o[31123] = i[60];
  assign o[31124] = i[60];
  assign o[31125] = i[60];
  assign o[31126] = i[60];
  assign o[31127] = i[60];
  assign o[31128] = i[60];
  assign o[31129] = i[60];
  assign o[31130] = i[60];
  assign o[31131] = i[60];
  assign o[31132] = i[60];
  assign o[31133] = i[60];
  assign o[31134] = i[60];
  assign o[31135] = i[60];
  assign o[31136] = i[60];
  assign o[31137] = i[60];
  assign o[31138] = i[60];
  assign o[31139] = i[60];
  assign o[31140] = i[60];
  assign o[31141] = i[60];
  assign o[31142] = i[60];
  assign o[31143] = i[60];
  assign o[31144] = i[60];
  assign o[31145] = i[60];
  assign o[31146] = i[60];
  assign o[31147] = i[60];
  assign o[31148] = i[60];
  assign o[31149] = i[60];
  assign o[31150] = i[60];
  assign o[31151] = i[60];
  assign o[31152] = i[60];
  assign o[31153] = i[60];
  assign o[31154] = i[60];
  assign o[31155] = i[60];
  assign o[31156] = i[60];
  assign o[31157] = i[60];
  assign o[31158] = i[60];
  assign o[31159] = i[60];
  assign o[31160] = i[60];
  assign o[31161] = i[60];
  assign o[31162] = i[60];
  assign o[31163] = i[60];
  assign o[31164] = i[60];
  assign o[31165] = i[60];
  assign o[31166] = i[60];
  assign o[31167] = i[60];
  assign o[31168] = i[60];
  assign o[31169] = i[60];
  assign o[31170] = i[60];
  assign o[31171] = i[60];
  assign o[31172] = i[60];
  assign o[31173] = i[60];
  assign o[31174] = i[60];
  assign o[31175] = i[60];
  assign o[31176] = i[60];
  assign o[31177] = i[60];
  assign o[31178] = i[60];
  assign o[31179] = i[60];
  assign o[31180] = i[60];
  assign o[31181] = i[60];
  assign o[31182] = i[60];
  assign o[31183] = i[60];
  assign o[31184] = i[60];
  assign o[31185] = i[60];
  assign o[31186] = i[60];
  assign o[31187] = i[60];
  assign o[31188] = i[60];
  assign o[31189] = i[60];
  assign o[31190] = i[60];
  assign o[31191] = i[60];
  assign o[31192] = i[60];
  assign o[31193] = i[60];
  assign o[31194] = i[60];
  assign o[31195] = i[60];
  assign o[31196] = i[60];
  assign o[31197] = i[60];
  assign o[31198] = i[60];
  assign o[31199] = i[60];
  assign o[31200] = i[60];
  assign o[31201] = i[60];
  assign o[31202] = i[60];
  assign o[31203] = i[60];
  assign o[31204] = i[60];
  assign o[31205] = i[60];
  assign o[31206] = i[60];
  assign o[31207] = i[60];
  assign o[31208] = i[60];
  assign o[31209] = i[60];
  assign o[31210] = i[60];
  assign o[31211] = i[60];
  assign o[31212] = i[60];
  assign o[31213] = i[60];
  assign o[31214] = i[60];
  assign o[31215] = i[60];
  assign o[31216] = i[60];
  assign o[31217] = i[60];
  assign o[31218] = i[60];
  assign o[31219] = i[60];
  assign o[31220] = i[60];
  assign o[31221] = i[60];
  assign o[31222] = i[60];
  assign o[31223] = i[60];
  assign o[31224] = i[60];
  assign o[31225] = i[60];
  assign o[31226] = i[60];
  assign o[31227] = i[60];
  assign o[31228] = i[60];
  assign o[31229] = i[60];
  assign o[31230] = i[60];
  assign o[31231] = i[60];
  assign o[30208] = i[59];
  assign o[30209] = i[59];
  assign o[30210] = i[59];
  assign o[30211] = i[59];
  assign o[30212] = i[59];
  assign o[30213] = i[59];
  assign o[30214] = i[59];
  assign o[30215] = i[59];
  assign o[30216] = i[59];
  assign o[30217] = i[59];
  assign o[30218] = i[59];
  assign o[30219] = i[59];
  assign o[30220] = i[59];
  assign o[30221] = i[59];
  assign o[30222] = i[59];
  assign o[30223] = i[59];
  assign o[30224] = i[59];
  assign o[30225] = i[59];
  assign o[30226] = i[59];
  assign o[30227] = i[59];
  assign o[30228] = i[59];
  assign o[30229] = i[59];
  assign o[30230] = i[59];
  assign o[30231] = i[59];
  assign o[30232] = i[59];
  assign o[30233] = i[59];
  assign o[30234] = i[59];
  assign o[30235] = i[59];
  assign o[30236] = i[59];
  assign o[30237] = i[59];
  assign o[30238] = i[59];
  assign o[30239] = i[59];
  assign o[30240] = i[59];
  assign o[30241] = i[59];
  assign o[30242] = i[59];
  assign o[30243] = i[59];
  assign o[30244] = i[59];
  assign o[30245] = i[59];
  assign o[30246] = i[59];
  assign o[30247] = i[59];
  assign o[30248] = i[59];
  assign o[30249] = i[59];
  assign o[30250] = i[59];
  assign o[30251] = i[59];
  assign o[30252] = i[59];
  assign o[30253] = i[59];
  assign o[30254] = i[59];
  assign o[30255] = i[59];
  assign o[30256] = i[59];
  assign o[30257] = i[59];
  assign o[30258] = i[59];
  assign o[30259] = i[59];
  assign o[30260] = i[59];
  assign o[30261] = i[59];
  assign o[30262] = i[59];
  assign o[30263] = i[59];
  assign o[30264] = i[59];
  assign o[30265] = i[59];
  assign o[30266] = i[59];
  assign o[30267] = i[59];
  assign o[30268] = i[59];
  assign o[30269] = i[59];
  assign o[30270] = i[59];
  assign o[30271] = i[59];
  assign o[30272] = i[59];
  assign o[30273] = i[59];
  assign o[30274] = i[59];
  assign o[30275] = i[59];
  assign o[30276] = i[59];
  assign o[30277] = i[59];
  assign o[30278] = i[59];
  assign o[30279] = i[59];
  assign o[30280] = i[59];
  assign o[30281] = i[59];
  assign o[30282] = i[59];
  assign o[30283] = i[59];
  assign o[30284] = i[59];
  assign o[30285] = i[59];
  assign o[30286] = i[59];
  assign o[30287] = i[59];
  assign o[30288] = i[59];
  assign o[30289] = i[59];
  assign o[30290] = i[59];
  assign o[30291] = i[59];
  assign o[30292] = i[59];
  assign o[30293] = i[59];
  assign o[30294] = i[59];
  assign o[30295] = i[59];
  assign o[30296] = i[59];
  assign o[30297] = i[59];
  assign o[30298] = i[59];
  assign o[30299] = i[59];
  assign o[30300] = i[59];
  assign o[30301] = i[59];
  assign o[30302] = i[59];
  assign o[30303] = i[59];
  assign o[30304] = i[59];
  assign o[30305] = i[59];
  assign o[30306] = i[59];
  assign o[30307] = i[59];
  assign o[30308] = i[59];
  assign o[30309] = i[59];
  assign o[30310] = i[59];
  assign o[30311] = i[59];
  assign o[30312] = i[59];
  assign o[30313] = i[59];
  assign o[30314] = i[59];
  assign o[30315] = i[59];
  assign o[30316] = i[59];
  assign o[30317] = i[59];
  assign o[30318] = i[59];
  assign o[30319] = i[59];
  assign o[30320] = i[59];
  assign o[30321] = i[59];
  assign o[30322] = i[59];
  assign o[30323] = i[59];
  assign o[30324] = i[59];
  assign o[30325] = i[59];
  assign o[30326] = i[59];
  assign o[30327] = i[59];
  assign o[30328] = i[59];
  assign o[30329] = i[59];
  assign o[30330] = i[59];
  assign o[30331] = i[59];
  assign o[30332] = i[59];
  assign o[30333] = i[59];
  assign o[30334] = i[59];
  assign o[30335] = i[59];
  assign o[30336] = i[59];
  assign o[30337] = i[59];
  assign o[30338] = i[59];
  assign o[30339] = i[59];
  assign o[30340] = i[59];
  assign o[30341] = i[59];
  assign o[30342] = i[59];
  assign o[30343] = i[59];
  assign o[30344] = i[59];
  assign o[30345] = i[59];
  assign o[30346] = i[59];
  assign o[30347] = i[59];
  assign o[30348] = i[59];
  assign o[30349] = i[59];
  assign o[30350] = i[59];
  assign o[30351] = i[59];
  assign o[30352] = i[59];
  assign o[30353] = i[59];
  assign o[30354] = i[59];
  assign o[30355] = i[59];
  assign o[30356] = i[59];
  assign o[30357] = i[59];
  assign o[30358] = i[59];
  assign o[30359] = i[59];
  assign o[30360] = i[59];
  assign o[30361] = i[59];
  assign o[30362] = i[59];
  assign o[30363] = i[59];
  assign o[30364] = i[59];
  assign o[30365] = i[59];
  assign o[30366] = i[59];
  assign o[30367] = i[59];
  assign o[30368] = i[59];
  assign o[30369] = i[59];
  assign o[30370] = i[59];
  assign o[30371] = i[59];
  assign o[30372] = i[59];
  assign o[30373] = i[59];
  assign o[30374] = i[59];
  assign o[30375] = i[59];
  assign o[30376] = i[59];
  assign o[30377] = i[59];
  assign o[30378] = i[59];
  assign o[30379] = i[59];
  assign o[30380] = i[59];
  assign o[30381] = i[59];
  assign o[30382] = i[59];
  assign o[30383] = i[59];
  assign o[30384] = i[59];
  assign o[30385] = i[59];
  assign o[30386] = i[59];
  assign o[30387] = i[59];
  assign o[30388] = i[59];
  assign o[30389] = i[59];
  assign o[30390] = i[59];
  assign o[30391] = i[59];
  assign o[30392] = i[59];
  assign o[30393] = i[59];
  assign o[30394] = i[59];
  assign o[30395] = i[59];
  assign o[30396] = i[59];
  assign o[30397] = i[59];
  assign o[30398] = i[59];
  assign o[30399] = i[59];
  assign o[30400] = i[59];
  assign o[30401] = i[59];
  assign o[30402] = i[59];
  assign o[30403] = i[59];
  assign o[30404] = i[59];
  assign o[30405] = i[59];
  assign o[30406] = i[59];
  assign o[30407] = i[59];
  assign o[30408] = i[59];
  assign o[30409] = i[59];
  assign o[30410] = i[59];
  assign o[30411] = i[59];
  assign o[30412] = i[59];
  assign o[30413] = i[59];
  assign o[30414] = i[59];
  assign o[30415] = i[59];
  assign o[30416] = i[59];
  assign o[30417] = i[59];
  assign o[30418] = i[59];
  assign o[30419] = i[59];
  assign o[30420] = i[59];
  assign o[30421] = i[59];
  assign o[30422] = i[59];
  assign o[30423] = i[59];
  assign o[30424] = i[59];
  assign o[30425] = i[59];
  assign o[30426] = i[59];
  assign o[30427] = i[59];
  assign o[30428] = i[59];
  assign o[30429] = i[59];
  assign o[30430] = i[59];
  assign o[30431] = i[59];
  assign o[30432] = i[59];
  assign o[30433] = i[59];
  assign o[30434] = i[59];
  assign o[30435] = i[59];
  assign o[30436] = i[59];
  assign o[30437] = i[59];
  assign o[30438] = i[59];
  assign o[30439] = i[59];
  assign o[30440] = i[59];
  assign o[30441] = i[59];
  assign o[30442] = i[59];
  assign o[30443] = i[59];
  assign o[30444] = i[59];
  assign o[30445] = i[59];
  assign o[30446] = i[59];
  assign o[30447] = i[59];
  assign o[30448] = i[59];
  assign o[30449] = i[59];
  assign o[30450] = i[59];
  assign o[30451] = i[59];
  assign o[30452] = i[59];
  assign o[30453] = i[59];
  assign o[30454] = i[59];
  assign o[30455] = i[59];
  assign o[30456] = i[59];
  assign o[30457] = i[59];
  assign o[30458] = i[59];
  assign o[30459] = i[59];
  assign o[30460] = i[59];
  assign o[30461] = i[59];
  assign o[30462] = i[59];
  assign o[30463] = i[59];
  assign o[30464] = i[59];
  assign o[30465] = i[59];
  assign o[30466] = i[59];
  assign o[30467] = i[59];
  assign o[30468] = i[59];
  assign o[30469] = i[59];
  assign o[30470] = i[59];
  assign o[30471] = i[59];
  assign o[30472] = i[59];
  assign o[30473] = i[59];
  assign o[30474] = i[59];
  assign o[30475] = i[59];
  assign o[30476] = i[59];
  assign o[30477] = i[59];
  assign o[30478] = i[59];
  assign o[30479] = i[59];
  assign o[30480] = i[59];
  assign o[30481] = i[59];
  assign o[30482] = i[59];
  assign o[30483] = i[59];
  assign o[30484] = i[59];
  assign o[30485] = i[59];
  assign o[30486] = i[59];
  assign o[30487] = i[59];
  assign o[30488] = i[59];
  assign o[30489] = i[59];
  assign o[30490] = i[59];
  assign o[30491] = i[59];
  assign o[30492] = i[59];
  assign o[30493] = i[59];
  assign o[30494] = i[59];
  assign o[30495] = i[59];
  assign o[30496] = i[59];
  assign o[30497] = i[59];
  assign o[30498] = i[59];
  assign o[30499] = i[59];
  assign o[30500] = i[59];
  assign o[30501] = i[59];
  assign o[30502] = i[59];
  assign o[30503] = i[59];
  assign o[30504] = i[59];
  assign o[30505] = i[59];
  assign o[30506] = i[59];
  assign o[30507] = i[59];
  assign o[30508] = i[59];
  assign o[30509] = i[59];
  assign o[30510] = i[59];
  assign o[30511] = i[59];
  assign o[30512] = i[59];
  assign o[30513] = i[59];
  assign o[30514] = i[59];
  assign o[30515] = i[59];
  assign o[30516] = i[59];
  assign o[30517] = i[59];
  assign o[30518] = i[59];
  assign o[30519] = i[59];
  assign o[30520] = i[59];
  assign o[30521] = i[59];
  assign o[30522] = i[59];
  assign o[30523] = i[59];
  assign o[30524] = i[59];
  assign o[30525] = i[59];
  assign o[30526] = i[59];
  assign o[30527] = i[59];
  assign o[30528] = i[59];
  assign o[30529] = i[59];
  assign o[30530] = i[59];
  assign o[30531] = i[59];
  assign o[30532] = i[59];
  assign o[30533] = i[59];
  assign o[30534] = i[59];
  assign o[30535] = i[59];
  assign o[30536] = i[59];
  assign o[30537] = i[59];
  assign o[30538] = i[59];
  assign o[30539] = i[59];
  assign o[30540] = i[59];
  assign o[30541] = i[59];
  assign o[30542] = i[59];
  assign o[30543] = i[59];
  assign o[30544] = i[59];
  assign o[30545] = i[59];
  assign o[30546] = i[59];
  assign o[30547] = i[59];
  assign o[30548] = i[59];
  assign o[30549] = i[59];
  assign o[30550] = i[59];
  assign o[30551] = i[59];
  assign o[30552] = i[59];
  assign o[30553] = i[59];
  assign o[30554] = i[59];
  assign o[30555] = i[59];
  assign o[30556] = i[59];
  assign o[30557] = i[59];
  assign o[30558] = i[59];
  assign o[30559] = i[59];
  assign o[30560] = i[59];
  assign o[30561] = i[59];
  assign o[30562] = i[59];
  assign o[30563] = i[59];
  assign o[30564] = i[59];
  assign o[30565] = i[59];
  assign o[30566] = i[59];
  assign o[30567] = i[59];
  assign o[30568] = i[59];
  assign o[30569] = i[59];
  assign o[30570] = i[59];
  assign o[30571] = i[59];
  assign o[30572] = i[59];
  assign o[30573] = i[59];
  assign o[30574] = i[59];
  assign o[30575] = i[59];
  assign o[30576] = i[59];
  assign o[30577] = i[59];
  assign o[30578] = i[59];
  assign o[30579] = i[59];
  assign o[30580] = i[59];
  assign o[30581] = i[59];
  assign o[30582] = i[59];
  assign o[30583] = i[59];
  assign o[30584] = i[59];
  assign o[30585] = i[59];
  assign o[30586] = i[59];
  assign o[30587] = i[59];
  assign o[30588] = i[59];
  assign o[30589] = i[59];
  assign o[30590] = i[59];
  assign o[30591] = i[59];
  assign o[30592] = i[59];
  assign o[30593] = i[59];
  assign o[30594] = i[59];
  assign o[30595] = i[59];
  assign o[30596] = i[59];
  assign o[30597] = i[59];
  assign o[30598] = i[59];
  assign o[30599] = i[59];
  assign o[30600] = i[59];
  assign o[30601] = i[59];
  assign o[30602] = i[59];
  assign o[30603] = i[59];
  assign o[30604] = i[59];
  assign o[30605] = i[59];
  assign o[30606] = i[59];
  assign o[30607] = i[59];
  assign o[30608] = i[59];
  assign o[30609] = i[59];
  assign o[30610] = i[59];
  assign o[30611] = i[59];
  assign o[30612] = i[59];
  assign o[30613] = i[59];
  assign o[30614] = i[59];
  assign o[30615] = i[59];
  assign o[30616] = i[59];
  assign o[30617] = i[59];
  assign o[30618] = i[59];
  assign o[30619] = i[59];
  assign o[30620] = i[59];
  assign o[30621] = i[59];
  assign o[30622] = i[59];
  assign o[30623] = i[59];
  assign o[30624] = i[59];
  assign o[30625] = i[59];
  assign o[30626] = i[59];
  assign o[30627] = i[59];
  assign o[30628] = i[59];
  assign o[30629] = i[59];
  assign o[30630] = i[59];
  assign o[30631] = i[59];
  assign o[30632] = i[59];
  assign o[30633] = i[59];
  assign o[30634] = i[59];
  assign o[30635] = i[59];
  assign o[30636] = i[59];
  assign o[30637] = i[59];
  assign o[30638] = i[59];
  assign o[30639] = i[59];
  assign o[30640] = i[59];
  assign o[30641] = i[59];
  assign o[30642] = i[59];
  assign o[30643] = i[59];
  assign o[30644] = i[59];
  assign o[30645] = i[59];
  assign o[30646] = i[59];
  assign o[30647] = i[59];
  assign o[30648] = i[59];
  assign o[30649] = i[59];
  assign o[30650] = i[59];
  assign o[30651] = i[59];
  assign o[30652] = i[59];
  assign o[30653] = i[59];
  assign o[30654] = i[59];
  assign o[30655] = i[59];
  assign o[30656] = i[59];
  assign o[30657] = i[59];
  assign o[30658] = i[59];
  assign o[30659] = i[59];
  assign o[30660] = i[59];
  assign o[30661] = i[59];
  assign o[30662] = i[59];
  assign o[30663] = i[59];
  assign o[30664] = i[59];
  assign o[30665] = i[59];
  assign o[30666] = i[59];
  assign o[30667] = i[59];
  assign o[30668] = i[59];
  assign o[30669] = i[59];
  assign o[30670] = i[59];
  assign o[30671] = i[59];
  assign o[30672] = i[59];
  assign o[30673] = i[59];
  assign o[30674] = i[59];
  assign o[30675] = i[59];
  assign o[30676] = i[59];
  assign o[30677] = i[59];
  assign o[30678] = i[59];
  assign o[30679] = i[59];
  assign o[30680] = i[59];
  assign o[30681] = i[59];
  assign o[30682] = i[59];
  assign o[30683] = i[59];
  assign o[30684] = i[59];
  assign o[30685] = i[59];
  assign o[30686] = i[59];
  assign o[30687] = i[59];
  assign o[30688] = i[59];
  assign o[30689] = i[59];
  assign o[30690] = i[59];
  assign o[30691] = i[59];
  assign o[30692] = i[59];
  assign o[30693] = i[59];
  assign o[30694] = i[59];
  assign o[30695] = i[59];
  assign o[30696] = i[59];
  assign o[30697] = i[59];
  assign o[30698] = i[59];
  assign o[30699] = i[59];
  assign o[30700] = i[59];
  assign o[30701] = i[59];
  assign o[30702] = i[59];
  assign o[30703] = i[59];
  assign o[30704] = i[59];
  assign o[30705] = i[59];
  assign o[30706] = i[59];
  assign o[30707] = i[59];
  assign o[30708] = i[59];
  assign o[30709] = i[59];
  assign o[30710] = i[59];
  assign o[30711] = i[59];
  assign o[30712] = i[59];
  assign o[30713] = i[59];
  assign o[30714] = i[59];
  assign o[30715] = i[59];
  assign o[30716] = i[59];
  assign o[30717] = i[59];
  assign o[30718] = i[59];
  assign o[30719] = i[59];
  assign o[29696] = i[58];
  assign o[29697] = i[58];
  assign o[29698] = i[58];
  assign o[29699] = i[58];
  assign o[29700] = i[58];
  assign o[29701] = i[58];
  assign o[29702] = i[58];
  assign o[29703] = i[58];
  assign o[29704] = i[58];
  assign o[29705] = i[58];
  assign o[29706] = i[58];
  assign o[29707] = i[58];
  assign o[29708] = i[58];
  assign o[29709] = i[58];
  assign o[29710] = i[58];
  assign o[29711] = i[58];
  assign o[29712] = i[58];
  assign o[29713] = i[58];
  assign o[29714] = i[58];
  assign o[29715] = i[58];
  assign o[29716] = i[58];
  assign o[29717] = i[58];
  assign o[29718] = i[58];
  assign o[29719] = i[58];
  assign o[29720] = i[58];
  assign o[29721] = i[58];
  assign o[29722] = i[58];
  assign o[29723] = i[58];
  assign o[29724] = i[58];
  assign o[29725] = i[58];
  assign o[29726] = i[58];
  assign o[29727] = i[58];
  assign o[29728] = i[58];
  assign o[29729] = i[58];
  assign o[29730] = i[58];
  assign o[29731] = i[58];
  assign o[29732] = i[58];
  assign o[29733] = i[58];
  assign o[29734] = i[58];
  assign o[29735] = i[58];
  assign o[29736] = i[58];
  assign o[29737] = i[58];
  assign o[29738] = i[58];
  assign o[29739] = i[58];
  assign o[29740] = i[58];
  assign o[29741] = i[58];
  assign o[29742] = i[58];
  assign o[29743] = i[58];
  assign o[29744] = i[58];
  assign o[29745] = i[58];
  assign o[29746] = i[58];
  assign o[29747] = i[58];
  assign o[29748] = i[58];
  assign o[29749] = i[58];
  assign o[29750] = i[58];
  assign o[29751] = i[58];
  assign o[29752] = i[58];
  assign o[29753] = i[58];
  assign o[29754] = i[58];
  assign o[29755] = i[58];
  assign o[29756] = i[58];
  assign o[29757] = i[58];
  assign o[29758] = i[58];
  assign o[29759] = i[58];
  assign o[29760] = i[58];
  assign o[29761] = i[58];
  assign o[29762] = i[58];
  assign o[29763] = i[58];
  assign o[29764] = i[58];
  assign o[29765] = i[58];
  assign o[29766] = i[58];
  assign o[29767] = i[58];
  assign o[29768] = i[58];
  assign o[29769] = i[58];
  assign o[29770] = i[58];
  assign o[29771] = i[58];
  assign o[29772] = i[58];
  assign o[29773] = i[58];
  assign o[29774] = i[58];
  assign o[29775] = i[58];
  assign o[29776] = i[58];
  assign o[29777] = i[58];
  assign o[29778] = i[58];
  assign o[29779] = i[58];
  assign o[29780] = i[58];
  assign o[29781] = i[58];
  assign o[29782] = i[58];
  assign o[29783] = i[58];
  assign o[29784] = i[58];
  assign o[29785] = i[58];
  assign o[29786] = i[58];
  assign o[29787] = i[58];
  assign o[29788] = i[58];
  assign o[29789] = i[58];
  assign o[29790] = i[58];
  assign o[29791] = i[58];
  assign o[29792] = i[58];
  assign o[29793] = i[58];
  assign o[29794] = i[58];
  assign o[29795] = i[58];
  assign o[29796] = i[58];
  assign o[29797] = i[58];
  assign o[29798] = i[58];
  assign o[29799] = i[58];
  assign o[29800] = i[58];
  assign o[29801] = i[58];
  assign o[29802] = i[58];
  assign o[29803] = i[58];
  assign o[29804] = i[58];
  assign o[29805] = i[58];
  assign o[29806] = i[58];
  assign o[29807] = i[58];
  assign o[29808] = i[58];
  assign o[29809] = i[58];
  assign o[29810] = i[58];
  assign o[29811] = i[58];
  assign o[29812] = i[58];
  assign o[29813] = i[58];
  assign o[29814] = i[58];
  assign o[29815] = i[58];
  assign o[29816] = i[58];
  assign o[29817] = i[58];
  assign o[29818] = i[58];
  assign o[29819] = i[58];
  assign o[29820] = i[58];
  assign o[29821] = i[58];
  assign o[29822] = i[58];
  assign o[29823] = i[58];
  assign o[29824] = i[58];
  assign o[29825] = i[58];
  assign o[29826] = i[58];
  assign o[29827] = i[58];
  assign o[29828] = i[58];
  assign o[29829] = i[58];
  assign o[29830] = i[58];
  assign o[29831] = i[58];
  assign o[29832] = i[58];
  assign o[29833] = i[58];
  assign o[29834] = i[58];
  assign o[29835] = i[58];
  assign o[29836] = i[58];
  assign o[29837] = i[58];
  assign o[29838] = i[58];
  assign o[29839] = i[58];
  assign o[29840] = i[58];
  assign o[29841] = i[58];
  assign o[29842] = i[58];
  assign o[29843] = i[58];
  assign o[29844] = i[58];
  assign o[29845] = i[58];
  assign o[29846] = i[58];
  assign o[29847] = i[58];
  assign o[29848] = i[58];
  assign o[29849] = i[58];
  assign o[29850] = i[58];
  assign o[29851] = i[58];
  assign o[29852] = i[58];
  assign o[29853] = i[58];
  assign o[29854] = i[58];
  assign o[29855] = i[58];
  assign o[29856] = i[58];
  assign o[29857] = i[58];
  assign o[29858] = i[58];
  assign o[29859] = i[58];
  assign o[29860] = i[58];
  assign o[29861] = i[58];
  assign o[29862] = i[58];
  assign o[29863] = i[58];
  assign o[29864] = i[58];
  assign o[29865] = i[58];
  assign o[29866] = i[58];
  assign o[29867] = i[58];
  assign o[29868] = i[58];
  assign o[29869] = i[58];
  assign o[29870] = i[58];
  assign o[29871] = i[58];
  assign o[29872] = i[58];
  assign o[29873] = i[58];
  assign o[29874] = i[58];
  assign o[29875] = i[58];
  assign o[29876] = i[58];
  assign o[29877] = i[58];
  assign o[29878] = i[58];
  assign o[29879] = i[58];
  assign o[29880] = i[58];
  assign o[29881] = i[58];
  assign o[29882] = i[58];
  assign o[29883] = i[58];
  assign o[29884] = i[58];
  assign o[29885] = i[58];
  assign o[29886] = i[58];
  assign o[29887] = i[58];
  assign o[29888] = i[58];
  assign o[29889] = i[58];
  assign o[29890] = i[58];
  assign o[29891] = i[58];
  assign o[29892] = i[58];
  assign o[29893] = i[58];
  assign o[29894] = i[58];
  assign o[29895] = i[58];
  assign o[29896] = i[58];
  assign o[29897] = i[58];
  assign o[29898] = i[58];
  assign o[29899] = i[58];
  assign o[29900] = i[58];
  assign o[29901] = i[58];
  assign o[29902] = i[58];
  assign o[29903] = i[58];
  assign o[29904] = i[58];
  assign o[29905] = i[58];
  assign o[29906] = i[58];
  assign o[29907] = i[58];
  assign o[29908] = i[58];
  assign o[29909] = i[58];
  assign o[29910] = i[58];
  assign o[29911] = i[58];
  assign o[29912] = i[58];
  assign o[29913] = i[58];
  assign o[29914] = i[58];
  assign o[29915] = i[58];
  assign o[29916] = i[58];
  assign o[29917] = i[58];
  assign o[29918] = i[58];
  assign o[29919] = i[58];
  assign o[29920] = i[58];
  assign o[29921] = i[58];
  assign o[29922] = i[58];
  assign o[29923] = i[58];
  assign o[29924] = i[58];
  assign o[29925] = i[58];
  assign o[29926] = i[58];
  assign o[29927] = i[58];
  assign o[29928] = i[58];
  assign o[29929] = i[58];
  assign o[29930] = i[58];
  assign o[29931] = i[58];
  assign o[29932] = i[58];
  assign o[29933] = i[58];
  assign o[29934] = i[58];
  assign o[29935] = i[58];
  assign o[29936] = i[58];
  assign o[29937] = i[58];
  assign o[29938] = i[58];
  assign o[29939] = i[58];
  assign o[29940] = i[58];
  assign o[29941] = i[58];
  assign o[29942] = i[58];
  assign o[29943] = i[58];
  assign o[29944] = i[58];
  assign o[29945] = i[58];
  assign o[29946] = i[58];
  assign o[29947] = i[58];
  assign o[29948] = i[58];
  assign o[29949] = i[58];
  assign o[29950] = i[58];
  assign o[29951] = i[58];
  assign o[29952] = i[58];
  assign o[29953] = i[58];
  assign o[29954] = i[58];
  assign o[29955] = i[58];
  assign o[29956] = i[58];
  assign o[29957] = i[58];
  assign o[29958] = i[58];
  assign o[29959] = i[58];
  assign o[29960] = i[58];
  assign o[29961] = i[58];
  assign o[29962] = i[58];
  assign o[29963] = i[58];
  assign o[29964] = i[58];
  assign o[29965] = i[58];
  assign o[29966] = i[58];
  assign o[29967] = i[58];
  assign o[29968] = i[58];
  assign o[29969] = i[58];
  assign o[29970] = i[58];
  assign o[29971] = i[58];
  assign o[29972] = i[58];
  assign o[29973] = i[58];
  assign o[29974] = i[58];
  assign o[29975] = i[58];
  assign o[29976] = i[58];
  assign o[29977] = i[58];
  assign o[29978] = i[58];
  assign o[29979] = i[58];
  assign o[29980] = i[58];
  assign o[29981] = i[58];
  assign o[29982] = i[58];
  assign o[29983] = i[58];
  assign o[29984] = i[58];
  assign o[29985] = i[58];
  assign o[29986] = i[58];
  assign o[29987] = i[58];
  assign o[29988] = i[58];
  assign o[29989] = i[58];
  assign o[29990] = i[58];
  assign o[29991] = i[58];
  assign o[29992] = i[58];
  assign o[29993] = i[58];
  assign o[29994] = i[58];
  assign o[29995] = i[58];
  assign o[29996] = i[58];
  assign o[29997] = i[58];
  assign o[29998] = i[58];
  assign o[29999] = i[58];
  assign o[30000] = i[58];
  assign o[30001] = i[58];
  assign o[30002] = i[58];
  assign o[30003] = i[58];
  assign o[30004] = i[58];
  assign o[30005] = i[58];
  assign o[30006] = i[58];
  assign o[30007] = i[58];
  assign o[30008] = i[58];
  assign o[30009] = i[58];
  assign o[30010] = i[58];
  assign o[30011] = i[58];
  assign o[30012] = i[58];
  assign o[30013] = i[58];
  assign o[30014] = i[58];
  assign o[30015] = i[58];
  assign o[30016] = i[58];
  assign o[30017] = i[58];
  assign o[30018] = i[58];
  assign o[30019] = i[58];
  assign o[30020] = i[58];
  assign o[30021] = i[58];
  assign o[30022] = i[58];
  assign o[30023] = i[58];
  assign o[30024] = i[58];
  assign o[30025] = i[58];
  assign o[30026] = i[58];
  assign o[30027] = i[58];
  assign o[30028] = i[58];
  assign o[30029] = i[58];
  assign o[30030] = i[58];
  assign o[30031] = i[58];
  assign o[30032] = i[58];
  assign o[30033] = i[58];
  assign o[30034] = i[58];
  assign o[30035] = i[58];
  assign o[30036] = i[58];
  assign o[30037] = i[58];
  assign o[30038] = i[58];
  assign o[30039] = i[58];
  assign o[30040] = i[58];
  assign o[30041] = i[58];
  assign o[30042] = i[58];
  assign o[30043] = i[58];
  assign o[30044] = i[58];
  assign o[30045] = i[58];
  assign o[30046] = i[58];
  assign o[30047] = i[58];
  assign o[30048] = i[58];
  assign o[30049] = i[58];
  assign o[30050] = i[58];
  assign o[30051] = i[58];
  assign o[30052] = i[58];
  assign o[30053] = i[58];
  assign o[30054] = i[58];
  assign o[30055] = i[58];
  assign o[30056] = i[58];
  assign o[30057] = i[58];
  assign o[30058] = i[58];
  assign o[30059] = i[58];
  assign o[30060] = i[58];
  assign o[30061] = i[58];
  assign o[30062] = i[58];
  assign o[30063] = i[58];
  assign o[30064] = i[58];
  assign o[30065] = i[58];
  assign o[30066] = i[58];
  assign o[30067] = i[58];
  assign o[30068] = i[58];
  assign o[30069] = i[58];
  assign o[30070] = i[58];
  assign o[30071] = i[58];
  assign o[30072] = i[58];
  assign o[30073] = i[58];
  assign o[30074] = i[58];
  assign o[30075] = i[58];
  assign o[30076] = i[58];
  assign o[30077] = i[58];
  assign o[30078] = i[58];
  assign o[30079] = i[58];
  assign o[30080] = i[58];
  assign o[30081] = i[58];
  assign o[30082] = i[58];
  assign o[30083] = i[58];
  assign o[30084] = i[58];
  assign o[30085] = i[58];
  assign o[30086] = i[58];
  assign o[30087] = i[58];
  assign o[30088] = i[58];
  assign o[30089] = i[58];
  assign o[30090] = i[58];
  assign o[30091] = i[58];
  assign o[30092] = i[58];
  assign o[30093] = i[58];
  assign o[30094] = i[58];
  assign o[30095] = i[58];
  assign o[30096] = i[58];
  assign o[30097] = i[58];
  assign o[30098] = i[58];
  assign o[30099] = i[58];
  assign o[30100] = i[58];
  assign o[30101] = i[58];
  assign o[30102] = i[58];
  assign o[30103] = i[58];
  assign o[30104] = i[58];
  assign o[30105] = i[58];
  assign o[30106] = i[58];
  assign o[30107] = i[58];
  assign o[30108] = i[58];
  assign o[30109] = i[58];
  assign o[30110] = i[58];
  assign o[30111] = i[58];
  assign o[30112] = i[58];
  assign o[30113] = i[58];
  assign o[30114] = i[58];
  assign o[30115] = i[58];
  assign o[30116] = i[58];
  assign o[30117] = i[58];
  assign o[30118] = i[58];
  assign o[30119] = i[58];
  assign o[30120] = i[58];
  assign o[30121] = i[58];
  assign o[30122] = i[58];
  assign o[30123] = i[58];
  assign o[30124] = i[58];
  assign o[30125] = i[58];
  assign o[30126] = i[58];
  assign o[30127] = i[58];
  assign o[30128] = i[58];
  assign o[30129] = i[58];
  assign o[30130] = i[58];
  assign o[30131] = i[58];
  assign o[30132] = i[58];
  assign o[30133] = i[58];
  assign o[30134] = i[58];
  assign o[30135] = i[58];
  assign o[30136] = i[58];
  assign o[30137] = i[58];
  assign o[30138] = i[58];
  assign o[30139] = i[58];
  assign o[30140] = i[58];
  assign o[30141] = i[58];
  assign o[30142] = i[58];
  assign o[30143] = i[58];
  assign o[30144] = i[58];
  assign o[30145] = i[58];
  assign o[30146] = i[58];
  assign o[30147] = i[58];
  assign o[30148] = i[58];
  assign o[30149] = i[58];
  assign o[30150] = i[58];
  assign o[30151] = i[58];
  assign o[30152] = i[58];
  assign o[30153] = i[58];
  assign o[30154] = i[58];
  assign o[30155] = i[58];
  assign o[30156] = i[58];
  assign o[30157] = i[58];
  assign o[30158] = i[58];
  assign o[30159] = i[58];
  assign o[30160] = i[58];
  assign o[30161] = i[58];
  assign o[30162] = i[58];
  assign o[30163] = i[58];
  assign o[30164] = i[58];
  assign o[30165] = i[58];
  assign o[30166] = i[58];
  assign o[30167] = i[58];
  assign o[30168] = i[58];
  assign o[30169] = i[58];
  assign o[30170] = i[58];
  assign o[30171] = i[58];
  assign o[30172] = i[58];
  assign o[30173] = i[58];
  assign o[30174] = i[58];
  assign o[30175] = i[58];
  assign o[30176] = i[58];
  assign o[30177] = i[58];
  assign o[30178] = i[58];
  assign o[30179] = i[58];
  assign o[30180] = i[58];
  assign o[30181] = i[58];
  assign o[30182] = i[58];
  assign o[30183] = i[58];
  assign o[30184] = i[58];
  assign o[30185] = i[58];
  assign o[30186] = i[58];
  assign o[30187] = i[58];
  assign o[30188] = i[58];
  assign o[30189] = i[58];
  assign o[30190] = i[58];
  assign o[30191] = i[58];
  assign o[30192] = i[58];
  assign o[30193] = i[58];
  assign o[30194] = i[58];
  assign o[30195] = i[58];
  assign o[30196] = i[58];
  assign o[30197] = i[58];
  assign o[30198] = i[58];
  assign o[30199] = i[58];
  assign o[30200] = i[58];
  assign o[30201] = i[58];
  assign o[30202] = i[58];
  assign o[30203] = i[58];
  assign o[30204] = i[58];
  assign o[30205] = i[58];
  assign o[30206] = i[58];
  assign o[30207] = i[58];
  assign o[29184] = i[57];
  assign o[29185] = i[57];
  assign o[29186] = i[57];
  assign o[29187] = i[57];
  assign o[29188] = i[57];
  assign o[29189] = i[57];
  assign o[29190] = i[57];
  assign o[29191] = i[57];
  assign o[29192] = i[57];
  assign o[29193] = i[57];
  assign o[29194] = i[57];
  assign o[29195] = i[57];
  assign o[29196] = i[57];
  assign o[29197] = i[57];
  assign o[29198] = i[57];
  assign o[29199] = i[57];
  assign o[29200] = i[57];
  assign o[29201] = i[57];
  assign o[29202] = i[57];
  assign o[29203] = i[57];
  assign o[29204] = i[57];
  assign o[29205] = i[57];
  assign o[29206] = i[57];
  assign o[29207] = i[57];
  assign o[29208] = i[57];
  assign o[29209] = i[57];
  assign o[29210] = i[57];
  assign o[29211] = i[57];
  assign o[29212] = i[57];
  assign o[29213] = i[57];
  assign o[29214] = i[57];
  assign o[29215] = i[57];
  assign o[29216] = i[57];
  assign o[29217] = i[57];
  assign o[29218] = i[57];
  assign o[29219] = i[57];
  assign o[29220] = i[57];
  assign o[29221] = i[57];
  assign o[29222] = i[57];
  assign o[29223] = i[57];
  assign o[29224] = i[57];
  assign o[29225] = i[57];
  assign o[29226] = i[57];
  assign o[29227] = i[57];
  assign o[29228] = i[57];
  assign o[29229] = i[57];
  assign o[29230] = i[57];
  assign o[29231] = i[57];
  assign o[29232] = i[57];
  assign o[29233] = i[57];
  assign o[29234] = i[57];
  assign o[29235] = i[57];
  assign o[29236] = i[57];
  assign o[29237] = i[57];
  assign o[29238] = i[57];
  assign o[29239] = i[57];
  assign o[29240] = i[57];
  assign o[29241] = i[57];
  assign o[29242] = i[57];
  assign o[29243] = i[57];
  assign o[29244] = i[57];
  assign o[29245] = i[57];
  assign o[29246] = i[57];
  assign o[29247] = i[57];
  assign o[29248] = i[57];
  assign o[29249] = i[57];
  assign o[29250] = i[57];
  assign o[29251] = i[57];
  assign o[29252] = i[57];
  assign o[29253] = i[57];
  assign o[29254] = i[57];
  assign o[29255] = i[57];
  assign o[29256] = i[57];
  assign o[29257] = i[57];
  assign o[29258] = i[57];
  assign o[29259] = i[57];
  assign o[29260] = i[57];
  assign o[29261] = i[57];
  assign o[29262] = i[57];
  assign o[29263] = i[57];
  assign o[29264] = i[57];
  assign o[29265] = i[57];
  assign o[29266] = i[57];
  assign o[29267] = i[57];
  assign o[29268] = i[57];
  assign o[29269] = i[57];
  assign o[29270] = i[57];
  assign o[29271] = i[57];
  assign o[29272] = i[57];
  assign o[29273] = i[57];
  assign o[29274] = i[57];
  assign o[29275] = i[57];
  assign o[29276] = i[57];
  assign o[29277] = i[57];
  assign o[29278] = i[57];
  assign o[29279] = i[57];
  assign o[29280] = i[57];
  assign o[29281] = i[57];
  assign o[29282] = i[57];
  assign o[29283] = i[57];
  assign o[29284] = i[57];
  assign o[29285] = i[57];
  assign o[29286] = i[57];
  assign o[29287] = i[57];
  assign o[29288] = i[57];
  assign o[29289] = i[57];
  assign o[29290] = i[57];
  assign o[29291] = i[57];
  assign o[29292] = i[57];
  assign o[29293] = i[57];
  assign o[29294] = i[57];
  assign o[29295] = i[57];
  assign o[29296] = i[57];
  assign o[29297] = i[57];
  assign o[29298] = i[57];
  assign o[29299] = i[57];
  assign o[29300] = i[57];
  assign o[29301] = i[57];
  assign o[29302] = i[57];
  assign o[29303] = i[57];
  assign o[29304] = i[57];
  assign o[29305] = i[57];
  assign o[29306] = i[57];
  assign o[29307] = i[57];
  assign o[29308] = i[57];
  assign o[29309] = i[57];
  assign o[29310] = i[57];
  assign o[29311] = i[57];
  assign o[29312] = i[57];
  assign o[29313] = i[57];
  assign o[29314] = i[57];
  assign o[29315] = i[57];
  assign o[29316] = i[57];
  assign o[29317] = i[57];
  assign o[29318] = i[57];
  assign o[29319] = i[57];
  assign o[29320] = i[57];
  assign o[29321] = i[57];
  assign o[29322] = i[57];
  assign o[29323] = i[57];
  assign o[29324] = i[57];
  assign o[29325] = i[57];
  assign o[29326] = i[57];
  assign o[29327] = i[57];
  assign o[29328] = i[57];
  assign o[29329] = i[57];
  assign o[29330] = i[57];
  assign o[29331] = i[57];
  assign o[29332] = i[57];
  assign o[29333] = i[57];
  assign o[29334] = i[57];
  assign o[29335] = i[57];
  assign o[29336] = i[57];
  assign o[29337] = i[57];
  assign o[29338] = i[57];
  assign o[29339] = i[57];
  assign o[29340] = i[57];
  assign o[29341] = i[57];
  assign o[29342] = i[57];
  assign o[29343] = i[57];
  assign o[29344] = i[57];
  assign o[29345] = i[57];
  assign o[29346] = i[57];
  assign o[29347] = i[57];
  assign o[29348] = i[57];
  assign o[29349] = i[57];
  assign o[29350] = i[57];
  assign o[29351] = i[57];
  assign o[29352] = i[57];
  assign o[29353] = i[57];
  assign o[29354] = i[57];
  assign o[29355] = i[57];
  assign o[29356] = i[57];
  assign o[29357] = i[57];
  assign o[29358] = i[57];
  assign o[29359] = i[57];
  assign o[29360] = i[57];
  assign o[29361] = i[57];
  assign o[29362] = i[57];
  assign o[29363] = i[57];
  assign o[29364] = i[57];
  assign o[29365] = i[57];
  assign o[29366] = i[57];
  assign o[29367] = i[57];
  assign o[29368] = i[57];
  assign o[29369] = i[57];
  assign o[29370] = i[57];
  assign o[29371] = i[57];
  assign o[29372] = i[57];
  assign o[29373] = i[57];
  assign o[29374] = i[57];
  assign o[29375] = i[57];
  assign o[29376] = i[57];
  assign o[29377] = i[57];
  assign o[29378] = i[57];
  assign o[29379] = i[57];
  assign o[29380] = i[57];
  assign o[29381] = i[57];
  assign o[29382] = i[57];
  assign o[29383] = i[57];
  assign o[29384] = i[57];
  assign o[29385] = i[57];
  assign o[29386] = i[57];
  assign o[29387] = i[57];
  assign o[29388] = i[57];
  assign o[29389] = i[57];
  assign o[29390] = i[57];
  assign o[29391] = i[57];
  assign o[29392] = i[57];
  assign o[29393] = i[57];
  assign o[29394] = i[57];
  assign o[29395] = i[57];
  assign o[29396] = i[57];
  assign o[29397] = i[57];
  assign o[29398] = i[57];
  assign o[29399] = i[57];
  assign o[29400] = i[57];
  assign o[29401] = i[57];
  assign o[29402] = i[57];
  assign o[29403] = i[57];
  assign o[29404] = i[57];
  assign o[29405] = i[57];
  assign o[29406] = i[57];
  assign o[29407] = i[57];
  assign o[29408] = i[57];
  assign o[29409] = i[57];
  assign o[29410] = i[57];
  assign o[29411] = i[57];
  assign o[29412] = i[57];
  assign o[29413] = i[57];
  assign o[29414] = i[57];
  assign o[29415] = i[57];
  assign o[29416] = i[57];
  assign o[29417] = i[57];
  assign o[29418] = i[57];
  assign o[29419] = i[57];
  assign o[29420] = i[57];
  assign o[29421] = i[57];
  assign o[29422] = i[57];
  assign o[29423] = i[57];
  assign o[29424] = i[57];
  assign o[29425] = i[57];
  assign o[29426] = i[57];
  assign o[29427] = i[57];
  assign o[29428] = i[57];
  assign o[29429] = i[57];
  assign o[29430] = i[57];
  assign o[29431] = i[57];
  assign o[29432] = i[57];
  assign o[29433] = i[57];
  assign o[29434] = i[57];
  assign o[29435] = i[57];
  assign o[29436] = i[57];
  assign o[29437] = i[57];
  assign o[29438] = i[57];
  assign o[29439] = i[57];
  assign o[29440] = i[57];
  assign o[29441] = i[57];
  assign o[29442] = i[57];
  assign o[29443] = i[57];
  assign o[29444] = i[57];
  assign o[29445] = i[57];
  assign o[29446] = i[57];
  assign o[29447] = i[57];
  assign o[29448] = i[57];
  assign o[29449] = i[57];
  assign o[29450] = i[57];
  assign o[29451] = i[57];
  assign o[29452] = i[57];
  assign o[29453] = i[57];
  assign o[29454] = i[57];
  assign o[29455] = i[57];
  assign o[29456] = i[57];
  assign o[29457] = i[57];
  assign o[29458] = i[57];
  assign o[29459] = i[57];
  assign o[29460] = i[57];
  assign o[29461] = i[57];
  assign o[29462] = i[57];
  assign o[29463] = i[57];
  assign o[29464] = i[57];
  assign o[29465] = i[57];
  assign o[29466] = i[57];
  assign o[29467] = i[57];
  assign o[29468] = i[57];
  assign o[29469] = i[57];
  assign o[29470] = i[57];
  assign o[29471] = i[57];
  assign o[29472] = i[57];
  assign o[29473] = i[57];
  assign o[29474] = i[57];
  assign o[29475] = i[57];
  assign o[29476] = i[57];
  assign o[29477] = i[57];
  assign o[29478] = i[57];
  assign o[29479] = i[57];
  assign o[29480] = i[57];
  assign o[29481] = i[57];
  assign o[29482] = i[57];
  assign o[29483] = i[57];
  assign o[29484] = i[57];
  assign o[29485] = i[57];
  assign o[29486] = i[57];
  assign o[29487] = i[57];
  assign o[29488] = i[57];
  assign o[29489] = i[57];
  assign o[29490] = i[57];
  assign o[29491] = i[57];
  assign o[29492] = i[57];
  assign o[29493] = i[57];
  assign o[29494] = i[57];
  assign o[29495] = i[57];
  assign o[29496] = i[57];
  assign o[29497] = i[57];
  assign o[29498] = i[57];
  assign o[29499] = i[57];
  assign o[29500] = i[57];
  assign o[29501] = i[57];
  assign o[29502] = i[57];
  assign o[29503] = i[57];
  assign o[29504] = i[57];
  assign o[29505] = i[57];
  assign o[29506] = i[57];
  assign o[29507] = i[57];
  assign o[29508] = i[57];
  assign o[29509] = i[57];
  assign o[29510] = i[57];
  assign o[29511] = i[57];
  assign o[29512] = i[57];
  assign o[29513] = i[57];
  assign o[29514] = i[57];
  assign o[29515] = i[57];
  assign o[29516] = i[57];
  assign o[29517] = i[57];
  assign o[29518] = i[57];
  assign o[29519] = i[57];
  assign o[29520] = i[57];
  assign o[29521] = i[57];
  assign o[29522] = i[57];
  assign o[29523] = i[57];
  assign o[29524] = i[57];
  assign o[29525] = i[57];
  assign o[29526] = i[57];
  assign o[29527] = i[57];
  assign o[29528] = i[57];
  assign o[29529] = i[57];
  assign o[29530] = i[57];
  assign o[29531] = i[57];
  assign o[29532] = i[57];
  assign o[29533] = i[57];
  assign o[29534] = i[57];
  assign o[29535] = i[57];
  assign o[29536] = i[57];
  assign o[29537] = i[57];
  assign o[29538] = i[57];
  assign o[29539] = i[57];
  assign o[29540] = i[57];
  assign o[29541] = i[57];
  assign o[29542] = i[57];
  assign o[29543] = i[57];
  assign o[29544] = i[57];
  assign o[29545] = i[57];
  assign o[29546] = i[57];
  assign o[29547] = i[57];
  assign o[29548] = i[57];
  assign o[29549] = i[57];
  assign o[29550] = i[57];
  assign o[29551] = i[57];
  assign o[29552] = i[57];
  assign o[29553] = i[57];
  assign o[29554] = i[57];
  assign o[29555] = i[57];
  assign o[29556] = i[57];
  assign o[29557] = i[57];
  assign o[29558] = i[57];
  assign o[29559] = i[57];
  assign o[29560] = i[57];
  assign o[29561] = i[57];
  assign o[29562] = i[57];
  assign o[29563] = i[57];
  assign o[29564] = i[57];
  assign o[29565] = i[57];
  assign o[29566] = i[57];
  assign o[29567] = i[57];
  assign o[29568] = i[57];
  assign o[29569] = i[57];
  assign o[29570] = i[57];
  assign o[29571] = i[57];
  assign o[29572] = i[57];
  assign o[29573] = i[57];
  assign o[29574] = i[57];
  assign o[29575] = i[57];
  assign o[29576] = i[57];
  assign o[29577] = i[57];
  assign o[29578] = i[57];
  assign o[29579] = i[57];
  assign o[29580] = i[57];
  assign o[29581] = i[57];
  assign o[29582] = i[57];
  assign o[29583] = i[57];
  assign o[29584] = i[57];
  assign o[29585] = i[57];
  assign o[29586] = i[57];
  assign o[29587] = i[57];
  assign o[29588] = i[57];
  assign o[29589] = i[57];
  assign o[29590] = i[57];
  assign o[29591] = i[57];
  assign o[29592] = i[57];
  assign o[29593] = i[57];
  assign o[29594] = i[57];
  assign o[29595] = i[57];
  assign o[29596] = i[57];
  assign o[29597] = i[57];
  assign o[29598] = i[57];
  assign o[29599] = i[57];
  assign o[29600] = i[57];
  assign o[29601] = i[57];
  assign o[29602] = i[57];
  assign o[29603] = i[57];
  assign o[29604] = i[57];
  assign o[29605] = i[57];
  assign o[29606] = i[57];
  assign o[29607] = i[57];
  assign o[29608] = i[57];
  assign o[29609] = i[57];
  assign o[29610] = i[57];
  assign o[29611] = i[57];
  assign o[29612] = i[57];
  assign o[29613] = i[57];
  assign o[29614] = i[57];
  assign o[29615] = i[57];
  assign o[29616] = i[57];
  assign o[29617] = i[57];
  assign o[29618] = i[57];
  assign o[29619] = i[57];
  assign o[29620] = i[57];
  assign o[29621] = i[57];
  assign o[29622] = i[57];
  assign o[29623] = i[57];
  assign o[29624] = i[57];
  assign o[29625] = i[57];
  assign o[29626] = i[57];
  assign o[29627] = i[57];
  assign o[29628] = i[57];
  assign o[29629] = i[57];
  assign o[29630] = i[57];
  assign o[29631] = i[57];
  assign o[29632] = i[57];
  assign o[29633] = i[57];
  assign o[29634] = i[57];
  assign o[29635] = i[57];
  assign o[29636] = i[57];
  assign o[29637] = i[57];
  assign o[29638] = i[57];
  assign o[29639] = i[57];
  assign o[29640] = i[57];
  assign o[29641] = i[57];
  assign o[29642] = i[57];
  assign o[29643] = i[57];
  assign o[29644] = i[57];
  assign o[29645] = i[57];
  assign o[29646] = i[57];
  assign o[29647] = i[57];
  assign o[29648] = i[57];
  assign o[29649] = i[57];
  assign o[29650] = i[57];
  assign o[29651] = i[57];
  assign o[29652] = i[57];
  assign o[29653] = i[57];
  assign o[29654] = i[57];
  assign o[29655] = i[57];
  assign o[29656] = i[57];
  assign o[29657] = i[57];
  assign o[29658] = i[57];
  assign o[29659] = i[57];
  assign o[29660] = i[57];
  assign o[29661] = i[57];
  assign o[29662] = i[57];
  assign o[29663] = i[57];
  assign o[29664] = i[57];
  assign o[29665] = i[57];
  assign o[29666] = i[57];
  assign o[29667] = i[57];
  assign o[29668] = i[57];
  assign o[29669] = i[57];
  assign o[29670] = i[57];
  assign o[29671] = i[57];
  assign o[29672] = i[57];
  assign o[29673] = i[57];
  assign o[29674] = i[57];
  assign o[29675] = i[57];
  assign o[29676] = i[57];
  assign o[29677] = i[57];
  assign o[29678] = i[57];
  assign o[29679] = i[57];
  assign o[29680] = i[57];
  assign o[29681] = i[57];
  assign o[29682] = i[57];
  assign o[29683] = i[57];
  assign o[29684] = i[57];
  assign o[29685] = i[57];
  assign o[29686] = i[57];
  assign o[29687] = i[57];
  assign o[29688] = i[57];
  assign o[29689] = i[57];
  assign o[29690] = i[57];
  assign o[29691] = i[57];
  assign o[29692] = i[57];
  assign o[29693] = i[57];
  assign o[29694] = i[57];
  assign o[29695] = i[57];
  assign o[28672] = i[56];
  assign o[28673] = i[56];
  assign o[28674] = i[56];
  assign o[28675] = i[56];
  assign o[28676] = i[56];
  assign o[28677] = i[56];
  assign o[28678] = i[56];
  assign o[28679] = i[56];
  assign o[28680] = i[56];
  assign o[28681] = i[56];
  assign o[28682] = i[56];
  assign o[28683] = i[56];
  assign o[28684] = i[56];
  assign o[28685] = i[56];
  assign o[28686] = i[56];
  assign o[28687] = i[56];
  assign o[28688] = i[56];
  assign o[28689] = i[56];
  assign o[28690] = i[56];
  assign o[28691] = i[56];
  assign o[28692] = i[56];
  assign o[28693] = i[56];
  assign o[28694] = i[56];
  assign o[28695] = i[56];
  assign o[28696] = i[56];
  assign o[28697] = i[56];
  assign o[28698] = i[56];
  assign o[28699] = i[56];
  assign o[28700] = i[56];
  assign o[28701] = i[56];
  assign o[28702] = i[56];
  assign o[28703] = i[56];
  assign o[28704] = i[56];
  assign o[28705] = i[56];
  assign o[28706] = i[56];
  assign o[28707] = i[56];
  assign o[28708] = i[56];
  assign o[28709] = i[56];
  assign o[28710] = i[56];
  assign o[28711] = i[56];
  assign o[28712] = i[56];
  assign o[28713] = i[56];
  assign o[28714] = i[56];
  assign o[28715] = i[56];
  assign o[28716] = i[56];
  assign o[28717] = i[56];
  assign o[28718] = i[56];
  assign o[28719] = i[56];
  assign o[28720] = i[56];
  assign o[28721] = i[56];
  assign o[28722] = i[56];
  assign o[28723] = i[56];
  assign o[28724] = i[56];
  assign o[28725] = i[56];
  assign o[28726] = i[56];
  assign o[28727] = i[56];
  assign o[28728] = i[56];
  assign o[28729] = i[56];
  assign o[28730] = i[56];
  assign o[28731] = i[56];
  assign o[28732] = i[56];
  assign o[28733] = i[56];
  assign o[28734] = i[56];
  assign o[28735] = i[56];
  assign o[28736] = i[56];
  assign o[28737] = i[56];
  assign o[28738] = i[56];
  assign o[28739] = i[56];
  assign o[28740] = i[56];
  assign o[28741] = i[56];
  assign o[28742] = i[56];
  assign o[28743] = i[56];
  assign o[28744] = i[56];
  assign o[28745] = i[56];
  assign o[28746] = i[56];
  assign o[28747] = i[56];
  assign o[28748] = i[56];
  assign o[28749] = i[56];
  assign o[28750] = i[56];
  assign o[28751] = i[56];
  assign o[28752] = i[56];
  assign o[28753] = i[56];
  assign o[28754] = i[56];
  assign o[28755] = i[56];
  assign o[28756] = i[56];
  assign o[28757] = i[56];
  assign o[28758] = i[56];
  assign o[28759] = i[56];
  assign o[28760] = i[56];
  assign o[28761] = i[56];
  assign o[28762] = i[56];
  assign o[28763] = i[56];
  assign o[28764] = i[56];
  assign o[28765] = i[56];
  assign o[28766] = i[56];
  assign o[28767] = i[56];
  assign o[28768] = i[56];
  assign o[28769] = i[56];
  assign o[28770] = i[56];
  assign o[28771] = i[56];
  assign o[28772] = i[56];
  assign o[28773] = i[56];
  assign o[28774] = i[56];
  assign o[28775] = i[56];
  assign o[28776] = i[56];
  assign o[28777] = i[56];
  assign o[28778] = i[56];
  assign o[28779] = i[56];
  assign o[28780] = i[56];
  assign o[28781] = i[56];
  assign o[28782] = i[56];
  assign o[28783] = i[56];
  assign o[28784] = i[56];
  assign o[28785] = i[56];
  assign o[28786] = i[56];
  assign o[28787] = i[56];
  assign o[28788] = i[56];
  assign o[28789] = i[56];
  assign o[28790] = i[56];
  assign o[28791] = i[56];
  assign o[28792] = i[56];
  assign o[28793] = i[56];
  assign o[28794] = i[56];
  assign o[28795] = i[56];
  assign o[28796] = i[56];
  assign o[28797] = i[56];
  assign o[28798] = i[56];
  assign o[28799] = i[56];
  assign o[28800] = i[56];
  assign o[28801] = i[56];
  assign o[28802] = i[56];
  assign o[28803] = i[56];
  assign o[28804] = i[56];
  assign o[28805] = i[56];
  assign o[28806] = i[56];
  assign o[28807] = i[56];
  assign o[28808] = i[56];
  assign o[28809] = i[56];
  assign o[28810] = i[56];
  assign o[28811] = i[56];
  assign o[28812] = i[56];
  assign o[28813] = i[56];
  assign o[28814] = i[56];
  assign o[28815] = i[56];
  assign o[28816] = i[56];
  assign o[28817] = i[56];
  assign o[28818] = i[56];
  assign o[28819] = i[56];
  assign o[28820] = i[56];
  assign o[28821] = i[56];
  assign o[28822] = i[56];
  assign o[28823] = i[56];
  assign o[28824] = i[56];
  assign o[28825] = i[56];
  assign o[28826] = i[56];
  assign o[28827] = i[56];
  assign o[28828] = i[56];
  assign o[28829] = i[56];
  assign o[28830] = i[56];
  assign o[28831] = i[56];
  assign o[28832] = i[56];
  assign o[28833] = i[56];
  assign o[28834] = i[56];
  assign o[28835] = i[56];
  assign o[28836] = i[56];
  assign o[28837] = i[56];
  assign o[28838] = i[56];
  assign o[28839] = i[56];
  assign o[28840] = i[56];
  assign o[28841] = i[56];
  assign o[28842] = i[56];
  assign o[28843] = i[56];
  assign o[28844] = i[56];
  assign o[28845] = i[56];
  assign o[28846] = i[56];
  assign o[28847] = i[56];
  assign o[28848] = i[56];
  assign o[28849] = i[56];
  assign o[28850] = i[56];
  assign o[28851] = i[56];
  assign o[28852] = i[56];
  assign o[28853] = i[56];
  assign o[28854] = i[56];
  assign o[28855] = i[56];
  assign o[28856] = i[56];
  assign o[28857] = i[56];
  assign o[28858] = i[56];
  assign o[28859] = i[56];
  assign o[28860] = i[56];
  assign o[28861] = i[56];
  assign o[28862] = i[56];
  assign o[28863] = i[56];
  assign o[28864] = i[56];
  assign o[28865] = i[56];
  assign o[28866] = i[56];
  assign o[28867] = i[56];
  assign o[28868] = i[56];
  assign o[28869] = i[56];
  assign o[28870] = i[56];
  assign o[28871] = i[56];
  assign o[28872] = i[56];
  assign o[28873] = i[56];
  assign o[28874] = i[56];
  assign o[28875] = i[56];
  assign o[28876] = i[56];
  assign o[28877] = i[56];
  assign o[28878] = i[56];
  assign o[28879] = i[56];
  assign o[28880] = i[56];
  assign o[28881] = i[56];
  assign o[28882] = i[56];
  assign o[28883] = i[56];
  assign o[28884] = i[56];
  assign o[28885] = i[56];
  assign o[28886] = i[56];
  assign o[28887] = i[56];
  assign o[28888] = i[56];
  assign o[28889] = i[56];
  assign o[28890] = i[56];
  assign o[28891] = i[56];
  assign o[28892] = i[56];
  assign o[28893] = i[56];
  assign o[28894] = i[56];
  assign o[28895] = i[56];
  assign o[28896] = i[56];
  assign o[28897] = i[56];
  assign o[28898] = i[56];
  assign o[28899] = i[56];
  assign o[28900] = i[56];
  assign o[28901] = i[56];
  assign o[28902] = i[56];
  assign o[28903] = i[56];
  assign o[28904] = i[56];
  assign o[28905] = i[56];
  assign o[28906] = i[56];
  assign o[28907] = i[56];
  assign o[28908] = i[56];
  assign o[28909] = i[56];
  assign o[28910] = i[56];
  assign o[28911] = i[56];
  assign o[28912] = i[56];
  assign o[28913] = i[56];
  assign o[28914] = i[56];
  assign o[28915] = i[56];
  assign o[28916] = i[56];
  assign o[28917] = i[56];
  assign o[28918] = i[56];
  assign o[28919] = i[56];
  assign o[28920] = i[56];
  assign o[28921] = i[56];
  assign o[28922] = i[56];
  assign o[28923] = i[56];
  assign o[28924] = i[56];
  assign o[28925] = i[56];
  assign o[28926] = i[56];
  assign o[28927] = i[56];
  assign o[28928] = i[56];
  assign o[28929] = i[56];
  assign o[28930] = i[56];
  assign o[28931] = i[56];
  assign o[28932] = i[56];
  assign o[28933] = i[56];
  assign o[28934] = i[56];
  assign o[28935] = i[56];
  assign o[28936] = i[56];
  assign o[28937] = i[56];
  assign o[28938] = i[56];
  assign o[28939] = i[56];
  assign o[28940] = i[56];
  assign o[28941] = i[56];
  assign o[28942] = i[56];
  assign o[28943] = i[56];
  assign o[28944] = i[56];
  assign o[28945] = i[56];
  assign o[28946] = i[56];
  assign o[28947] = i[56];
  assign o[28948] = i[56];
  assign o[28949] = i[56];
  assign o[28950] = i[56];
  assign o[28951] = i[56];
  assign o[28952] = i[56];
  assign o[28953] = i[56];
  assign o[28954] = i[56];
  assign o[28955] = i[56];
  assign o[28956] = i[56];
  assign o[28957] = i[56];
  assign o[28958] = i[56];
  assign o[28959] = i[56];
  assign o[28960] = i[56];
  assign o[28961] = i[56];
  assign o[28962] = i[56];
  assign o[28963] = i[56];
  assign o[28964] = i[56];
  assign o[28965] = i[56];
  assign o[28966] = i[56];
  assign o[28967] = i[56];
  assign o[28968] = i[56];
  assign o[28969] = i[56];
  assign o[28970] = i[56];
  assign o[28971] = i[56];
  assign o[28972] = i[56];
  assign o[28973] = i[56];
  assign o[28974] = i[56];
  assign o[28975] = i[56];
  assign o[28976] = i[56];
  assign o[28977] = i[56];
  assign o[28978] = i[56];
  assign o[28979] = i[56];
  assign o[28980] = i[56];
  assign o[28981] = i[56];
  assign o[28982] = i[56];
  assign o[28983] = i[56];
  assign o[28984] = i[56];
  assign o[28985] = i[56];
  assign o[28986] = i[56];
  assign o[28987] = i[56];
  assign o[28988] = i[56];
  assign o[28989] = i[56];
  assign o[28990] = i[56];
  assign o[28991] = i[56];
  assign o[28992] = i[56];
  assign o[28993] = i[56];
  assign o[28994] = i[56];
  assign o[28995] = i[56];
  assign o[28996] = i[56];
  assign o[28997] = i[56];
  assign o[28998] = i[56];
  assign o[28999] = i[56];
  assign o[29000] = i[56];
  assign o[29001] = i[56];
  assign o[29002] = i[56];
  assign o[29003] = i[56];
  assign o[29004] = i[56];
  assign o[29005] = i[56];
  assign o[29006] = i[56];
  assign o[29007] = i[56];
  assign o[29008] = i[56];
  assign o[29009] = i[56];
  assign o[29010] = i[56];
  assign o[29011] = i[56];
  assign o[29012] = i[56];
  assign o[29013] = i[56];
  assign o[29014] = i[56];
  assign o[29015] = i[56];
  assign o[29016] = i[56];
  assign o[29017] = i[56];
  assign o[29018] = i[56];
  assign o[29019] = i[56];
  assign o[29020] = i[56];
  assign o[29021] = i[56];
  assign o[29022] = i[56];
  assign o[29023] = i[56];
  assign o[29024] = i[56];
  assign o[29025] = i[56];
  assign o[29026] = i[56];
  assign o[29027] = i[56];
  assign o[29028] = i[56];
  assign o[29029] = i[56];
  assign o[29030] = i[56];
  assign o[29031] = i[56];
  assign o[29032] = i[56];
  assign o[29033] = i[56];
  assign o[29034] = i[56];
  assign o[29035] = i[56];
  assign o[29036] = i[56];
  assign o[29037] = i[56];
  assign o[29038] = i[56];
  assign o[29039] = i[56];
  assign o[29040] = i[56];
  assign o[29041] = i[56];
  assign o[29042] = i[56];
  assign o[29043] = i[56];
  assign o[29044] = i[56];
  assign o[29045] = i[56];
  assign o[29046] = i[56];
  assign o[29047] = i[56];
  assign o[29048] = i[56];
  assign o[29049] = i[56];
  assign o[29050] = i[56];
  assign o[29051] = i[56];
  assign o[29052] = i[56];
  assign o[29053] = i[56];
  assign o[29054] = i[56];
  assign o[29055] = i[56];
  assign o[29056] = i[56];
  assign o[29057] = i[56];
  assign o[29058] = i[56];
  assign o[29059] = i[56];
  assign o[29060] = i[56];
  assign o[29061] = i[56];
  assign o[29062] = i[56];
  assign o[29063] = i[56];
  assign o[29064] = i[56];
  assign o[29065] = i[56];
  assign o[29066] = i[56];
  assign o[29067] = i[56];
  assign o[29068] = i[56];
  assign o[29069] = i[56];
  assign o[29070] = i[56];
  assign o[29071] = i[56];
  assign o[29072] = i[56];
  assign o[29073] = i[56];
  assign o[29074] = i[56];
  assign o[29075] = i[56];
  assign o[29076] = i[56];
  assign o[29077] = i[56];
  assign o[29078] = i[56];
  assign o[29079] = i[56];
  assign o[29080] = i[56];
  assign o[29081] = i[56];
  assign o[29082] = i[56];
  assign o[29083] = i[56];
  assign o[29084] = i[56];
  assign o[29085] = i[56];
  assign o[29086] = i[56];
  assign o[29087] = i[56];
  assign o[29088] = i[56];
  assign o[29089] = i[56];
  assign o[29090] = i[56];
  assign o[29091] = i[56];
  assign o[29092] = i[56];
  assign o[29093] = i[56];
  assign o[29094] = i[56];
  assign o[29095] = i[56];
  assign o[29096] = i[56];
  assign o[29097] = i[56];
  assign o[29098] = i[56];
  assign o[29099] = i[56];
  assign o[29100] = i[56];
  assign o[29101] = i[56];
  assign o[29102] = i[56];
  assign o[29103] = i[56];
  assign o[29104] = i[56];
  assign o[29105] = i[56];
  assign o[29106] = i[56];
  assign o[29107] = i[56];
  assign o[29108] = i[56];
  assign o[29109] = i[56];
  assign o[29110] = i[56];
  assign o[29111] = i[56];
  assign o[29112] = i[56];
  assign o[29113] = i[56];
  assign o[29114] = i[56];
  assign o[29115] = i[56];
  assign o[29116] = i[56];
  assign o[29117] = i[56];
  assign o[29118] = i[56];
  assign o[29119] = i[56];
  assign o[29120] = i[56];
  assign o[29121] = i[56];
  assign o[29122] = i[56];
  assign o[29123] = i[56];
  assign o[29124] = i[56];
  assign o[29125] = i[56];
  assign o[29126] = i[56];
  assign o[29127] = i[56];
  assign o[29128] = i[56];
  assign o[29129] = i[56];
  assign o[29130] = i[56];
  assign o[29131] = i[56];
  assign o[29132] = i[56];
  assign o[29133] = i[56];
  assign o[29134] = i[56];
  assign o[29135] = i[56];
  assign o[29136] = i[56];
  assign o[29137] = i[56];
  assign o[29138] = i[56];
  assign o[29139] = i[56];
  assign o[29140] = i[56];
  assign o[29141] = i[56];
  assign o[29142] = i[56];
  assign o[29143] = i[56];
  assign o[29144] = i[56];
  assign o[29145] = i[56];
  assign o[29146] = i[56];
  assign o[29147] = i[56];
  assign o[29148] = i[56];
  assign o[29149] = i[56];
  assign o[29150] = i[56];
  assign o[29151] = i[56];
  assign o[29152] = i[56];
  assign o[29153] = i[56];
  assign o[29154] = i[56];
  assign o[29155] = i[56];
  assign o[29156] = i[56];
  assign o[29157] = i[56];
  assign o[29158] = i[56];
  assign o[29159] = i[56];
  assign o[29160] = i[56];
  assign o[29161] = i[56];
  assign o[29162] = i[56];
  assign o[29163] = i[56];
  assign o[29164] = i[56];
  assign o[29165] = i[56];
  assign o[29166] = i[56];
  assign o[29167] = i[56];
  assign o[29168] = i[56];
  assign o[29169] = i[56];
  assign o[29170] = i[56];
  assign o[29171] = i[56];
  assign o[29172] = i[56];
  assign o[29173] = i[56];
  assign o[29174] = i[56];
  assign o[29175] = i[56];
  assign o[29176] = i[56];
  assign o[29177] = i[56];
  assign o[29178] = i[56];
  assign o[29179] = i[56];
  assign o[29180] = i[56];
  assign o[29181] = i[56];
  assign o[29182] = i[56];
  assign o[29183] = i[56];
  assign o[28160] = i[55];
  assign o[28161] = i[55];
  assign o[28162] = i[55];
  assign o[28163] = i[55];
  assign o[28164] = i[55];
  assign o[28165] = i[55];
  assign o[28166] = i[55];
  assign o[28167] = i[55];
  assign o[28168] = i[55];
  assign o[28169] = i[55];
  assign o[28170] = i[55];
  assign o[28171] = i[55];
  assign o[28172] = i[55];
  assign o[28173] = i[55];
  assign o[28174] = i[55];
  assign o[28175] = i[55];
  assign o[28176] = i[55];
  assign o[28177] = i[55];
  assign o[28178] = i[55];
  assign o[28179] = i[55];
  assign o[28180] = i[55];
  assign o[28181] = i[55];
  assign o[28182] = i[55];
  assign o[28183] = i[55];
  assign o[28184] = i[55];
  assign o[28185] = i[55];
  assign o[28186] = i[55];
  assign o[28187] = i[55];
  assign o[28188] = i[55];
  assign o[28189] = i[55];
  assign o[28190] = i[55];
  assign o[28191] = i[55];
  assign o[28192] = i[55];
  assign o[28193] = i[55];
  assign o[28194] = i[55];
  assign o[28195] = i[55];
  assign o[28196] = i[55];
  assign o[28197] = i[55];
  assign o[28198] = i[55];
  assign o[28199] = i[55];
  assign o[28200] = i[55];
  assign o[28201] = i[55];
  assign o[28202] = i[55];
  assign o[28203] = i[55];
  assign o[28204] = i[55];
  assign o[28205] = i[55];
  assign o[28206] = i[55];
  assign o[28207] = i[55];
  assign o[28208] = i[55];
  assign o[28209] = i[55];
  assign o[28210] = i[55];
  assign o[28211] = i[55];
  assign o[28212] = i[55];
  assign o[28213] = i[55];
  assign o[28214] = i[55];
  assign o[28215] = i[55];
  assign o[28216] = i[55];
  assign o[28217] = i[55];
  assign o[28218] = i[55];
  assign o[28219] = i[55];
  assign o[28220] = i[55];
  assign o[28221] = i[55];
  assign o[28222] = i[55];
  assign o[28223] = i[55];
  assign o[28224] = i[55];
  assign o[28225] = i[55];
  assign o[28226] = i[55];
  assign o[28227] = i[55];
  assign o[28228] = i[55];
  assign o[28229] = i[55];
  assign o[28230] = i[55];
  assign o[28231] = i[55];
  assign o[28232] = i[55];
  assign o[28233] = i[55];
  assign o[28234] = i[55];
  assign o[28235] = i[55];
  assign o[28236] = i[55];
  assign o[28237] = i[55];
  assign o[28238] = i[55];
  assign o[28239] = i[55];
  assign o[28240] = i[55];
  assign o[28241] = i[55];
  assign o[28242] = i[55];
  assign o[28243] = i[55];
  assign o[28244] = i[55];
  assign o[28245] = i[55];
  assign o[28246] = i[55];
  assign o[28247] = i[55];
  assign o[28248] = i[55];
  assign o[28249] = i[55];
  assign o[28250] = i[55];
  assign o[28251] = i[55];
  assign o[28252] = i[55];
  assign o[28253] = i[55];
  assign o[28254] = i[55];
  assign o[28255] = i[55];
  assign o[28256] = i[55];
  assign o[28257] = i[55];
  assign o[28258] = i[55];
  assign o[28259] = i[55];
  assign o[28260] = i[55];
  assign o[28261] = i[55];
  assign o[28262] = i[55];
  assign o[28263] = i[55];
  assign o[28264] = i[55];
  assign o[28265] = i[55];
  assign o[28266] = i[55];
  assign o[28267] = i[55];
  assign o[28268] = i[55];
  assign o[28269] = i[55];
  assign o[28270] = i[55];
  assign o[28271] = i[55];
  assign o[28272] = i[55];
  assign o[28273] = i[55];
  assign o[28274] = i[55];
  assign o[28275] = i[55];
  assign o[28276] = i[55];
  assign o[28277] = i[55];
  assign o[28278] = i[55];
  assign o[28279] = i[55];
  assign o[28280] = i[55];
  assign o[28281] = i[55];
  assign o[28282] = i[55];
  assign o[28283] = i[55];
  assign o[28284] = i[55];
  assign o[28285] = i[55];
  assign o[28286] = i[55];
  assign o[28287] = i[55];
  assign o[28288] = i[55];
  assign o[28289] = i[55];
  assign o[28290] = i[55];
  assign o[28291] = i[55];
  assign o[28292] = i[55];
  assign o[28293] = i[55];
  assign o[28294] = i[55];
  assign o[28295] = i[55];
  assign o[28296] = i[55];
  assign o[28297] = i[55];
  assign o[28298] = i[55];
  assign o[28299] = i[55];
  assign o[28300] = i[55];
  assign o[28301] = i[55];
  assign o[28302] = i[55];
  assign o[28303] = i[55];
  assign o[28304] = i[55];
  assign o[28305] = i[55];
  assign o[28306] = i[55];
  assign o[28307] = i[55];
  assign o[28308] = i[55];
  assign o[28309] = i[55];
  assign o[28310] = i[55];
  assign o[28311] = i[55];
  assign o[28312] = i[55];
  assign o[28313] = i[55];
  assign o[28314] = i[55];
  assign o[28315] = i[55];
  assign o[28316] = i[55];
  assign o[28317] = i[55];
  assign o[28318] = i[55];
  assign o[28319] = i[55];
  assign o[28320] = i[55];
  assign o[28321] = i[55];
  assign o[28322] = i[55];
  assign o[28323] = i[55];
  assign o[28324] = i[55];
  assign o[28325] = i[55];
  assign o[28326] = i[55];
  assign o[28327] = i[55];
  assign o[28328] = i[55];
  assign o[28329] = i[55];
  assign o[28330] = i[55];
  assign o[28331] = i[55];
  assign o[28332] = i[55];
  assign o[28333] = i[55];
  assign o[28334] = i[55];
  assign o[28335] = i[55];
  assign o[28336] = i[55];
  assign o[28337] = i[55];
  assign o[28338] = i[55];
  assign o[28339] = i[55];
  assign o[28340] = i[55];
  assign o[28341] = i[55];
  assign o[28342] = i[55];
  assign o[28343] = i[55];
  assign o[28344] = i[55];
  assign o[28345] = i[55];
  assign o[28346] = i[55];
  assign o[28347] = i[55];
  assign o[28348] = i[55];
  assign o[28349] = i[55];
  assign o[28350] = i[55];
  assign o[28351] = i[55];
  assign o[28352] = i[55];
  assign o[28353] = i[55];
  assign o[28354] = i[55];
  assign o[28355] = i[55];
  assign o[28356] = i[55];
  assign o[28357] = i[55];
  assign o[28358] = i[55];
  assign o[28359] = i[55];
  assign o[28360] = i[55];
  assign o[28361] = i[55];
  assign o[28362] = i[55];
  assign o[28363] = i[55];
  assign o[28364] = i[55];
  assign o[28365] = i[55];
  assign o[28366] = i[55];
  assign o[28367] = i[55];
  assign o[28368] = i[55];
  assign o[28369] = i[55];
  assign o[28370] = i[55];
  assign o[28371] = i[55];
  assign o[28372] = i[55];
  assign o[28373] = i[55];
  assign o[28374] = i[55];
  assign o[28375] = i[55];
  assign o[28376] = i[55];
  assign o[28377] = i[55];
  assign o[28378] = i[55];
  assign o[28379] = i[55];
  assign o[28380] = i[55];
  assign o[28381] = i[55];
  assign o[28382] = i[55];
  assign o[28383] = i[55];
  assign o[28384] = i[55];
  assign o[28385] = i[55];
  assign o[28386] = i[55];
  assign o[28387] = i[55];
  assign o[28388] = i[55];
  assign o[28389] = i[55];
  assign o[28390] = i[55];
  assign o[28391] = i[55];
  assign o[28392] = i[55];
  assign o[28393] = i[55];
  assign o[28394] = i[55];
  assign o[28395] = i[55];
  assign o[28396] = i[55];
  assign o[28397] = i[55];
  assign o[28398] = i[55];
  assign o[28399] = i[55];
  assign o[28400] = i[55];
  assign o[28401] = i[55];
  assign o[28402] = i[55];
  assign o[28403] = i[55];
  assign o[28404] = i[55];
  assign o[28405] = i[55];
  assign o[28406] = i[55];
  assign o[28407] = i[55];
  assign o[28408] = i[55];
  assign o[28409] = i[55];
  assign o[28410] = i[55];
  assign o[28411] = i[55];
  assign o[28412] = i[55];
  assign o[28413] = i[55];
  assign o[28414] = i[55];
  assign o[28415] = i[55];
  assign o[28416] = i[55];
  assign o[28417] = i[55];
  assign o[28418] = i[55];
  assign o[28419] = i[55];
  assign o[28420] = i[55];
  assign o[28421] = i[55];
  assign o[28422] = i[55];
  assign o[28423] = i[55];
  assign o[28424] = i[55];
  assign o[28425] = i[55];
  assign o[28426] = i[55];
  assign o[28427] = i[55];
  assign o[28428] = i[55];
  assign o[28429] = i[55];
  assign o[28430] = i[55];
  assign o[28431] = i[55];
  assign o[28432] = i[55];
  assign o[28433] = i[55];
  assign o[28434] = i[55];
  assign o[28435] = i[55];
  assign o[28436] = i[55];
  assign o[28437] = i[55];
  assign o[28438] = i[55];
  assign o[28439] = i[55];
  assign o[28440] = i[55];
  assign o[28441] = i[55];
  assign o[28442] = i[55];
  assign o[28443] = i[55];
  assign o[28444] = i[55];
  assign o[28445] = i[55];
  assign o[28446] = i[55];
  assign o[28447] = i[55];
  assign o[28448] = i[55];
  assign o[28449] = i[55];
  assign o[28450] = i[55];
  assign o[28451] = i[55];
  assign o[28452] = i[55];
  assign o[28453] = i[55];
  assign o[28454] = i[55];
  assign o[28455] = i[55];
  assign o[28456] = i[55];
  assign o[28457] = i[55];
  assign o[28458] = i[55];
  assign o[28459] = i[55];
  assign o[28460] = i[55];
  assign o[28461] = i[55];
  assign o[28462] = i[55];
  assign o[28463] = i[55];
  assign o[28464] = i[55];
  assign o[28465] = i[55];
  assign o[28466] = i[55];
  assign o[28467] = i[55];
  assign o[28468] = i[55];
  assign o[28469] = i[55];
  assign o[28470] = i[55];
  assign o[28471] = i[55];
  assign o[28472] = i[55];
  assign o[28473] = i[55];
  assign o[28474] = i[55];
  assign o[28475] = i[55];
  assign o[28476] = i[55];
  assign o[28477] = i[55];
  assign o[28478] = i[55];
  assign o[28479] = i[55];
  assign o[28480] = i[55];
  assign o[28481] = i[55];
  assign o[28482] = i[55];
  assign o[28483] = i[55];
  assign o[28484] = i[55];
  assign o[28485] = i[55];
  assign o[28486] = i[55];
  assign o[28487] = i[55];
  assign o[28488] = i[55];
  assign o[28489] = i[55];
  assign o[28490] = i[55];
  assign o[28491] = i[55];
  assign o[28492] = i[55];
  assign o[28493] = i[55];
  assign o[28494] = i[55];
  assign o[28495] = i[55];
  assign o[28496] = i[55];
  assign o[28497] = i[55];
  assign o[28498] = i[55];
  assign o[28499] = i[55];
  assign o[28500] = i[55];
  assign o[28501] = i[55];
  assign o[28502] = i[55];
  assign o[28503] = i[55];
  assign o[28504] = i[55];
  assign o[28505] = i[55];
  assign o[28506] = i[55];
  assign o[28507] = i[55];
  assign o[28508] = i[55];
  assign o[28509] = i[55];
  assign o[28510] = i[55];
  assign o[28511] = i[55];
  assign o[28512] = i[55];
  assign o[28513] = i[55];
  assign o[28514] = i[55];
  assign o[28515] = i[55];
  assign o[28516] = i[55];
  assign o[28517] = i[55];
  assign o[28518] = i[55];
  assign o[28519] = i[55];
  assign o[28520] = i[55];
  assign o[28521] = i[55];
  assign o[28522] = i[55];
  assign o[28523] = i[55];
  assign o[28524] = i[55];
  assign o[28525] = i[55];
  assign o[28526] = i[55];
  assign o[28527] = i[55];
  assign o[28528] = i[55];
  assign o[28529] = i[55];
  assign o[28530] = i[55];
  assign o[28531] = i[55];
  assign o[28532] = i[55];
  assign o[28533] = i[55];
  assign o[28534] = i[55];
  assign o[28535] = i[55];
  assign o[28536] = i[55];
  assign o[28537] = i[55];
  assign o[28538] = i[55];
  assign o[28539] = i[55];
  assign o[28540] = i[55];
  assign o[28541] = i[55];
  assign o[28542] = i[55];
  assign o[28543] = i[55];
  assign o[28544] = i[55];
  assign o[28545] = i[55];
  assign o[28546] = i[55];
  assign o[28547] = i[55];
  assign o[28548] = i[55];
  assign o[28549] = i[55];
  assign o[28550] = i[55];
  assign o[28551] = i[55];
  assign o[28552] = i[55];
  assign o[28553] = i[55];
  assign o[28554] = i[55];
  assign o[28555] = i[55];
  assign o[28556] = i[55];
  assign o[28557] = i[55];
  assign o[28558] = i[55];
  assign o[28559] = i[55];
  assign o[28560] = i[55];
  assign o[28561] = i[55];
  assign o[28562] = i[55];
  assign o[28563] = i[55];
  assign o[28564] = i[55];
  assign o[28565] = i[55];
  assign o[28566] = i[55];
  assign o[28567] = i[55];
  assign o[28568] = i[55];
  assign o[28569] = i[55];
  assign o[28570] = i[55];
  assign o[28571] = i[55];
  assign o[28572] = i[55];
  assign o[28573] = i[55];
  assign o[28574] = i[55];
  assign o[28575] = i[55];
  assign o[28576] = i[55];
  assign o[28577] = i[55];
  assign o[28578] = i[55];
  assign o[28579] = i[55];
  assign o[28580] = i[55];
  assign o[28581] = i[55];
  assign o[28582] = i[55];
  assign o[28583] = i[55];
  assign o[28584] = i[55];
  assign o[28585] = i[55];
  assign o[28586] = i[55];
  assign o[28587] = i[55];
  assign o[28588] = i[55];
  assign o[28589] = i[55];
  assign o[28590] = i[55];
  assign o[28591] = i[55];
  assign o[28592] = i[55];
  assign o[28593] = i[55];
  assign o[28594] = i[55];
  assign o[28595] = i[55];
  assign o[28596] = i[55];
  assign o[28597] = i[55];
  assign o[28598] = i[55];
  assign o[28599] = i[55];
  assign o[28600] = i[55];
  assign o[28601] = i[55];
  assign o[28602] = i[55];
  assign o[28603] = i[55];
  assign o[28604] = i[55];
  assign o[28605] = i[55];
  assign o[28606] = i[55];
  assign o[28607] = i[55];
  assign o[28608] = i[55];
  assign o[28609] = i[55];
  assign o[28610] = i[55];
  assign o[28611] = i[55];
  assign o[28612] = i[55];
  assign o[28613] = i[55];
  assign o[28614] = i[55];
  assign o[28615] = i[55];
  assign o[28616] = i[55];
  assign o[28617] = i[55];
  assign o[28618] = i[55];
  assign o[28619] = i[55];
  assign o[28620] = i[55];
  assign o[28621] = i[55];
  assign o[28622] = i[55];
  assign o[28623] = i[55];
  assign o[28624] = i[55];
  assign o[28625] = i[55];
  assign o[28626] = i[55];
  assign o[28627] = i[55];
  assign o[28628] = i[55];
  assign o[28629] = i[55];
  assign o[28630] = i[55];
  assign o[28631] = i[55];
  assign o[28632] = i[55];
  assign o[28633] = i[55];
  assign o[28634] = i[55];
  assign o[28635] = i[55];
  assign o[28636] = i[55];
  assign o[28637] = i[55];
  assign o[28638] = i[55];
  assign o[28639] = i[55];
  assign o[28640] = i[55];
  assign o[28641] = i[55];
  assign o[28642] = i[55];
  assign o[28643] = i[55];
  assign o[28644] = i[55];
  assign o[28645] = i[55];
  assign o[28646] = i[55];
  assign o[28647] = i[55];
  assign o[28648] = i[55];
  assign o[28649] = i[55];
  assign o[28650] = i[55];
  assign o[28651] = i[55];
  assign o[28652] = i[55];
  assign o[28653] = i[55];
  assign o[28654] = i[55];
  assign o[28655] = i[55];
  assign o[28656] = i[55];
  assign o[28657] = i[55];
  assign o[28658] = i[55];
  assign o[28659] = i[55];
  assign o[28660] = i[55];
  assign o[28661] = i[55];
  assign o[28662] = i[55];
  assign o[28663] = i[55];
  assign o[28664] = i[55];
  assign o[28665] = i[55];
  assign o[28666] = i[55];
  assign o[28667] = i[55];
  assign o[28668] = i[55];
  assign o[28669] = i[55];
  assign o[28670] = i[55];
  assign o[28671] = i[55];
  assign o[27648] = i[54];
  assign o[27649] = i[54];
  assign o[27650] = i[54];
  assign o[27651] = i[54];
  assign o[27652] = i[54];
  assign o[27653] = i[54];
  assign o[27654] = i[54];
  assign o[27655] = i[54];
  assign o[27656] = i[54];
  assign o[27657] = i[54];
  assign o[27658] = i[54];
  assign o[27659] = i[54];
  assign o[27660] = i[54];
  assign o[27661] = i[54];
  assign o[27662] = i[54];
  assign o[27663] = i[54];
  assign o[27664] = i[54];
  assign o[27665] = i[54];
  assign o[27666] = i[54];
  assign o[27667] = i[54];
  assign o[27668] = i[54];
  assign o[27669] = i[54];
  assign o[27670] = i[54];
  assign o[27671] = i[54];
  assign o[27672] = i[54];
  assign o[27673] = i[54];
  assign o[27674] = i[54];
  assign o[27675] = i[54];
  assign o[27676] = i[54];
  assign o[27677] = i[54];
  assign o[27678] = i[54];
  assign o[27679] = i[54];
  assign o[27680] = i[54];
  assign o[27681] = i[54];
  assign o[27682] = i[54];
  assign o[27683] = i[54];
  assign o[27684] = i[54];
  assign o[27685] = i[54];
  assign o[27686] = i[54];
  assign o[27687] = i[54];
  assign o[27688] = i[54];
  assign o[27689] = i[54];
  assign o[27690] = i[54];
  assign o[27691] = i[54];
  assign o[27692] = i[54];
  assign o[27693] = i[54];
  assign o[27694] = i[54];
  assign o[27695] = i[54];
  assign o[27696] = i[54];
  assign o[27697] = i[54];
  assign o[27698] = i[54];
  assign o[27699] = i[54];
  assign o[27700] = i[54];
  assign o[27701] = i[54];
  assign o[27702] = i[54];
  assign o[27703] = i[54];
  assign o[27704] = i[54];
  assign o[27705] = i[54];
  assign o[27706] = i[54];
  assign o[27707] = i[54];
  assign o[27708] = i[54];
  assign o[27709] = i[54];
  assign o[27710] = i[54];
  assign o[27711] = i[54];
  assign o[27712] = i[54];
  assign o[27713] = i[54];
  assign o[27714] = i[54];
  assign o[27715] = i[54];
  assign o[27716] = i[54];
  assign o[27717] = i[54];
  assign o[27718] = i[54];
  assign o[27719] = i[54];
  assign o[27720] = i[54];
  assign o[27721] = i[54];
  assign o[27722] = i[54];
  assign o[27723] = i[54];
  assign o[27724] = i[54];
  assign o[27725] = i[54];
  assign o[27726] = i[54];
  assign o[27727] = i[54];
  assign o[27728] = i[54];
  assign o[27729] = i[54];
  assign o[27730] = i[54];
  assign o[27731] = i[54];
  assign o[27732] = i[54];
  assign o[27733] = i[54];
  assign o[27734] = i[54];
  assign o[27735] = i[54];
  assign o[27736] = i[54];
  assign o[27737] = i[54];
  assign o[27738] = i[54];
  assign o[27739] = i[54];
  assign o[27740] = i[54];
  assign o[27741] = i[54];
  assign o[27742] = i[54];
  assign o[27743] = i[54];
  assign o[27744] = i[54];
  assign o[27745] = i[54];
  assign o[27746] = i[54];
  assign o[27747] = i[54];
  assign o[27748] = i[54];
  assign o[27749] = i[54];
  assign o[27750] = i[54];
  assign o[27751] = i[54];
  assign o[27752] = i[54];
  assign o[27753] = i[54];
  assign o[27754] = i[54];
  assign o[27755] = i[54];
  assign o[27756] = i[54];
  assign o[27757] = i[54];
  assign o[27758] = i[54];
  assign o[27759] = i[54];
  assign o[27760] = i[54];
  assign o[27761] = i[54];
  assign o[27762] = i[54];
  assign o[27763] = i[54];
  assign o[27764] = i[54];
  assign o[27765] = i[54];
  assign o[27766] = i[54];
  assign o[27767] = i[54];
  assign o[27768] = i[54];
  assign o[27769] = i[54];
  assign o[27770] = i[54];
  assign o[27771] = i[54];
  assign o[27772] = i[54];
  assign o[27773] = i[54];
  assign o[27774] = i[54];
  assign o[27775] = i[54];
  assign o[27776] = i[54];
  assign o[27777] = i[54];
  assign o[27778] = i[54];
  assign o[27779] = i[54];
  assign o[27780] = i[54];
  assign o[27781] = i[54];
  assign o[27782] = i[54];
  assign o[27783] = i[54];
  assign o[27784] = i[54];
  assign o[27785] = i[54];
  assign o[27786] = i[54];
  assign o[27787] = i[54];
  assign o[27788] = i[54];
  assign o[27789] = i[54];
  assign o[27790] = i[54];
  assign o[27791] = i[54];
  assign o[27792] = i[54];
  assign o[27793] = i[54];
  assign o[27794] = i[54];
  assign o[27795] = i[54];
  assign o[27796] = i[54];
  assign o[27797] = i[54];
  assign o[27798] = i[54];
  assign o[27799] = i[54];
  assign o[27800] = i[54];
  assign o[27801] = i[54];
  assign o[27802] = i[54];
  assign o[27803] = i[54];
  assign o[27804] = i[54];
  assign o[27805] = i[54];
  assign o[27806] = i[54];
  assign o[27807] = i[54];
  assign o[27808] = i[54];
  assign o[27809] = i[54];
  assign o[27810] = i[54];
  assign o[27811] = i[54];
  assign o[27812] = i[54];
  assign o[27813] = i[54];
  assign o[27814] = i[54];
  assign o[27815] = i[54];
  assign o[27816] = i[54];
  assign o[27817] = i[54];
  assign o[27818] = i[54];
  assign o[27819] = i[54];
  assign o[27820] = i[54];
  assign o[27821] = i[54];
  assign o[27822] = i[54];
  assign o[27823] = i[54];
  assign o[27824] = i[54];
  assign o[27825] = i[54];
  assign o[27826] = i[54];
  assign o[27827] = i[54];
  assign o[27828] = i[54];
  assign o[27829] = i[54];
  assign o[27830] = i[54];
  assign o[27831] = i[54];
  assign o[27832] = i[54];
  assign o[27833] = i[54];
  assign o[27834] = i[54];
  assign o[27835] = i[54];
  assign o[27836] = i[54];
  assign o[27837] = i[54];
  assign o[27838] = i[54];
  assign o[27839] = i[54];
  assign o[27840] = i[54];
  assign o[27841] = i[54];
  assign o[27842] = i[54];
  assign o[27843] = i[54];
  assign o[27844] = i[54];
  assign o[27845] = i[54];
  assign o[27846] = i[54];
  assign o[27847] = i[54];
  assign o[27848] = i[54];
  assign o[27849] = i[54];
  assign o[27850] = i[54];
  assign o[27851] = i[54];
  assign o[27852] = i[54];
  assign o[27853] = i[54];
  assign o[27854] = i[54];
  assign o[27855] = i[54];
  assign o[27856] = i[54];
  assign o[27857] = i[54];
  assign o[27858] = i[54];
  assign o[27859] = i[54];
  assign o[27860] = i[54];
  assign o[27861] = i[54];
  assign o[27862] = i[54];
  assign o[27863] = i[54];
  assign o[27864] = i[54];
  assign o[27865] = i[54];
  assign o[27866] = i[54];
  assign o[27867] = i[54];
  assign o[27868] = i[54];
  assign o[27869] = i[54];
  assign o[27870] = i[54];
  assign o[27871] = i[54];
  assign o[27872] = i[54];
  assign o[27873] = i[54];
  assign o[27874] = i[54];
  assign o[27875] = i[54];
  assign o[27876] = i[54];
  assign o[27877] = i[54];
  assign o[27878] = i[54];
  assign o[27879] = i[54];
  assign o[27880] = i[54];
  assign o[27881] = i[54];
  assign o[27882] = i[54];
  assign o[27883] = i[54];
  assign o[27884] = i[54];
  assign o[27885] = i[54];
  assign o[27886] = i[54];
  assign o[27887] = i[54];
  assign o[27888] = i[54];
  assign o[27889] = i[54];
  assign o[27890] = i[54];
  assign o[27891] = i[54];
  assign o[27892] = i[54];
  assign o[27893] = i[54];
  assign o[27894] = i[54];
  assign o[27895] = i[54];
  assign o[27896] = i[54];
  assign o[27897] = i[54];
  assign o[27898] = i[54];
  assign o[27899] = i[54];
  assign o[27900] = i[54];
  assign o[27901] = i[54];
  assign o[27902] = i[54];
  assign o[27903] = i[54];
  assign o[27904] = i[54];
  assign o[27905] = i[54];
  assign o[27906] = i[54];
  assign o[27907] = i[54];
  assign o[27908] = i[54];
  assign o[27909] = i[54];
  assign o[27910] = i[54];
  assign o[27911] = i[54];
  assign o[27912] = i[54];
  assign o[27913] = i[54];
  assign o[27914] = i[54];
  assign o[27915] = i[54];
  assign o[27916] = i[54];
  assign o[27917] = i[54];
  assign o[27918] = i[54];
  assign o[27919] = i[54];
  assign o[27920] = i[54];
  assign o[27921] = i[54];
  assign o[27922] = i[54];
  assign o[27923] = i[54];
  assign o[27924] = i[54];
  assign o[27925] = i[54];
  assign o[27926] = i[54];
  assign o[27927] = i[54];
  assign o[27928] = i[54];
  assign o[27929] = i[54];
  assign o[27930] = i[54];
  assign o[27931] = i[54];
  assign o[27932] = i[54];
  assign o[27933] = i[54];
  assign o[27934] = i[54];
  assign o[27935] = i[54];
  assign o[27936] = i[54];
  assign o[27937] = i[54];
  assign o[27938] = i[54];
  assign o[27939] = i[54];
  assign o[27940] = i[54];
  assign o[27941] = i[54];
  assign o[27942] = i[54];
  assign o[27943] = i[54];
  assign o[27944] = i[54];
  assign o[27945] = i[54];
  assign o[27946] = i[54];
  assign o[27947] = i[54];
  assign o[27948] = i[54];
  assign o[27949] = i[54];
  assign o[27950] = i[54];
  assign o[27951] = i[54];
  assign o[27952] = i[54];
  assign o[27953] = i[54];
  assign o[27954] = i[54];
  assign o[27955] = i[54];
  assign o[27956] = i[54];
  assign o[27957] = i[54];
  assign o[27958] = i[54];
  assign o[27959] = i[54];
  assign o[27960] = i[54];
  assign o[27961] = i[54];
  assign o[27962] = i[54];
  assign o[27963] = i[54];
  assign o[27964] = i[54];
  assign o[27965] = i[54];
  assign o[27966] = i[54];
  assign o[27967] = i[54];
  assign o[27968] = i[54];
  assign o[27969] = i[54];
  assign o[27970] = i[54];
  assign o[27971] = i[54];
  assign o[27972] = i[54];
  assign o[27973] = i[54];
  assign o[27974] = i[54];
  assign o[27975] = i[54];
  assign o[27976] = i[54];
  assign o[27977] = i[54];
  assign o[27978] = i[54];
  assign o[27979] = i[54];
  assign o[27980] = i[54];
  assign o[27981] = i[54];
  assign o[27982] = i[54];
  assign o[27983] = i[54];
  assign o[27984] = i[54];
  assign o[27985] = i[54];
  assign o[27986] = i[54];
  assign o[27987] = i[54];
  assign o[27988] = i[54];
  assign o[27989] = i[54];
  assign o[27990] = i[54];
  assign o[27991] = i[54];
  assign o[27992] = i[54];
  assign o[27993] = i[54];
  assign o[27994] = i[54];
  assign o[27995] = i[54];
  assign o[27996] = i[54];
  assign o[27997] = i[54];
  assign o[27998] = i[54];
  assign o[27999] = i[54];
  assign o[28000] = i[54];
  assign o[28001] = i[54];
  assign o[28002] = i[54];
  assign o[28003] = i[54];
  assign o[28004] = i[54];
  assign o[28005] = i[54];
  assign o[28006] = i[54];
  assign o[28007] = i[54];
  assign o[28008] = i[54];
  assign o[28009] = i[54];
  assign o[28010] = i[54];
  assign o[28011] = i[54];
  assign o[28012] = i[54];
  assign o[28013] = i[54];
  assign o[28014] = i[54];
  assign o[28015] = i[54];
  assign o[28016] = i[54];
  assign o[28017] = i[54];
  assign o[28018] = i[54];
  assign o[28019] = i[54];
  assign o[28020] = i[54];
  assign o[28021] = i[54];
  assign o[28022] = i[54];
  assign o[28023] = i[54];
  assign o[28024] = i[54];
  assign o[28025] = i[54];
  assign o[28026] = i[54];
  assign o[28027] = i[54];
  assign o[28028] = i[54];
  assign o[28029] = i[54];
  assign o[28030] = i[54];
  assign o[28031] = i[54];
  assign o[28032] = i[54];
  assign o[28033] = i[54];
  assign o[28034] = i[54];
  assign o[28035] = i[54];
  assign o[28036] = i[54];
  assign o[28037] = i[54];
  assign o[28038] = i[54];
  assign o[28039] = i[54];
  assign o[28040] = i[54];
  assign o[28041] = i[54];
  assign o[28042] = i[54];
  assign o[28043] = i[54];
  assign o[28044] = i[54];
  assign o[28045] = i[54];
  assign o[28046] = i[54];
  assign o[28047] = i[54];
  assign o[28048] = i[54];
  assign o[28049] = i[54];
  assign o[28050] = i[54];
  assign o[28051] = i[54];
  assign o[28052] = i[54];
  assign o[28053] = i[54];
  assign o[28054] = i[54];
  assign o[28055] = i[54];
  assign o[28056] = i[54];
  assign o[28057] = i[54];
  assign o[28058] = i[54];
  assign o[28059] = i[54];
  assign o[28060] = i[54];
  assign o[28061] = i[54];
  assign o[28062] = i[54];
  assign o[28063] = i[54];
  assign o[28064] = i[54];
  assign o[28065] = i[54];
  assign o[28066] = i[54];
  assign o[28067] = i[54];
  assign o[28068] = i[54];
  assign o[28069] = i[54];
  assign o[28070] = i[54];
  assign o[28071] = i[54];
  assign o[28072] = i[54];
  assign o[28073] = i[54];
  assign o[28074] = i[54];
  assign o[28075] = i[54];
  assign o[28076] = i[54];
  assign o[28077] = i[54];
  assign o[28078] = i[54];
  assign o[28079] = i[54];
  assign o[28080] = i[54];
  assign o[28081] = i[54];
  assign o[28082] = i[54];
  assign o[28083] = i[54];
  assign o[28084] = i[54];
  assign o[28085] = i[54];
  assign o[28086] = i[54];
  assign o[28087] = i[54];
  assign o[28088] = i[54];
  assign o[28089] = i[54];
  assign o[28090] = i[54];
  assign o[28091] = i[54];
  assign o[28092] = i[54];
  assign o[28093] = i[54];
  assign o[28094] = i[54];
  assign o[28095] = i[54];
  assign o[28096] = i[54];
  assign o[28097] = i[54];
  assign o[28098] = i[54];
  assign o[28099] = i[54];
  assign o[28100] = i[54];
  assign o[28101] = i[54];
  assign o[28102] = i[54];
  assign o[28103] = i[54];
  assign o[28104] = i[54];
  assign o[28105] = i[54];
  assign o[28106] = i[54];
  assign o[28107] = i[54];
  assign o[28108] = i[54];
  assign o[28109] = i[54];
  assign o[28110] = i[54];
  assign o[28111] = i[54];
  assign o[28112] = i[54];
  assign o[28113] = i[54];
  assign o[28114] = i[54];
  assign o[28115] = i[54];
  assign o[28116] = i[54];
  assign o[28117] = i[54];
  assign o[28118] = i[54];
  assign o[28119] = i[54];
  assign o[28120] = i[54];
  assign o[28121] = i[54];
  assign o[28122] = i[54];
  assign o[28123] = i[54];
  assign o[28124] = i[54];
  assign o[28125] = i[54];
  assign o[28126] = i[54];
  assign o[28127] = i[54];
  assign o[28128] = i[54];
  assign o[28129] = i[54];
  assign o[28130] = i[54];
  assign o[28131] = i[54];
  assign o[28132] = i[54];
  assign o[28133] = i[54];
  assign o[28134] = i[54];
  assign o[28135] = i[54];
  assign o[28136] = i[54];
  assign o[28137] = i[54];
  assign o[28138] = i[54];
  assign o[28139] = i[54];
  assign o[28140] = i[54];
  assign o[28141] = i[54];
  assign o[28142] = i[54];
  assign o[28143] = i[54];
  assign o[28144] = i[54];
  assign o[28145] = i[54];
  assign o[28146] = i[54];
  assign o[28147] = i[54];
  assign o[28148] = i[54];
  assign o[28149] = i[54];
  assign o[28150] = i[54];
  assign o[28151] = i[54];
  assign o[28152] = i[54];
  assign o[28153] = i[54];
  assign o[28154] = i[54];
  assign o[28155] = i[54];
  assign o[28156] = i[54];
  assign o[28157] = i[54];
  assign o[28158] = i[54];
  assign o[28159] = i[54];
  assign o[27136] = i[53];
  assign o[27137] = i[53];
  assign o[27138] = i[53];
  assign o[27139] = i[53];
  assign o[27140] = i[53];
  assign o[27141] = i[53];
  assign o[27142] = i[53];
  assign o[27143] = i[53];
  assign o[27144] = i[53];
  assign o[27145] = i[53];
  assign o[27146] = i[53];
  assign o[27147] = i[53];
  assign o[27148] = i[53];
  assign o[27149] = i[53];
  assign o[27150] = i[53];
  assign o[27151] = i[53];
  assign o[27152] = i[53];
  assign o[27153] = i[53];
  assign o[27154] = i[53];
  assign o[27155] = i[53];
  assign o[27156] = i[53];
  assign o[27157] = i[53];
  assign o[27158] = i[53];
  assign o[27159] = i[53];
  assign o[27160] = i[53];
  assign o[27161] = i[53];
  assign o[27162] = i[53];
  assign o[27163] = i[53];
  assign o[27164] = i[53];
  assign o[27165] = i[53];
  assign o[27166] = i[53];
  assign o[27167] = i[53];
  assign o[27168] = i[53];
  assign o[27169] = i[53];
  assign o[27170] = i[53];
  assign o[27171] = i[53];
  assign o[27172] = i[53];
  assign o[27173] = i[53];
  assign o[27174] = i[53];
  assign o[27175] = i[53];
  assign o[27176] = i[53];
  assign o[27177] = i[53];
  assign o[27178] = i[53];
  assign o[27179] = i[53];
  assign o[27180] = i[53];
  assign o[27181] = i[53];
  assign o[27182] = i[53];
  assign o[27183] = i[53];
  assign o[27184] = i[53];
  assign o[27185] = i[53];
  assign o[27186] = i[53];
  assign o[27187] = i[53];
  assign o[27188] = i[53];
  assign o[27189] = i[53];
  assign o[27190] = i[53];
  assign o[27191] = i[53];
  assign o[27192] = i[53];
  assign o[27193] = i[53];
  assign o[27194] = i[53];
  assign o[27195] = i[53];
  assign o[27196] = i[53];
  assign o[27197] = i[53];
  assign o[27198] = i[53];
  assign o[27199] = i[53];
  assign o[27200] = i[53];
  assign o[27201] = i[53];
  assign o[27202] = i[53];
  assign o[27203] = i[53];
  assign o[27204] = i[53];
  assign o[27205] = i[53];
  assign o[27206] = i[53];
  assign o[27207] = i[53];
  assign o[27208] = i[53];
  assign o[27209] = i[53];
  assign o[27210] = i[53];
  assign o[27211] = i[53];
  assign o[27212] = i[53];
  assign o[27213] = i[53];
  assign o[27214] = i[53];
  assign o[27215] = i[53];
  assign o[27216] = i[53];
  assign o[27217] = i[53];
  assign o[27218] = i[53];
  assign o[27219] = i[53];
  assign o[27220] = i[53];
  assign o[27221] = i[53];
  assign o[27222] = i[53];
  assign o[27223] = i[53];
  assign o[27224] = i[53];
  assign o[27225] = i[53];
  assign o[27226] = i[53];
  assign o[27227] = i[53];
  assign o[27228] = i[53];
  assign o[27229] = i[53];
  assign o[27230] = i[53];
  assign o[27231] = i[53];
  assign o[27232] = i[53];
  assign o[27233] = i[53];
  assign o[27234] = i[53];
  assign o[27235] = i[53];
  assign o[27236] = i[53];
  assign o[27237] = i[53];
  assign o[27238] = i[53];
  assign o[27239] = i[53];
  assign o[27240] = i[53];
  assign o[27241] = i[53];
  assign o[27242] = i[53];
  assign o[27243] = i[53];
  assign o[27244] = i[53];
  assign o[27245] = i[53];
  assign o[27246] = i[53];
  assign o[27247] = i[53];
  assign o[27248] = i[53];
  assign o[27249] = i[53];
  assign o[27250] = i[53];
  assign o[27251] = i[53];
  assign o[27252] = i[53];
  assign o[27253] = i[53];
  assign o[27254] = i[53];
  assign o[27255] = i[53];
  assign o[27256] = i[53];
  assign o[27257] = i[53];
  assign o[27258] = i[53];
  assign o[27259] = i[53];
  assign o[27260] = i[53];
  assign o[27261] = i[53];
  assign o[27262] = i[53];
  assign o[27263] = i[53];
  assign o[27264] = i[53];
  assign o[27265] = i[53];
  assign o[27266] = i[53];
  assign o[27267] = i[53];
  assign o[27268] = i[53];
  assign o[27269] = i[53];
  assign o[27270] = i[53];
  assign o[27271] = i[53];
  assign o[27272] = i[53];
  assign o[27273] = i[53];
  assign o[27274] = i[53];
  assign o[27275] = i[53];
  assign o[27276] = i[53];
  assign o[27277] = i[53];
  assign o[27278] = i[53];
  assign o[27279] = i[53];
  assign o[27280] = i[53];
  assign o[27281] = i[53];
  assign o[27282] = i[53];
  assign o[27283] = i[53];
  assign o[27284] = i[53];
  assign o[27285] = i[53];
  assign o[27286] = i[53];
  assign o[27287] = i[53];
  assign o[27288] = i[53];
  assign o[27289] = i[53];
  assign o[27290] = i[53];
  assign o[27291] = i[53];
  assign o[27292] = i[53];
  assign o[27293] = i[53];
  assign o[27294] = i[53];
  assign o[27295] = i[53];
  assign o[27296] = i[53];
  assign o[27297] = i[53];
  assign o[27298] = i[53];
  assign o[27299] = i[53];
  assign o[27300] = i[53];
  assign o[27301] = i[53];
  assign o[27302] = i[53];
  assign o[27303] = i[53];
  assign o[27304] = i[53];
  assign o[27305] = i[53];
  assign o[27306] = i[53];
  assign o[27307] = i[53];
  assign o[27308] = i[53];
  assign o[27309] = i[53];
  assign o[27310] = i[53];
  assign o[27311] = i[53];
  assign o[27312] = i[53];
  assign o[27313] = i[53];
  assign o[27314] = i[53];
  assign o[27315] = i[53];
  assign o[27316] = i[53];
  assign o[27317] = i[53];
  assign o[27318] = i[53];
  assign o[27319] = i[53];
  assign o[27320] = i[53];
  assign o[27321] = i[53];
  assign o[27322] = i[53];
  assign o[27323] = i[53];
  assign o[27324] = i[53];
  assign o[27325] = i[53];
  assign o[27326] = i[53];
  assign o[27327] = i[53];
  assign o[27328] = i[53];
  assign o[27329] = i[53];
  assign o[27330] = i[53];
  assign o[27331] = i[53];
  assign o[27332] = i[53];
  assign o[27333] = i[53];
  assign o[27334] = i[53];
  assign o[27335] = i[53];
  assign o[27336] = i[53];
  assign o[27337] = i[53];
  assign o[27338] = i[53];
  assign o[27339] = i[53];
  assign o[27340] = i[53];
  assign o[27341] = i[53];
  assign o[27342] = i[53];
  assign o[27343] = i[53];
  assign o[27344] = i[53];
  assign o[27345] = i[53];
  assign o[27346] = i[53];
  assign o[27347] = i[53];
  assign o[27348] = i[53];
  assign o[27349] = i[53];
  assign o[27350] = i[53];
  assign o[27351] = i[53];
  assign o[27352] = i[53];
  assign o[27353] = i[53];
  assign o[27354] = i[53];
  assign o[27355] = i[53];
  assign o[27356] = i[53];
  assign o[27357] = i[53];
  assign o[27358] = i[53];
  assign o[27359] = i[53];
  assign o[27360] = i[53];
  assign o[27361] = i[53];
  assign o[27362] = i[53];
  assign o[27363] = i[53];
  assign o[27364] = i[53];
  assign o[27365] = i[53];
  assign o[27366] = i[53];
  assign o[27367] = i[53];
  assign o[27368] = i[53];
  assign o[27369] = i[53];
  assign o[27370] = i[53];
  assign o[27371] = i[53];
  assign o[27372] = i[53];
  assign o[27373] = i[53];
  assign o[27374] = i[53];
  assign o[27375] = i[53];
  assign o[27376] = i[53];
  assign o[27377] = i[53];
  assign o[27378] = i[53];
  assign o[27379] = i[53];
  assign o[27380] = i[53];
  assign o[27381] = i[53];
  assign o[27382] = i[53];
  assign o[27383] = i[53];
  assign o[27384] = i[53];
  assign o[27385] = i[53];
  assign o[27386] = i[53];
  assign o[27387] = i[53];
  assign o[27388] = i[53];
  assign o[27389] = i[53];
  assign o[27390] = i[53];
  assign o[27391] = i[53];
  assign o[27392] = i[53];
  assign o[27393] = i[53];
  assign o[27394] = i[53];
  assign o[27395] = i[53];
  assign o[27396] = i[53];
  assign o[27397] = i[53];
  assign o[27398] = i[53];
  assign o[27399] = i[53];
  assign o[27400] = i[53];
  assign o[27401] = i[53];
  assign o[27402] = i[53];
  assign o[27403] = i[53];
  assign o[27404] = i[53];
  assign o[27405] = i[53];
  assign o[27406] = i[53];
  assign o[27407] = i[53];
  assign o[27408] = i[53];
  assign o[27409] = i[53];
  assign o[27410] = i[53];
  assign o[27411] = i[53];
  assign o[27412] = i[53];
  assign o[27413] = i[53];
  assign o[27414] = i[53];
  assign o[27415] = i[53];
  assign o[27416] = i[53];
  assign o[27417] = i[53];
  assign o[27418] = i[53];
  assign o[27419] = i[53];
  assign o[27420] = i[53];
  assign o[27421] = i[53];
  assign o[27422] = i[53];
  assign o[27423] = i[53];
  assign o[27424] = i[53];
  assign o[27425] = i[53];
  assign o[27426] = i[53];
  assign o[27427] = i[53];
  assign o[27428] = i[53];
  assign o[27429] = i[53];
  assign o[27430] = i[53];
  assign o[27431] = i[53];
  assign o[27432] = i[53];
  assign o[27433] = i[53];
  assign o[27434] = i[53];
  assign o[27435] = i[53];
  assign o[27436] = i[53];
  assign o[27437] = i[53];
  assign o[27438] = i[53];
  assign o[27439] = i[53];
  assign o[27440] = i[53];
  assign o[27441] = i[53];
  assign o[27442] = i[53];
  assign o[27443] = i[53];
  assign o[27444] = i[53];
  assign o[27445] = i[53];
  assign o[27446] = i[53];
  assign o[27447] = i[53];
  assign o[27448] = i[53];
  assign o[27449] = i[53];
  assign o[27450] = i[53];
  assign o[27451] = i[53];
  assign o[27452] = i[53];
  assign o[27453] = i[53];
  assign o[27454] = i[53];
  assign o[27455] = i[53];
  assign o[27456] = i[53];
  assign o[27457] = i[53];
  assign o[27458] = i[53];
  assign o[27459] = i[53];
  assign o[27460] = i[53];
  assign o[27461] = i[53];
  assign o[27462] = i[53];
  assign o[27463] = i[53];
  assign o[27464] = i[53];
  assign o[27465] = i[53];
  assign o[27466] = i[53];
  assign o[27467] = i[53];
  assign o[27468] = i[53];
  assign o[27469] = i[53];
  assign o[27470] = i[53];
  assign o[27471] = i[53];
  assign o[27472] = i[53];
  assign o[27473] = i[53];
  assign o[27474] = i[53];
  assign o[27475] = i[53];
  assign o[27476] = i[53];
  assign o[27477] = i[53];
  assign o[27478] = i[53];
  assign o[27479] = i[53];
  assign o[27480] = i[53];
  assign o[27481] = i[53];
  assign o[27482] = i[53];
  assign o[27483] = i[53];
  assign o[27484] = i[53];
  assign o[27485] = i[53];
  assign o[27486] = i[53];
  assign o[27487] = i[53];
  assign o[27488] = i[53];
  assign o[27489] = i[53];
  assign o[27490] = i[53];
  assign o[27491] = i[53];
  assign o[27492] = i[53];
  assign o[27493] = i[53];
  assign o[27494] = i[53];
  assign o[27495] = i[53];
  assign o[27496] = i[53];
  assign o[27497] = i[53];
  assign o[27498] = i[53];
  assign o[27499] = i[53];
  assign o[27500] = i[53];
  assign o[27501] = i[53];
  assign o[27502] = i[53];
  assign o[27503] = i[53];
  assign o[27504] = i[53];
  assign o[27505] = i[53];
  assign o[27506] = i[53];
  assign o[27507] = i[53];
  assign o[27508] = i[53];
  assign o[27509] = i[53];
  assign o[27510] = i[53];
  assign o[27511] = i[53];
  assign o[27512] = i[53];
  assign o[27513] = i[53];
  assign o[27514] = i[53];
  assign o[27515] = i[53];
  assign o[27516] = i[53];
  assign o[27517] = i[53];
  assign o[27518] = i[53];
  assign o[27519] = i[53];
  assign o[27520] = i[53];
  assign o[27521] = i[53];
  assign o[27522] = i[53];
  assign o[27523] = i[53];
  assign o[27524] = i[53];
  assign o[27525] = i[53];
  assign o[27526] = i[53];
  assign o[27527] = i[53];
  assign o[27528] = i[53];
  assign o[27529] = i[53];
  assign o[27530] = i[53];
  assign o[27531] = i[53];
  assign o[27532] = i[53];
  assign o[27533] = i[53];
  assign o[27534] = i[53];
  assign o[27535] = i[53];
  assign o[27536] = i[53];
  assign o[27537] = i[53];
  assign o[27538] = i[53];
  assign o[27539] = i[53];
  assign o[27540] = i[53];
  assign o[27541] = i[53];
  assign o[27542] = i[53];
  assign o[27543] = i[53];
  assign o[27544] = i[53];
  assign o[27545] = i[53];
  assign o[27546] = i[53];
  assign o[27547] = i[53];
  assign o[27548] = i[53];
  assign o[27549] = i[53];
  assign o[27550] = i[53];
  assign o[27551] = i[53];
  assign o[27552] = i[53];
  assign o[27553] = i[53];
  assign o[27554] = i[53];
  assign o[27555] = i[53];
  assign o[27556] = i[53];
  assign o[27557] = i[53];
  assign o[27558] = i[53];
  assign o[27559] = i[53];
  assign o[27560] = i[53];
  assign o[27561] = i[53];
  assign o[27562] = i[53];
  assign o[27563] = i[53];
  assign o[27564] = i[53];
  assign o[27565] = i[53];
  assign o[27566] = i[53];
  assign o[27567] = i[53];
  assign o[27568] = i[53];
  assign o[27569] = i[53];
  assign o[27570] = i[53];
  assign o[27571] = i[53];
  assign o[27572] = i[53];
  assign o[27573] = i[53];
  assign o[27574] = i[53];
  assign o[27575] = i[53];
  assign o[27576] = i[53];
  assign o[27577] = i[53];
  assign o[27578] = i[53];
  assign o[27579] = i[53];
  assign o[27580] = i[53];
  assign o[27581] = i[53];
  assign o[27582] = i[53];
  assign o[27583] = i[53];
  assign o[27584] = i[53];
  assign o[27585] = i[53];
  assign o[27586] = i[53];
  assign o[27587] = i[53];
  assign o[27588] = i[53];
  assign o[27589] = i[53];
  assign o[27590] = i[53];
  assign o[27591] = i[53];
  assign o[27592] = i[53];
  assign o[27593] = i[53];
  assign o[27594] = i[53];
  assign o[27595] = i[53];
  assign o[27596] = i[53];
  assign o[27597] = i[53];
  assign o[27598] = i[53];
  assign o[27599] = i[53];
  assign o[27600] = i[53];
  assign o[27601] = i[53];
  assign o[27602] = i[53];
  assign o[27603] = i[53];
  assign o[27604] = i[53];
  assign o[27605] = i[53];
  assign o[27606] = i[53];
  assign o[27607] = i[53];
  assign o[27608] = i[53];
  assign o[27609] = i[53];
  assign o[27610] = i[53];
  assign o[27611] = i[53];
  assign o[27612] = i[53];
  assign o[27613] = i[53];
  assign o[27614] = i[53];
  assign o[27615] = i[53];
  assign o[27616] = i[53];
  assign o[27617] = i[53];
  assign o[27618] = i[53];
  assign o[27619] = i[53];
  assign o[27620] = i[53];
  assign o[27621] = i[53];
  assign o[27622] = i[53];
  assign o[27623] = i[53];
  assign o[27624] = i[53];
  assign o[27625] = i[53];
  assign o[27626] = i[53];
  assign o[27627] = i[53];
  assign o[27628] = i[53];
  assign o[27629] = i[53];
  assign o[27630] = i[53];
  assign o[27631] = i[53];
  assign o[27632] = i[53];
  assign o[27633] = i[53];
  assign o[27634] = i[53];
  assign o[27635] = i[53];
  assign o[27636] = i[53];
  assign o[27637] = i[53];
  assign o[27638] = i[53];
  assign o[27639] = i[53];
  assign o[27640] = i[53];
  assign o[27641] = i[53];
  assign o[27642] = i[53];
  assign o[27643] = i[53];
  assign o[27644] = i[53];
  assign o[27645] = i[53];
  assign o[27646] = i[53];
  assign o[27647] = i[53];
  assign o[26624] = i[52];
  assign o[26625] = i[52];
  assign o[26626] = i[52];
  assign o[26627] = i[52];
  assign o[26628] = i[52];
  assign o[26629] = i[52];
  assign o[26630] = i[52];
  assign o[26631] = i[52];
  assign o[26632] = i[52];
  assign o[26633] = i[52];
  assign o[26634] = i[52];
  assign o[26635] = i[52];
  assign o[26636] = i[52];
  assign o[26637] = i[52];
  assign o[26638] = i[52];
  assign o[26639] = i[52];
  assign o[26640] = i[52];
  assign o[26641] = i[52];
  assign o[26642] = i[52];
  assign o[26643] = i[52];
  assign o[26644] = i[52];
  assign o[26645] = i[52];
  assign o[26646] = i[52];
  assign o[26647] = i[52];
  assign o[26648] = i[52];
  assign o[26649] = i[52];
  assign o[26650] = i[52];
  assign o[26651] = i[52];
  assign o[26652] = i[52];
  assign o[26653] = i[52];
  assign o[26654] = i[52];
  assign o[26655] = i[52];
  assign o[26656] = i[52];
  assign o[26657] = i[52];
  assign o[26658] = i[52];
  assign o[26659] = i[52];
  assign o[26660] = i[52];
  assign o[26661] = i[52];
  assign o[26662] = i[52];
  assign o[26663] = i[52];
  assign o[26664] = i[52];
  assign o[26665] = i[52];
  assign o[26666] = i[52];
  assign o[26667] = i[52];
  assign o[26668] = i[52];
  assign o[26669] = i[52];
  assign o[26670] = i[52];
  assign o[26671] = i[52];
  assign o[26672] = i[52];
  assign o[26673] = i[52];
  assign o[26674] = i[52];
  assign o[26675] = i[52];
  assign o[26676] = i[52];
  assign o[26677] = i[52];
  assign o[26678] = i[52];
  assign o[26679] = i[52];
  assign o[26680] = i[52];
  assign o[26681] = i[52];
  assign o[26682] = i[52];
  assign o[26683] = i[52];
  assign o[26684] = i[52];
  assign o[26685] = i[52];
  assign o[26686] = i[52];
  assign o[26687] = i[52];
  assign o[26688] = i[52];
  assign o[26689] = i[52];
  assign o[26690] = i[52];
  assign o[26691] = i[52];
  assign o[26692] = i[52];
  assign o[26693] = i[52];
  assign o[26694] = i[52];
  assign o[26695] = i[52];
  assign o[26696] = i[52];
  assign o[26697] = i[52];
  assign o[26698] = i[52];
  assign o[26699] = i[52];
  assign o[26700] = i[52];
  assign o[26701] = i[52];
  assign o[26702] = i[52];
  assign o[26703] = i[52];
  assign o[26704] = i[52];
  assign o[26705] = i[52];
  assign o[26706] = i[52];
  assign o[26707] = i[52];
  assign o[26708] = i[52];
  assign o[26709] = i[52];
  assign o[26710] = i[52];
  assign o[26711] = i[52];
  assign o[26712] = i[52];
  assign o[26713] = i[52];
  assign o[26714] = i[52];
  assign o[26715] = i[52];
  assign o[26716] = i[52];
  assign o[26717] = i[52];
  assign o[26718] = i[52];
  assign o[26719] = i[52];
  assign o[26720] = i[52];
  assign o[26721] = i[52];
  assign o[26722] = i[52];
  assign o[26723] = i[52];
  assign o[26724] = i[52];
  assign o[26725] = i[52];
  assign o[26726] = i[52];
  assign o[26727] = i[52];
  assign o[26728] = i[52];
  assign o[26729] = i[52];
  assign o[26730] = i[52];
  assign o[26731] = i[52];
  assign o[26732] = i[52];
  assign o[26733] = i[52];
  assign o[26734] = i[52];
  assign o[26735] = i[52];
  assign o[26736] = i[52];
  assign o[26737] = i[52];
  assign o[26738] = i[52];
  assign o[26739] = i[52];
  assign o[26740] = i[52];
  assign o[26741] = i[52];
  assign o[26742] = i[52];
  assign o[26743] = i[52];
  assign o[26744] = i[52];
  assign o[26745] = i[52];
  assign o[26746] = i[52];
  assign o[26747] = i[52];
  assign o[26748] = i[52];
  assign o[26749] = i[52];
  assign o[26750] = i[52];
  assign o[26751] = i[52];
  assign o[26752] = i[52];
  assign o[26753] = i[52];
  assign o[26754] = i[52];
  assign o[26755] = i[52];
  assign o[26756] = i[52];
  assign o[26757] = i[52];
  assign o[26758] = i[52];
  assign o[26759] = i[52];
  assign o[26760] = i[52];
  assign o[26761] = i[52];
  assign o[26762] = i[52];
  assign o[26763] = i[52];
  assign o[26764] = i[52];
  assign o[26765] = i[52];
  assign o[26766] = i[52];
  assign o[26767] = i[52];
  assign o[26768] = i[52];
  assign o[26769] = i[52];
  assign o[26770] = i[52];
  assign o[26771] = i[52];
  assign o[26772] = i[52];
  assign o[26773] = i[52];
  assign o[26774] = i[52];
  assign o[26775] = i[52];
  assign o[26776] = i[52];
  assign o[26777] = i[52];
  assign o[26778] = i[52];
  assign o[26779] = i[52];
  assign o[26780] = i[52];
  assign o[26781] = i[52];
  assign o[26782] = i[52];
  assign o[26783] = i[52];
  assign o[26784] = i[52];
  assign o[26785] = i[52];
  assign o[26786] = i[52];
  assign o[26787] = i[52];
  assign o[26788] = i[52];
  assign o[26789] = i[52];
  assign o[26790] = i[52];
  assign o[26791] = i[52];
  assign o[26792] = i[52];
  assign o[26793] = i[52];
  assign o[26794] = i[52];
  assign o[26795] = i[52];
  assign o[26796] = i[52];
  assign o[26797] = i[52];
  assign o[26798] = i[52];
  assign o[26799] = i[52];
  assign o[26800] = i[52];
  assign o[26801] = i[52];
  assign o[26802] = i[52];
  assign o[26803] = i[52];
  assign o[26804] = i[52];
  assign o[26805] = i[52];
  assign o[26806] = i[52];
  assign o[26807] = i[52];
  assign o[26808] = i[52];
  assign o[26809] = i[52];
  assign o[26810] = i[52];
  assign o[26811] = i[52];
  assign o[26812] = i[52];
  assign o[26813] = i[52];
  assign o[26814] = i[52];
  assign o[26815] = i[52];
  assign o[26816] = i[52];
  assign o[26817] = i[52];
  assign o[26818] = i[52];
  assign o[26819] = i[52];
  assign o[26820] = i[52];
  assign o[26821] = i[52];
  assign o[26822] = i[52];
  assign o[26823] = i[52];
  assign o[26824] = i[52];
  assign o[26825] = i[52];
  assign o[26826] = i[52];
  assign o[26827] = i[52];
  assign o[26828] = i[52];
  assign o[26829] = i[52];
  assign o[26830] = i[52];
  assign o[26831] = i[52];
  assign o[26832] = i[52];
  assign o[26833] = i[52];
  assign o[26834] = i[52];
  assign o[26835] = i[52];
  assign o[26836] = i[52];
  assign o[26837] = i[52];
  assign o[26838] = i[52];
  assign o[26839] = i[52];
  assign o[26840] = i[52];
  assign o[26841] = i[52];
  assign o[26842] = i[52];
  assign o[26843] = i[52];
  assign o[26844] = i[52];
  assign o[26845] = i[52];
  assign o[26846] = i[52];
  assign o[26847] = i[52];
  assign o[26848] = i[52];
  assign o[26849] = i[52];
  assign o[26850] = i[52];
  assign o[26851] = i[52];
  assign o[26852] = i[52];
  assign o[26853] = i[52];
  assign o[26854] = i[52];
  assign o[26855] = i[52];
  assign o[26856] = i[52];
  assign o[26857] = i[52];
  assign o[26858] = i[52];
  assign o[26859] = i[52];
  assign o[26860] = i[52];
  assign o[26861] = i[52];
  assign o[26862] = i[52];
  assign o[26863] = i[52];
  assign o[26864] = i[52];
  assign o[26865] = i[52];
  assign o[26866] = i[52];
  assign o[26867] = i[52];
  assign o[26868] = i[52];
  assign o[26869] = i[52];
  assign o[26870] = i[52];
  assign o[26871] = i[52];
  assign o[26872] = i[52];
  assign o[26873] = i[52];
  assign o[26874] = i[52];
  assign o[26875] = i[52];
  assign o[26876] = i[52];
  assign o[26877] = i[52];
  assign o[26878] = i[52];
  assign o[26879] = i[52];
  assign o[26880] = i[52];
  assign o[26881] = i[52];
  assign o[26882] = i[52];
  assign o[26883] = i[52];
  assign o[26884] = i[52];
  assign o[26885] = i[52];
  assign o[26886] = i[52];
  assign o[26887] = i[52];
  assign o[26888] = i[52];
  assign o[26889] = i[52];
  assign o[26890] = i[52];
  assign o[26891] = i[52];
  assign o[26892] = i[52];
  assign o[26893] = i[52];
  assign o[26894] = i[52];
  assign o[26895] = i[52];
  assign o[26896] = i[52];
  assign o[26897] = i[52];
  assign o[26898] = i[52];
  assign o[26899] = i[52];
  assign o[26900] = i[52];
  assign o[26901] = i[52];
  assign o[26902] = i[52];
  assign o[26903] = i[52];
  assign o[26904] = i[52];
  assign o[26905] = i[52];
  assign o[26906] = i[52];
  assign o[26907] = i[52];
  assign o[26908] = i[52];
  assign o[26909] = i[52];
  assign o[26910] = i[52];
  assign o[26911] = i[52];
  assign o[26912] = i[52];
  assign o[26913] = i[52];
  assign o[26914] = i[52];
  assign o[26915] = i[52];
  assign o[26916] = i[52];
  assign o[26917] = i[52];
  assign o[26918] = i[52];
  assign o[26919] = i[52];
  assign o[26920] = i[52];
  assign o[26921] = i[52];
  assign o[26922] = i[52];
  assign o[26923] = i[52];
  assign o[26924] = i[52];
  assign o[26925] = i[52];
  assign o[26926] = i[52];
  assign o[26927] = i[52];
  assign o[26928] = i[52];
  assign o[26929] = i[52];
  assign o[26930] = i[52];
  assign o[26931] = i[52];
  assign o[26932] = i[52];
  assign o[26933] = i[52];
  assign o[26934] = i[52];
  assign o[26935] = i[52];
  assign o[26936] = i[52];
  assign o[26937] = i[52];
  assign o[26938] = i[52];
  assign o[26939] = i[52];
  assign o[26940] = i[52];
  assign o[26941] = i[52];
  assign o[26942] = i[52];
  assign o[26943] = i[52];
  assign o[26944] = i[52];
  assign o[26945] = i[52];
  assign o[26946] = i[52];
  assign o[26947] = i[52];
  assign o[26948] = i[52];
  assign o[26949] = i[52];
  assign o[26950] = i[52];
  assign o[26951] = i[52];
  assign o[26952] = i[52];
  assign o[26953] = i[52];
  assign o[26954] = i[52];
  assign o[26955] = i[52];
  assign o[26956] = i[52];
  assign o[26957] = i[52];
  assign o[26958] = i[52];
  assign o[26959] = i[52];
  assign o[26960] = i[52];
  assign o[26961] = i[52];
  assign o[26962] = i[52];
  assign o[26963] = i[52];
  assign o[26964] = i[52];
  assign o[26965] = i[52];
  assign o[26966] = i[52];
  assign o[26967] = i[52];
  assign o[26968] = i[52];
  assign o[26969] = i[52];
  assign o[26970] = i[52];
  assign o[26971] = i[52];
  assign o[26972] = i[52];
  assign o[26973] = i[52];
  assign o[26974] = i[52];
  assign o[26975] = i[52];
  assign o[26976] = i[52];
  assign o[26977] = i[52];
  assign o[26978] = i[52];
  assign o[26979] = i[52];
  assign o[26980] = i[52];
  assign o[26981] = i[52];
  assign o[26982] = i[52];
  assign o[26983] = i[52];
  assign o[26984] = i[52];
  assign o[26985] = i[52];
  assign o[26986] = i[52];
  assign o[26987] = i[52];
  assign o[26988] = i[52];
  assign o[26989] = i[52];
  assign o[26990] = i[52];
  assign o[26991] = i[52];
  assign o[26992] = i[52];
  assign o[26993] = i[52];
  assign o[26994] = i[52];
  assign o[26995] = i[52];
  assign o[26996] = i[52];
  assign o[26997] = i[52];
  assign o[26998] = i[52];
  assign o[26999] = i[52];
  assign o[27000] = i[52];
  assign o[27001] = i[52];
  assign o[27002] = i[52];
  assign o[27003] = i[52];
  assign o[27004] = i[52];
  assign o[27005] = i[52];
  assign o[27006] = i[52];
  assign o[27007] = i[52];
  assign o[27008] = i[52];
  assign o[27009] = i[52];
  assign o[27010] = i[52];
  assign o[27011] = i[52];
  assign o[27012] = i[52];
  assign o[27013] = i[52];
  assign o[27014] = i[52];
  assign o[27015] = i[52];
  assign o[27016] = i[52];
  assign o[27017] = i[52];
  assign o[27018] = i[52];
  assign o[27019] = i[52];
  assign o[27020] = i[52];
  assign o[27021] = i[52];
  assign o[27022] = i[52];
  assign o[27023] = i[52];
  assign o[27024] = i[52];
  assign o[27025] = i[52];
  assign o[27026] = i[52];
  assign o[27027] = i[52];
  assign o[27028] = i[52];
  assign o[27029] = i[52];
  assign o[27030] = i[52];
  assign o[27031] = i[52];
  assign o[27032] = i[52];
  assign o[27033] = i[52];
  assign o[27034] = i[52];
  assign o[27035] = i[52];
  assign o[27036] = i[52];
  assign o[27037] = i[52];
  assign o[27038] = i[52];
  assign o[27039] = i[52];
  assign o[27040] = i[52];
  assign o[27041] = i[52];
  assign o[27042] = i[52];
  assign o[27043] = i[52];
  assign o[27044] = i[52];
  assign o[27045] = i[52];
  assign o[27046] = i[52];
  assign o[27047] = i[52];
  assign o[27048] = i[52];
  assign o[27049] = i[52];
  assign o[27050] = i[52];
  assign o[27051] = i[52];
  assign o[27052] = i[52];
  assign o[27053] = i[52];
  assign o[27054] = i[52];
  assign o[27055] = i[52];
  assign o[27056] = i[52];
  assign o[27057] = i[52];
  assign o[27058] = i[52];
  assign o[27059] = i[52];
  assign o[27060] = i[52];
  assign o[27061] = i[52];
  assign o[27062] = i[52];
  assign o[27063] = i[52];
  assign o[27064] = i[52];
  assign o[27065] = i[52];
  assign o[27066] = i[52];
  assign o[27067] = i[52];
  assign o[27068] = i[52];
  assign o[27069] = i[52];
  assign o[27070] = i[52];
  assign o[27071] = i[52];
  assign o[27072] = i[52];
  assign o[27073] = i[52];
  assign o[27074] = i[52];
  assign o[27075] = i[52];
  assign o[27076] = i[52];
  assign o[27077] = i[52];
  assign o[27078] = i[52];
  assign o[27079] = i[52];
  assign o[27080] = i[52];
  assign o[27081] = i[52];
  assign o[27082] = i[52];
  assign o[27083] = i[52];
  assign o[27084] = i[52];
  assign o[27085] = i[52];
  assign o[27086] = i[52];
  assign o[27087] = i[52];
  assign o[27088] = i[52];
  assign o[27089] = i[52];
  assign o[27090] = i[52];
  assign o[27091] = i[52];
  assign o[27092] = i[52];
  assign o[27093] = i[52];
  assign o[27094] = i[52];
  assign o[27095] = i[52];
  assign o[27096] = i[52];
  assign o[27097] = i[52];
  assign o[27098] = i[52];
  assign o[27099] = i[52];
  assign o[27100] = i[52];
  assign o[27101] = i[52];
  assign o[27102] = i[52];
  assign o[27103] = i[52];
  assign o[27104] = i[52];
  assign o[27105] = i[52];
  assign o[27106] = i[52];
  assign o[27107] = i[52];
  assign o[27108] = i[52];
  assign o[27109] = i[52];
  assign o[27110] = i[52];
  assign o[27111] = i[52];
  assign o[27112] = i[52];
  assign o[27113] = i[52];
  assign o[27114] = i[52];
  assign o[27115] = i[52];
  assign o[27116] = i[52];
  assign o[27117] = i[52];
  assign o[27118] = i[52];
  assign o[27119] = i[52];
  assign o[27120] = i[52];
  assign o[27121] = i[52];
  assign o[27122] = i[52];
  assign o[27123] = i[52];
  assign o[27124] = i[52];
  assign o[27125] = i[52];
  assign o[27126] = i[52];
  assign o[27127] = i[52];
  assign o[27128] = i[52];
  assign o[27129] = i[52];
  assign o[27130] = i[52];
  assign o[27131] = i[52];
  assign o[27132] = i[52];
  assign o[27133] = i[52];
  assign o[27134] = i[52];
  assign o[27135] = i[52];
  assign o[26112] = i[51];
  assign o[26113] = i[51];
  assign o[26114] = i[51];
  assign o[26115] = i[51];
  assign o[26116] = i[51];
  assign o[26117] = i[51];
  assign o[26118] = i[51];
  assign o[26119] = i[51];
  assign o[26120] = i[51];
  assign o[26121] = i[51];
  assign o[26122] = i[51];
  assign o[26123] = i[51];
  assign o[26124] = i[51];
  assign o[26125] = i[51];
  assign o[26126] = i[51];
  assign o[26127] = i[51];
  assign o[26128] = i[51];
  assign o[26129] = i[51];
  assign o[26130] = i[51];
  assign o[26131] = i[51];
  assign o[26132] = i[51];
  assign o[26133] = i[51];
  assign o[26134] = i[51];
  assign o[26135] = i[51];
  assign o[26136] = i[51];
  assign o[26137] = i[51];
  assign o[26138] = i[51];
  assign o[26139] = i[51];
  assign o[26140] = i[51];
  assign o[26141] = i[51];
  assign o[26142] = i[51];
  assign o[26143] = i[51];
  assign o[26144] = i[51];
  assign o[26145] = i[51];
  assign o[26146] = i[51];
  assign o[26147] = i[51];
  assign o[26148] = i[51];
  assign o[26149] = i[51];
  assign o[26150] = i[51];
  assign o[26151] = i[51];
  assign o[26152] = i[51];
  assign o[26153] = i[51];
  assign o[26154] = i[51];
  assign o[26155] = i[51];
  assign o[26156] = i[51];
  assign o[26157] = i[51];
  assign o[26158] = i[51];
  assign o[26159] = i[51];
  assign o[26160] = i[51];
  assign o[26161] = i[51];
  assign o[26162] = i[51];
  assign o[26163] = i[51];
  assign o[26164] = i[51];
  assign o[26165] = i[51];
  assign o[26166] = i[51];
  assign o[26167] = i[51];
  assign o[26168] = i[51];
  assign o[26169] = i[51];
  assign o[26170] = i[51];
  assign o[26171] = i[51];
  assign o[26172] = i[51];
  assign o[26173] = i[51];
  assign o[26174] = i[51];
  assign o[26175] = i[51];
  assign o[26176] = i[51];
  assign o[26177] = i[51];
  assign o[26178] = i[51];
  assign o[26179] = i[51];
  assign o[26180] = i[51];
  assign o[26181] = i[51];
  assign o[26182] = i[51];
  assign o[26183] = i[51];
  assign o[26184] = i[51];
  assign o[26185] = i[51];
  assign o[26186] = i[51];
  assign o[26187] = i[51];
  assign o[26188] = i[51];
  assign o[26189] = i[51];
  assign o[26190] = i[51];
  assign o[26191] = i[51];
  assign o[26192] = i[51];
  assign o[26193] = i[51];
  assign o[26194] = i[51];
  assign o[26195] = i[51];
  assign o[26196] = i[51];
  assign o[26197] = i[51];
  assign o[26198] = i[51];
  assign o[26199] = i[51];
  assign o[26200] = i[51];
  assign o[26201] = i[51];
  assign o[26202] = i[51];
  assign o[26203] = i[51];
  assign o[26204] = i[51];
  assign o[26205] = i[51];
  assign o[26206] = i[51];
  assign o[26207] = i[51];
  assign o[26208] = i[51];
  assign o[26209] = i[51];
  assign o[26210] = i[51];
  assign o[26211] = i[51];
  assign o[26212] = i[51];
  assign o[26213] = i[51];
  assign o[26214] = i[51];
  assign o[26215] = i[51];
  assign o[26216] = i[51];
  assign o[26217] = i[51];
  assign o[26218] = i[51];
  assign o[26219] = i[51];
  assign o[26220] = i[51];
  assign o[26221] = i[51];
  assign o[26222] = i[51];
  assign o[26223] = i[51];
  assign o[26224] = i[51];
  assign o[26225] = i[51];
  assign o[26226] = i[51];
  assign o[26227] = i[51];
  assign o[26228] = i[51];
  assign o[26229] = i[51];
  assign o[26230] = i[51];
  assign o[26231] = i[51];
  assign o[26232] = i[51];
  assign o[26233] = i[51];
  assign o[26234] = i[51];
  assign o[26235] = i[51];
  assign o[26236] = i[51];
  assign o[26237] = i[51];
  assign o[26238] = i[51];
  assign o[26239] = i[51];
  assign o[26240] = i[51];
  assign o[26241] = i[51];
  assign o[26242] = i[51];
  assign o[26243] = i[51];
  assign o[26244] = i[51];
  assign o[26245] = i[51];
  assign o[26246] = i[51];
  assign o[26247] = i[51];
  assign o[26248] = i[51];
  assign o[26249] = i[51];
  assign o[26250] = i[51];
  assign o[26251] = i[51];
  assign o[26252] = i[51];
  assign o[26253] = i[51];
  assign o[26254] = i[51];
  assign o[26255] = i[51];
  assign o[26256] = i[51];
  assign o[26257] = i[51];
  assign o[26258] = i[51];
  assign o[26259] = i[51];
  assign o[26260] = i[51];
  assign o[26261] = i[51];
  assign o[26262] = i[51];
  assign o[26263] = i[51];
  assign o[26264] = i[51];
  assign o[26265] = i[51];
  assign o[26266] = i[51];
  assign o[26267] = i[51];
  assign o[26268] = i[51];
  assign o[26269] = i[51];
  assign o[26270] = i[51];
  assign o[26271] = i[51];
  assign o[26272] = i[51];
  assign o[26273] = i[51];
  assign o[26274] = i[51];
  assign o[26275] = i[51];
  assign o[26276] = i[51];
  assign o[26277] = i[51];
  assign o[26278] = i[51];
  assign o[26279] = i[51];
  assign o[26280] = i[51];
  assign o[26281] = i[51];
  assign o[26282] = i[51];
  assign o[26283] = i[51];
  assign o[26284] = i[51];
  assign o[26285] = i[51];
  assign o[26286] = i[51];
  assign o[26287] = i[51];
  assign o[26288] = i[51];
  assign o[26289] = i[51];
  assign o[26290] = i[51];
  assign o[26291] = i[51];
  assign o[26292] = i[51];
  assign o[26293] = i[51];
  assign o[26294] = i[51];
  assign o[26295] = i[51];
  assign o[26296] = i[51];
  assign o[26297] = i[51];
  assign o[26298] = i[51];
  assign o[26299] = i[51];
  assign o[26300] = i[51];
  assign o[26301] = i[51];
  assign o[26302] = i[51];
  assign o[26303] = i[51];
  assign o[26304] = i[51];
  assign o[26305] = i[51];
  assign o[26306] = i[51];
  assign o[26307] = i[51];
  assign o[26308] = i[51];
  assign o[26309] = i[51];
  assign o[26310] = i[51];
  assign o[26311] = i[51];
  assign o[26312] = i[51];
  assign o[26313] = i[51];
  assign o[26314] = i[51];
  assign o[26315] = i[51];
  assign o[26316] = i[51];
  assign o[26317] = i[51];
  assign o[26318] = i[51];
  assign o[26319] = i[51];
  assign o[26320] = i[51];
  assign o[26321] = i[51];
  assign o[26322] = i[51];
  assign o[26323] = i[51];
  assign o[26324] = i[51];
  assign o[26325] = i[51];
  assign o[26326] = i[51];
  assign o[26327] = i[51];
  assign o[26328] = i[51];
  assign o[26329] = i[51];
  assign o[26330] = i[51];
  assign o[26331] = i[51];
  assign o[26332] = i[51];
  assign o[26333] = i[51];
  assign o[26334] = i[51];
  assign o[26335] = i[51];
  assign o[26336] = i[51];
  assign o[26337] = i[51];
  assign o[26338] = i[51];
  assign o[26339] = i[51];
  assign o[26340] = i[51];
  assign o[26341] = i[51];
  assign o[26342] = i[51];
  assign o[26343] = i[51];
  assign o[26344] = i[51];
  assign o[26345] = i[51];
  assign o[26346] = i[51];
  assign o[26347] = i[51];
  assign o[26348] = i[51];
  assign o[26349] = i[51];
  assign o[26350] = i[51];
  assign o[26351] = i[51];
  assign o[26352] = i[51];
  assign o[26353] = i[51];
  assign o[26354] = i[51];
  assign o[26355] = i[51];
  assign o[26356] = i[51];
  assign o[26357] = i[51];
  assign o[26358] = i[51];
  assign o[26359] = i[51];
  assign o[26360] = i[51];
  assign o[26361] = i[51];
  assign o[26362] = i[51];
  assign o[26363] = i[51];
  assign o[26364] = i[51];
  assign o[26365] = i[51];
  assign o[26366] = i[51];
  assign o[26367] = i[51];
  assign o[26368] = i[51];
  assign o[26369] = i[51];
  assign o[26370] = i[51];
  assign o[26371] = i[51];
  assign o[26372] = i[51];
  assign o[26373] = i[51];
  assign o[26374] = i[51];
  assign o[26375] = i[51];
  assign o[26376] = i[51];
  assign o[26377] = i[51];
  assign o[26378] = i[51];
  assign o[26379] = i[51];
  assign o[26380] = i[51];
  assign o[26381] = i[51];
  assign o[26382] = i[51];
  assign o[26383] = i[51];
  assign o[26384] = i[51];
  assign o[26385] = i[51];
  assign o[26386] = i[51];
  assign o[26387] = i[51];
  assign o[26388] = i[51];
  assign o[26389] = i[51];
  assign o[26390] = i[51];
  assign o[26391] = i[51];
  assign o[26392] = i[51];
  assign o[26393] = i[51];
  assign o[26394] = i[51];
  assign o[26395] = i[51];
  assign o[26396] = i[51];
  assign o[26397] = i[51];
  assign o[26398] = i[51];
  assign o[26399] = i[51];
  assign o[26400] = i[51];
  assign o[26401] = i[51];
  assign o[26402] = i[51];
  assign o[26403] = i[51];
  assign o[26404] = i[51];
  assign o[26405] = i[51];
  assign o[26406] = i[51];
  assign o[26407] = i[51];
  assign o[26408] = i[51];
  assign o[26409] = i[51];
  assign o[26410] = i[51];
  assign o[26411] = i[51];
  assign o[26412] = i[51];
  assign o[26413] = i[51];
  assign o[26414] = i[51];
  assign o[26415] = i[51];
  assign o[26416] = i[51];
  assign o[26417] = i[51];
  assign o[26418] = i[51];
  assign o[26419] = i[51];
  assign o[26420] = i[51];
  assign o[26421] = i[51];
  assign o[26422] = i[51];
  assign o[26423] = i[51];
  assign o[26424] = i[51];
  assign o[26425] = i[51];
  assign o[26426] = i[51];
  assign o[26427] = i[51];
  assign o[26428] = i[51];
  assign o[26429] = i[51];
  assign o[26430] = i[51];
  assign o[26431] = i[51];
  assign o[26432] = i[51];
  assign o[26433] = i[51];
  assign o[26434] = i[51];
  assign o[26435] = i[51];
  assign o[26436] = i[51];
  assign o[26437] = i[51];
  assign o[26438] = i[51];
  assign o[26439] = i[51];
  assign o[26440] = i[51];
  assign o[26441] = i[51];
  assign o[26442] = i[51];
  assign o[26443] = i[51];
  assign o[26444] = i[51];
  assign o[26445] = i[51];
  assign o[26446] = i[51];
  assign o[26447] = i[51];
  assign o[26448] = i[51];
  assign o[26449] = i[51];
  assign o[26450] = i[51];
  assign o[26451] = i[51];
  assign o[26452] = i[51];
  assign o[26453] = i[51];
  assign o[26454] = i[51];
  assign o[26455] = i[51];
  assign o[26456] = i[51];
  assign o[26457] = i[51];
  assign o[26458] = i[51];
  assign o[26459] = i[51];
  assign o[26460] = i[51];
  assign o[26461] = i[51];
  assign o[26462] = i[51];
  assign o[26463] = i[51];
  assign o[26464] = i[51];
  assign o[26465] = i[51];
  assign o[26466] = i[51];
  assign o[26467] = i[51];
  assign o[26468] = i[51];
  assign o[26469] = i[51];
  assign o[26470] = i[51];
  assign o[26471] = i[51];
  assign o[26472] = i[51];
  assign o[26473] = i[51];
  assign o[26474] = i[51];
  assign o[26475] = i[51];
  assign o[26476] = i[51];
  assign o[26477] = i[51];
  assign o[26478] = i[51];
  assign o[26479] = i[51];
  assign o[26480] = i[51];
  assign o[26481] = i[51];
  assign o[26482] = i[51];
  assign o[26483] = i[51];
  assign o[26484] = i[51];
  assign o[26485] = i[51];
  assign o[26486] = i[51];
  assign o[26487] = i[51];
  assign o[26488] = i[51];
  assign o[26489] = i[51];
  assign o[26490] = i[51];
  assign o[26491] = i[51];
  assign o[26492] = i[51];
  assign o[26493] = i[51];
  assign o[26494] = i[51];
  assign o[26495] = i[51];
  assign o[26496] = i[51];
  assign o[26497] = i[51];
  assign o[26498] = i[51];
  assign o[26499] = i[51];
  assign o[26500] = i[51];
  assign o[26501] = i[51];
  assign o[26502] = i[51];
  assign o[26503] = i[51];
  assign o[26504] = i[51];
  assign o[26505] = i[51];
  assign o[26506] = i[51];
  assign o[26507] = i[51];
  assign o[26508] = i[51];
  assign o[26509] = i[51];
  assign o[26510] = i[51];
  assign o[26511] = i[51];
  assign o[26512] = i[51];
  assign o[26513] = i[51];
  assign o[26514] = i[51];
  assign o[26515] = i[51];
  assign o[26516] = i[51];
  assign o[26517] = i[51];
  assign o[26518] = i[51];
  assign o[26519] = i[51];
  assign o[26520] = i[51];
  assign o[26521] = i[51];
  assign o[26522] = i[51];
  assign o[26523] = i[51];
  assign o[26524] = i[51];
  assign o[26525] = i[51];
  assign o[26526] = i[51];
  assign o[26527] = i[51];
  assign o[26528] = i[51];
  assign o[26529] = i[51];
  assign o[26530] = i[51];
  assign o[26531] = i[51];
  assign o[26532] = i[51];
  assign o[26533] = i[51];
  assign o[26534] = i[51];
  assign o[26535] = i[51];
  assign o[26536] = i[51];
  assign o[26537] = i[51];
  assign o[26538] = i[51];
  assign o[26539] = i[51];
  assign o[26540] = i[51];
  assign o[26541] = i[51];
  assign o[26542] = i[51];
  assign o[26543] = i[51];
  assign o[26544] = i[51];
  assign o[26545] = i[51];
  assign o[26546] = i[51];
  assign o[26547] = i[51];
  assign o[26548] = i[51];
  assign o[26549] = i[51];
  assign o[26550] = i[51];
  assign o[26551] = i[51];
  assign o[26552] = i[51];
  assign o[26553] = i[51];
  assign o[26554] = i[51];
  assign o[26555] = i[51];
  assign o[26556] = i[51];
  assign o[26557] = i[51];
  assign o[26558] = i[51];
  assign o[26559] = i[51];
  assign o[26560] = i[51];
  assign o[26561] = i[51];
  assign o[26562] = i[51];
  assign o[26563] = i[51];
  assign o[26564] = i[51];
  assign o[26565] = i[51];
  assign o[26566] = i[51];
  assign o[26567] = i[51];
  assign o[26568] = i[51];
  assign o[26569] = i[51];
  assign o[26570] = i[51];
  assign o[26571] = i[51];
  assign o[26572] = i[51];
  assign o[26573] = i[51];
  assign o[26574] = i[51];
  assign o[26575] = i[51];
  assign o[26576] = i[51];
  assign o[26577] = i[51];
  assign o[26578] = i[51];
  assign o[26579] = i[51];
  assign o[26580] = i[51];
  assign o[26581] = i[51];
  assign o[26582] = i[51];
  assign o[26583] = i[51];
  assign o[26584] = i[51];
  assign o[26585] = i[51];
  assign o[26586] = i[51];
  assign o[26587] = i[51];
  assign o[26588] = i[51];
  assign o[26589] = i[51];
  assign o[26590] = i[51];
  assign o[26591] = i[51];
  assign o[26592] = i[51];
  assign o[26593] = i[51];
  assign o[26594] = i[51];
  assign o[26595] = i[51];
  assign o[26596] = i[51];
  assign o[26597] = i[51];
  assign o[26598] = i[51];
  assign o[26599] = i[51];
  assign o[26600] = i[51];
  assign o[26601] = i[51];
  assign o[26602] = i[51];
  assign o[26603] = i[51];
  assign o[26604] = i[51];
  assign o[26605] = i[51];
  assign o[26606] = i[51];
  assign o[26607] = i[51];
  assign o[26608] = i[51];
  assign o[26609] = i[51];
  assign o[26610] = i[51];
  assign o[26611] = i[51];
  assign o[26612] = i[51];
  assign o[26613] = i[51];
  assign o[26614] = i[51];
  assign o[26615] = i[51];
  assign o[26616] = i[51];
  assign o[26617] = i[51];
  assign o[26618] = i[51];
  assign o[26619] = i[51];
  assign o[26620] = i[51];
  assign o[26621] = i[51];
  assign o[26622] = i[51];
  assign o[26623] = i[51];
  assign o[25600] = i[50];
  assign o[25601] = i[50];
  assign o[25602] = i[50];
  assign o[25603] = i[50];
  assign o[25604] = i[50];
  assign o[25605] = i[50];
  assign o[25606] = i[50];
  assign o[25607] = i[50];
  assign o[25608] = i[50];
  assign o[25609] = i[50];
  assign o[25610] = i[50];
  assign o[25611] = i[50];
  assign o[25612] = i[50];
  assign o[25613] = i[50];
  assign o[25614] = i[50];
  assign o[25615] = i[50];
  assign o[25616] = i[50];
  assign o[25617] = i[50];
  assign o[25618] = i[50];
  assign o[25619] = i[50];
  assign o[25620] = i[50];
  assign o[25621] = i[50];
  assign o[25622] = i[50];
  assign o[25623] = i[50];
  assign o[25624] = i[50];
  assign o[25625] = i[50];
  assign o[25626] = i[50];
  assign o[25627] = i[50];
  assign o[25628] = i[50];
  assign o[25629] = i[50];
  assign o[25630] = i[50];
  assign o[25631] = i[50];
  assign o[25632] = i[50];
  assign o[25633] = i[50];
  assign o[25634] = i[50];
  assign o[25635] = i[50];
  assign o[25636] = i[50];
  assign o[25637] = i[50];
  assign o[25638] = i[50];
  assign o[25639] = i[50];
  assign o[25640] = i[50];
  assign o[25641] = i[50];
  assign o[25642] = i[50];
  assign o[25643] = i[50];
  assign o[25644] = i[50];
  assign o[25645] = i[50];
  assign o[25646] = i[50];
  assign o[25647] = i[50];
  assign o[25648] = i[50];
  assign o[25649] = i[50];
  assign o[25650] = i[50];
  assign o[25651] = i[50];
  assign o[25652] = i[50];
  assign o[25653] = i[50];
  assign o[25654] = i[50];
  assign o[25655] = i[50];
  assign o[25656] = i[50];
  assign o[25657] = i[50];
  assign o[25658] = i[50];
  assign o[25659] = i[50];
  assign o[25660] = i[50];
  assign o[25661] = i[50];
  assign o[25662] = i[50];
  assign o[25663] = i[50];
  assign o[25664] = i[50];
  assign o[25665] = i[50];
  assign o[25666] = i[50];
  assign o[25667] = i[50];
  assign o[25668] = i[50];
  assign o[25669] = i[50];
  assign o[25670] = i[50];
  assign o[25671] = i[50];
  assign o[25672] = i[50];
  assign o[25673] = i[50];
  assign o[25674] = i[50];
  assign o[25675] = i[50];
  assign o[25676] = i[50];
  assign o[25677] = i[50];
  assign o[25678] = i[50];
  assign o[25679] = i[50];
  assign o[25680] = i[50];
  assign o[25681] = i[50];
  assign o[25682] = i[50];
  assign o[25683] = i[50];
  assign o[25684] = i[50];
  assign o[25685] = i[50];
  assign o[25686] = i[50];
  assign o[25687] = i[50];
  assign o[25688] = i[50];
  assign o[25689] = i[50];
  assign o[25690] = i[50];
  assign o[25691] = i[50];
  assign o[25692] = i[50];
  assign o[25693] = i[50];
  assign o[25694] = i[50];
  assign o[25695] = i[50];
  assign o[25696] = i[50];
  assign o[25697] = i[50];
  assign o[25698] = i[50];
  assign o[25699] = i[50];
  assign o[25700] = i[50];
  assign o[25701] = i[50];
  assign o[25702] = i[50];
  assign o[25703] = i[50];
  assign o[25704] = i[50];
  assign o[25705] = i[50];
  assign o[25706] = i[50];
  assign o[25707] = i[50];
  assign o[25708] = i[50];
  assign o[25709] = i[50];
  assign o[25710] = i[50];
  assign o[25711] = i[50];
  assign o[25712] = i[50];
  assign o[25713] = i[50];
  assign o[25714] = i[50];
  assign o[25715] = i[50];
  assign o[25716] = i[50];
  assign o[25717] = i[50];
  assign o[25718] = i[50];
  assign o[25719] = i[50];
  assign o[25720] = i[50];
  assign o[25721] = i[50];
  assign o[25722] = i[50];
  assign o[25723] = i[50];
  assign o[25724] = i[50];
  assign o[25725] = i[50];
  assign o[25726] = i[50];
  assign o[25727] = i[50];
  assign o[25728] = i[50];
  assign o[25729] = i[50];
  assign o[25730] = i[50];
  assign o[25731] = i[50];
  assign o[25732] = i[50];
  assign o[25733] = i[50];
  assign o[25734] = i[50];
  assign o[25735] = i[50];
  assign o[25736] = i[50];
  assign o[25737] = i[50];
  assign o[25738] = i[50];
  assign o[25739] = i[50];
  assign o[25740] = i[50];
  assign o[25741] = i[50];
  assign o[25742] = i[50];
  assign o[25743] = i[50];
  assign o[25744] = i[50];
  assign o[25745] = i[50];
  assign o[25746] = i[50];
  assign o[25747] = i[50];
  assign o[25748] = i[50];
  assign o[25749] = i[50];
  assign o[25750] = i[50];
  assign o[25751] = i[50];
  assign o[25752] = i[50];
  assign o[25753] = i[50];
  assign o[25754] = i[50];
  assign o[25755] = i[50];
  assign o[25756] = i[50];
  assign o[25757] = i[50];
  assign o[25758] = i[50];
  assign o[25759] = i[50];
  assign o[25760] = i[50];
  assign o[25761] = i[50];
  assign o[25762] = i[50];
  assign o[25763] = i[50];
  assign o[25764] = i[50];
  assign o[25765] = i[50];
  assign o[25766] = i[50];
  assign o[25767] = i[50];
  assign o[25768] = i[50];
  assign o[25769] = i[50];
  assign o[25770] = i[50];
  assign o[25771] = i[50];
  assign o[25772] = i[50];
  assign o[25773] = i[50];
  assign o[25774] = i[50];
  assign o[25775] = i[50];
  assign o[25776] = i[50];
  assign o[25777] = i[50];
  assign o[25778] = i[50];
  assign o[25779] = i[50];
  assign o[25780] = i[50];
  assign o[25781] = i[50];
  assign o[25782] = i[50];
  assign o[25783] = i[50];
  assign o[25784] = i[50];
  assign o[25785] = i[50];
  assign o[25786] = i[50];
  assign o[25787] = i[50];
  assign o[25788] = i[50];
  assign o[25789] = i[50];
  assign o[25790] = i[50];
  assign o[25791] = i[50];
  assign o[25792] = i[50];
  assign o[25793] = i[50];
  assign o[25794] = i[50];
  assign o[25795] = i[50];
  assign o[25796] = i[50];
  assign o[25797] = i[50];
  assign o[25798] = i[50];
  assign o[25799] = i[50];
  assign o[25800] = i[50];
  assign o[25801] = i[50];
  assign o[25802] = i[50];
  assign o[25803] = i[50];
  assign o[25804] = i[50];
  assign o[25805] = i[50];
  assign o[25806] = i[50];
  assign o[25807] = i[50];
  assign o[25808] = i[50];
  assign o[25809] = i[50];
  assign o[25810] = i[50];
  assign o[25811] = i[50];
  assign o[25812] = i[50];
  assign o[25813] = i[50];
  assign o[25814] = i[50];
  assign o[25815] = i[50];
  assign o[25816] = i[50];
  assign o[25817] = i[50];
  assign o[25818] = i[50];
  assign o[25819] = i[50];
  assign o[25820] = i[50];
  assign o[25821] = i[50];
  assign o[25822] = i[50];
  assign o[25823] = i[50];
  assign o[25824] = i[50];
  assign o[25825] = i[50];
  assign o[25826] = i[50];
  assign o[25827] = i[50];
  assign o[25828] = i[50];
  assign o[25829] = i[50];
  assign o[25830] = i[50];
  assign o[25831] = i[50];
  assign o[25832] = i[50];
  assign o[25833] = i[50];
  assign o[25834] = i[50];
  assign o[25835] = i[50];
  assign o[25836] = i[50];
  assign o[25837] = i[50];
  assign o[25838] = i[50];
  assign o[25839] = i[50];
  assign o[25840] = i[50];
  assign o[25841] = i[50];
  assign o[25842] = i[50];
  assign o[25843] = i[50];
  assign o[25844] = i[50];
  assign o[25845] = i[50];
  assign o[25846] = i[50];
  assign o[25847] = i[50];
  assign o[25848] = i[50];
  assign o[25849] = i[50];
  assign o[25850] = i[50];
  assign o[25851] = i[50];
  assign o[25852] = i[50];
  assign o[25853] = i[50];
  assign o[25854] = i[50];
  assign o[25855] = i[50];
  assign o[25856] = i[50];
  assign o[25857] = i[50];
  assign o[25858] = i[50];
  assign o[25859] = i[50];
  assign o[25860] = i[50];
  assign o[25861] = i[50];
  assign o[25862] = i[50];
  assign o[25863] = i[50];
  assign o[25864] = i[50];
  assign o[25865] = i[50];
  assign o[25866] = i[50];
  assign o[25867] = i[50];
  assign o[25868] = i[50];
  assign o[25869] = i[50];
  assign o[25870] = i[50];
  assign o[25871] = i[50];
  assign o[25872] = i[50];
  assign o[25873] = i[50];
  assign o[25874] = i[50];
  assign o[25875] = i[50];
  assign o[25876] = i[50];
  assign o[25877] = i[50];
  assign o[25878] = i[50];
  assign o[25879] = i[50];
  assign o[25880] = i[50];
  assign o[25881] = i[50];
  assign o[25882] = i[50];
  assign o[25883] = i[50];
  assign o[25884] = i[50];
  assign o[25885] = i[50];
  assign o[25886] = i[50];
  assign o[25887] = i[50];
  assign o[25888] = i[50];
  assign o[25889] = i[50];
  assign o[25890] = i[50];
  assign o[25891] = i[50];
  assign o[25892] = i[50];
  assign o[25893] = i[50];
  assign o[25894] = i[50];
  assign o[25895] = i[50];
  assign o[25896] = i[50];
  assign o[25897] = i[50];
  assign o[25898] = i[50];
  assign o[25899] = i[50];
  assign o[25900] = i[50];
  assign o[25901] = i[50];
  assign o[25902] = i[50];
  assign o[25903] = i[50];
  assign o[25904] = i[50];
  assign o[25905] = i[50];
  assign o[25906] = i[50];
  assign o[25907] = i[50];
  assign o[25908] = i[50];
  assign o[25909] = i[50];
  assign o[25910] = i[50];
  assign o[25911] = i[50];
  assign o[25912] = i[50];
  assign o[25913] = i[50];
  assign o[25914] = i[50];
  assign o[25915] = i[50];
  assign o[25916] = i[50];
  assign o[25917] = i[50];
  assign o[25918] = i[50];
  assign o[25919] = i[50];
  assign o[25920] = i[50];
  assign o[25921] = i[50];
  assign o[25922] = i[50];
  assign o[25923] = i[50];
  assign o[25924] = i[50];
  assign o[25925] = i[50];
  assign o[25926] = i[50];
  assign o[25927] = i[50];
  assign o[25928] = i[50];
  assign o[25929] = i[50];
  assign o[25930] = i[50];
  assign o[25931] = i[50];
  assign o[25932] = i[50];
  assign o[25933] = i[50];
  assign o[25934] = i[50];
  assign o[25935] = i[50];
  assign o[25936] = i[50];
  assign o[25937] = i[50];
  assign o[25938] = i[50];
  assign o[25939] = i[50];
  assign o[25940] = i[50];
  assign o[25941] = i[50];
  assign o[25942] = i[50];
  assign o[25943] = i[50];
  assign o[25944] = i[50];
  assign o[25945] = i[50];
  assign o[25946] = i[50];
  assign o[25947] = i[50];
  assign o[25948] = i[50];
  assign o[25949] = i[50];
  assign o[25950] = i[50];
  assign o[25951] = i[50];
  assign o[25952] = i[50];
  assign o[25953] = i[50];
  assign o[25954] = i[50];
  assign o[25955] = i[50];
  assign o[25956] = i[50];
  assign o[25957] = i[50];
  assign o[25958] = i[50];
  assign o[25959] = i[50];
  assign o[25960] = i[50];
  assign o[25961] = i[50];
  assign o[25962] = i[50];
  assign o[25963] = i[50];
  assign o[25964] = i[50];
  assign o[25965] = i[50];
  assign o[25966] = i[50];
  assign o[25967] = i[50];
  assign o[25968] = i[50];
  assign o[25969] = i[50];
  assign o[25970] = i[50];
  assign o[25971] = i[50];
  assign o[25972] = i[50];
  assign o[25973] = i[50];
  assign o[25974] = i[50];
  assign o[25975] = i[50];
  assign o[25976] = i[50];
  assign o[25977] = i[50];
  assign o[25978] = i[50];
  assign o[25979] = i[50];
  assign o[25980] = i[50];
  assign o[25981] = i[50];
  assign o[25982] = i[50];
  assign o[25983] = i[50];
  assign o[25984] = i[50];
  assign o[25985] = i[50];
  assign o[25986] = i[50];
  assign o[25987] = i[50];
  assign o[25988] = i[50];
  assign o[25989] = i[50];
  assign o[25990] = i[50];
  assign o[25991] = i[50];
  assign o[25992] = i[50];
  assign o[25993] = i[50];
  assign o[25994] = i[50];
  assign o[25995] = i[50];
  assign o[25996] = i[50];
  assign o[25997] = i[50];
  assign o[25998] = i[50];
  assign o[25999] = i[50];
  assign o[26000] = i[50];
  assign o[26001] = i[50];
  assign o[26002] = i[50];
  assign o[26003] = i[50];
  assign o[26004] = i[50];
  assign o[26005] = i[50];
  assign o[26006] = i[50];
  assign o[26007] = i[50];
  assign o[26008] = i[50];
  assign o[26009] = i[50];
  assign o[26010] = i[50];
  assign o[26011] = i[50];
  assign o[26012] = i[50];
  assign o[26013] = i[50];
  assign o[26014] = i[50];
  assign o[26015] = i[50];
  assign o[26016] = i[50];
  assign o[26017] = i[50];
  assign o[26018] = i[50];
  assign o[26019] = i[50];
  assign o[26020] = i[50];
  assign o[26021] = i[50];
  assign o[26022] = i[50];
  assign o[26023] = i[50];
  assign o[26024] = i[50];
  assign o[26025] = i[50];
  assign o[26026] = i[50];
  assign o[26027] = i[50];
  assign o[26028] = i[50];
  assign o[26029] = i[50];
  assign o[26030] = i[50];
  assign o[26031] = i[50];
  assign o[26032] = i[50];
  assign o[26033] = i[50];
  assign o[26034] = i[50];
  assign o[26035] = i[50];
  assign o[26036] = i[50];
  assign o[26037] = i[50];
  assign o[26038] = i[50];
  assign o[26039] = i[50];
  assign o[26040] = i[50];
  assign o[26041] = i[50];
  assign o[26042] = i[50];
  assign o[26043] = i[50];
  assign o[26044] = i[50];
  assign o[26045] = i[50];
  assign o[26046] = i[50];
  assign o[26047] = i[50];
  assign o[26048] = i[50];
  assign o[26049] = i[50];
  assign o[26050] = i[50];
  assign o[26051] = i[50];
  assign o[26052] = i[50];
  assign o[26053] = i[50];
  assign o[26054] = i[50];
  assign o[26055] = i[50];
  assign o[26056] = i[50];
  assign o[26057] = i[50];
  assign o[26058] = i[50];
  assign o[26059] = i[50];
  assign o[26060] = i[50];
  assign o[26061] = i[50];
  assign o[26062] = i[50];
  assign o[26063] = i[50];
  assign o[26064] = i[50];
  assign o[26065] = i[50];
  assign o[26066] = i[50];
  assign o[26067] = i[50];
  assign o[26068] = i[50];
  assign o[26069] = i[50];
  assign o[26070] = i[50];
  assign o[26071] = i[50];
  assign o[26072] = i[50];
  assign o[26073] = i[50];
  assign o[26074] = i[50];
  assign o[26075] = i[50];
  assign o[26076] = i[50];
  assign o[26077] = i[50];
  assign o[26078] = i[50];
  assign o[26079] = i[50];
  assign o[26080] = i[50];
  assign o[26081] = i[50];
  assign o[26082] = i[50];
  assign o[26083] = i[50];
  assign o[26084] = i[50];
  assign o[26085] = i[50];
  assign o[26086] = i[50];
  assign o[26087] = i[50];
  assign o[26088] = i[50];
  assign o[26089] = i[50];
  assign o[26090] = i[50];
  assign o[26091] = i[50];
  assign o[26092] = i[50];
  assign o[26093] = i[50];
  assign o[26094] = i[50];
  assign o[26095] = i[50];
  assign o[26096] = i[50];
  assign o[26097] = i[50];
  assign o[26098] = i[50];
  assign o[26099] = i[50];
  assign o[26100] = i[50];
  assign o[26101] = i[50];
  assign o[26102] = i[50];
  assign o[26103] = i[50];
  assign o[26104] = i[50];
  assign o[26105] = i[50];
  assign o[26106] = i[50];
  assign o[26107] = i[50];
  assign o[26108] = i[50];
  assign o[26109] = i[50];
  assign o[26110] = i[50];
  assign o[26111] = i[50];
  assign o[25088] = i[49];
  assign o[25089] = i[49];
  assign o[25090] = i[49];
  assign o[25091] = i[49];
  assign o[25092] = i[49];
  assign o[25093] = i[49];
  assign o[25094] = i[49];
  assign o[25095] = i[49];
  assign o[25096] = i[49];
  assign o[25097] = i[49];
  assign o[25098] = i[49];
  assign o[25099] = i[49];
  assign o[25100] = i[49];
  assign o[25101] = i[49];
  assign o[25102] = i[49];
  assign o[25103] = i[49];
  assign o[25104] = i[49];
  assign o[25105] = i[49];
  assign o[25106] = i[49];
  assign o[25107] = i[49];
  assign o[25108] = i[49];
  assign o[25109] = i[49];
  assign o[25110] = i[49];
  assign o[25111] = i[49];
  assign o[25112] = i[49];
  assign o[25113] = i[49];
  assign o[25114] = i[49];
  assign o[25115] = i[49];
  assign o[25116] = i[49];
  assign o[25117] = i[49];
  assign o[25118] = i[49];
  assign o[25119] = i[49];
  assign o[25120] = i[49];
  assign o[25121] = i[49];
  assign o[25122] = i[49];
  assign o[25123] = i[49];
  assign o[25124] = i[49];
  assign o[25125] = i[49];
  assign o[25126] = i[49];
  assign o[25127] = i[49];
  assign o[25128] = i[49];
  assign o[25129] = i[49];
  assign o[25130] = i[49];
  assign o[25131] = i[49];
  assign o[25132] = i[49];
  assign o[25133] = i[49];
  assign o[25134] = i[49];
  assign o[25135] = i[49];
  assign o[25136] = i[49];
  assign o[25137] = i[49];
  assign o[25138] = i[49];
  assign o[25139] = i[49];
  assign o[25140] = i[49];
  assign o[25141] = i[49];
  assign o[25142] = i[49];
  assign o[25143] = i[49];
  assign o[25144] = i[49];
  assign o[25145] = i[49];
  assign o[25146] = i[49];
  assign o[25147] = i[49];
  assign o[25148] = i[49];
  assign o[25149] = i[49];
  assign o[25150] = i[49];
  assign o[25151] = i[49];
  assign o[25152] = i[49];
  assign o[25153] = i[49];
  assign o[25154] = i[49];
  assign o[25155] = i[49];
  assign o[25156] = i[49];
  assign o[25157] = i[49];
  assign o[25158] = i[49];
  assign o[25159] = i[49];
  assign o[25160] = i[49];
  assign o[25161] = i[49];
  assign o[25162] = i[49];
  assign o[25163] = i[49];
  assign o[25164] = i[49];
  assign o[25165] = i[49];
  assign o[25166] = i[49];
  assign o[25167] = i[49];
  assign o[25168] = i[49];
  assign o[25169] = i[49];
  assign o[25170] = i[49];
  assign o[25171] = i[49];
  assign o[25172] = i[49];
  assign o[25173] = i[49];
  assign o[25174] = i[49];
  assign o[25175] = i[49];
  assign o[25176] = i[49];
  assign o[25177] = i[49];
  assign o[25178] = i[49];
  assign o[25179] = i[49];
  assign o[25180] = i[49];
  assign o[25181] = i[49];
  assign o[25182] = i[49];
  assign o[25183] = i[49];
  assign o[25184] = i[49];
  assign o[25185] = i[49];
  assign o[25186] = i[49];
  assign o[25187] = i[49];
  assign o[25188] = i[49];
  assign o[25189] = i[49];
  assign o[25190] = i[49];
  assign o[25191] = i[49];
  assign o[25192] = i[49];
  assign o[25193] = i[49];
  assign o[25194] = i[49];
  assign o[25195] = i[49];
  assign o[25196] = i[49];
  assign o[25197] = i[49];
  assign o[25198] = i[49];
  assign o[25199] = i[49];
  assign o[25200] = i[49];
  assign o[25201] = i[49];
  assign o[25202] = i[49];
  assign o[25203] = i[49];
  assign o[25204] = i[49];
  assign o[25205] = i[49];
  assign o[25206] = i[49];
  assign o[25207] = i[49];
  assign o[25208] = i[49];
  assign o[25209] = i[49];
  assign o[25210] = i[49];
  assign o[25211] = i[49];
  assign o[25212] = i[49];
  assign o[25213] = i[49];
  assign o[25214] = i[49];
  assign o[25215] = i[49];
  assign o[25216] = i[49];
  assign o[25217] = i[49];
  assign o[25218] = i[49];
  assign o[25219] = i[49];
  assign o[25220] = i[49];
  assign o[25221] = i[49];
  assign o[25222] = i[49];
  assign o[25223] = i[49];
  assign o[25224] = i[49];
  assign o[25225] = i[49];
  assign o[25226] = i[49];
  assign o[25227] = i[49];
  assign o[25228] = i[49];
  assign o[25229] = i[49];
  assign o[25230] = i[49];
  assign o[25231] = i[49];
  assign o[25232] = i[49];
  assign o[25233] = i[49];
  assign o[25234] = i[49];
  assign o[25235] = i[49];
  assign o[25236] = i[49];
  assign o[25237] = i[49];
  assign o[25238] = i[49];
  assign o[25239] = i[49];
  assign o[25240] = i[49];
  assign o[25241] = i[49];
  assign o[25242] = i[49];
  assign o[25243] = i[49];
  assign o[25244] = i[49];
  assign o[25245] = i[49];
  assign o[25246] = i[49];
  assign o[25247] = i[49];
  assign o[25248] = i[49];
  assign o[25249] = i[49];
  assign o[25250] = i[49];
  assign o[25251] = i[49];
  assign o[25252] = i[49];
  assign o[25253] = i[49];
  assign o[25254] = i[49];
  assign o[25255] = i[49];
  assign o[25256] = i[49];
  assign o[25257] = i[49];
  assign o[25258] = i[49];
  assign o[25259] = i[49];
  assign o[25260] = i[49];
  assign o[25261] = i[49];
  assign o[25262] = i[49];
  assign o[25263] = i[49];
  assign o[25264] = i[49];
  assign o[25265] = i[49];
  assign o[25266] = i[49];
  assign o[25267] = i[49];
  assign o[25268] = i[49];
  assign o[25269] = i[49];
  assign o[25270] = i[49];
  assign o[25271] = i[49];
  assign o[25272] = i[49];
  assign o[25273] = i[49];
  assign o[25274] = i[49];
  assign o[25275] = i[49];
  assign o[25276] = i[49];
  assign o[25277] = i[49];
  assign o[25278] = i[49];
  assign o[25279] = i[49];
  assign o[25280] = i[49];
  assign o[25281] = i[49];
  assign o[25282] = i[49];
  assign o[25283] = i[49];
  assign o[25284] = i[49];
  assign o[25285] = i[49];
  assign o[25286] = i[49];
  assign o[25287] = i[49];
  assign o[25288] = i[49];
  assign o[25289] = i[49];
  assign o[25290] = i[49];
  assign o[25291] = i[49];
  assign o[25292] = i[49];
  assign o[25293] = i[49];
  assign o[25294] = i[49];
  assign o[25295] = i[49];
  assign o[25296] = i[49];
  assign o[25297] = i[49];
  assign o[25298] = i[49];
  assign o[25299] = i[49];
  assign o[25300] = i[49];
  assign o[25301] = i[49];
  assign o[25302] = i[49];
  assign o[25303] = i[49];
  assign o[25304] = i[49];
  assign o[25305] = i[49];
  assign o[25306] = i[49];
  assign o[25307] = i[49];
  assign o[25308] = i[49];
  assign o[25309] = i[49];
  assign o[25310] = i[49];
  assign o[25311] = i[49];
  assign o[25312] = i[49];
  assign o[25313] = i[49];
  assign o[25314] = i[49];
  assign o[25315] = i[49];
  assign o[25316] = i[49];
  assign o[25317] = i[49];
  assign o[25318] = i[49];
  assign o[25319] = i[49];
  assign o[25320] = i[49];
  assign o[25321] = i[49];
  assign o[25322] = i[49];
  assign o[25323] = i[49];
  assign o[25324] = i[49];
  assign o[25325] = i[49];
  assign o[25326] = i[49];
  assign o[25327] = i[49];
  assign o[25328] = i[49];
  assign o[25329] = i[49];
  assign o[25330] = i[49];
  assign o[25331] = i[49];
  assign o[25332] = i[49];
  assign o[25333] = i[49];
  assign o[25334] = i[49];
  assign o[25335] = i[49];
  assign o[25336] = i[49];
  assign o[25337] = i[49];
  assign o[25338] = i[49];
  assign o[25339] = i[49];
  assign o[25340] = i[49];
  assign o[25341] = i[49];
  assign o[25342] = i[49];
  assign o[25343] = i[49];
  assign o[25344] = i[49];
  assign o[25345] = i[49];
  assign o[25346] = i[49];
  assign o[25347] = i[49];
  assign o[25348] = i[49];
  assign o[25349] = i[49];
  assign o[25350] = i[49];
  assign o[25351] = i[49];
  assign o[25352] = i[49];
  assign o[25353] = i[49];
  assign o[25354] = i[49];
  assign o[25355] = i[49];
  assign o[25356] = i[49];
  assign o[25357] = i[49];
  assign o[25358] = i[49];
  assign o[25359] = i[49];
  assign o[25360] = i[49];
  assign o[25361] = i[49];
  assign o[25362] = i[49];
  assign o[25363] = i[49];
  assign o[25364] = i[49];
  assign o[25365] = i[49];
  assign o[25366] = i[49];
  assign o[25367] = i[49];
  assign o[25368] = i[49];
  assign o[25369] = i[49];
  assign o[25370] = i[49];
  assign o[25371] = i[49];
  assign o[25372] = i[49];
  assign o[25373] = i[49];
  assign o[25374] = i[49];
  assign o[25375] = i[49];
  assign o[25376] = i[49];
  assign o[25377] = i[49];
  assign o[25378] = i[49];
  assign o[25379] = i[49];
  assign o[25380] = i[49];
  assign o[25381] = i[49];
  assign o[25382] = i[49];
  assign o[25383] = i[49];
  assign o[25384] = i[49];
  assign o[25385] = i[49];
  assign o[25386] = i[49];
  assign o[25387] = i[49];
  assign o[25388] = i[49];
  assign o[25389] = i[49];
  assign o[25390] = i[49];
  assign o[25391] = i[49];
  assign o[25392] = i[49];
  assign o[25393] = i[49];
  assign o[25394] = i[49];
  assign o[25395] = i[49];
  assign o[25396] = i[49];
  assign o[25397] = i[49];
  assign o[25398] = i[49];
  assign o[25399] = i[49];
  assign o[25400] = i[49];
  assign o[25401] = i[49];
  assign o[25402] = i[49];
  assign o[25403] = i[49];
  assign o[25404] = i[49];
  assign o[25405] = i[49];
  assign o[25406] = i[49];
  assign o[25407] = i[49];
  assign o[25408] = i[49];
  assign o[25409] = i[49];
  assign o[25410] = i[49];
  assign o[25411] = i[49];
  assign o[25412] = i[49];
  assign o[25413] = i[49];
  assign o[25414] = i[49];
  assign o[25415] = i[49];
  assign o[25416] = i[49];
  assign o[25417] = i[49];
  assign o[25418] = i[49];
  assign o[25419] = i[49];
  assign o[25420] = i[49];
  assign o[25421] = i[49];
  assign o[25422] = i[49];
  assign o[25423] = i[49];
  assign o[25424] = i[49];
  assign o[25425] = i[49];
  assign o[25426] = i[49];
  assign o[25427] = i[49];
  assign o[25428] = i[49];
  assign o[25429] = i[49];
  assign o[25430] = i[49];
  assign o[25431] = i[49];
  assign o[25432] = i[49];
  assign o[25433] = i[49];
  assign o[25434] = i[49];
  assign o[25435] = i[49];
  assign o[25436] = i[49];
  assign o[25437] = i[49];
  assign o[25438] = i[49];
  assign o[25439] = i[49];
  assign o[25440] = i[49];
  assign o[25441] = i[49];
  assign o[25442] = i[49];
  assign o[25443] = i[49];
  assign o[25444] = i[49];
  assign o[25445] = i[49];
  assign o[25446] = i[49];
  assign o[25447] = i[49];
  assign o[25448] = i[49];
  assign o[25449] = i[49];
  assign o[25450] = i[49];
  assign o[25451] = i[49];
  assign o[25452] = i[49];
  assign o[25453] = i[49];
  assign o[25454] = i[49];
  assign o[25455] = i[49];
  assign o[25456] = i[49];
  assign o[25457] = i[49];
  assign o[25458] = i[49];
  assign o[25459] = i[49];
  assign o[25460] = i[49];
  assign o[25461] = i[49];
  assign o[25462] = i[49];
  assign o[25463] = i[49];
  assign o[25464] = i[49];
  assign o[25465] = i[49];
  assign o[25466] = i[49];
  assign o[25467] = i[49];
  assign o[25468] = i[49];
  assign o[25469] = i[49];
  assign o[25470] = i[49];
  assign o[25471] = i[49];
  assign o[25472] = i[49];
  assign o[25473] = i[49];
  assign o[25474] = i[49];
  assign o[25475] = i[49];
  assign o[25476] = i[49];
  assign o[25477] = i[49];
  assign o[25478] = i[49];
  assign o[25479] = i[49];
  assign o[25480] = i[49];
  assign o[25481] = i[49];
  assign o[25482] = i[49];
  assign o[25483] = i[49];
  assign o[25484] = i[49];
  assign o[25485] = i[49];
  assign o[25486] = i[49];
  assign o[25487] = i[49];
  assign o[25488] = i[49];
  assign o[25489] = i[49];
  assign o[25490] = i[49];
  assign o[25491] = i[49];
  assign o[25492] = i[49];
  assign o[25493] = i[49];
  assign o[25494] = i[49];
  assign o[25495] = i[49];
  assign o[25496] = i[49];
  assign o[25497] = i[49];
  assign o[25498] = i[49];
  assign o[25499] = i[49];
  assign o[25500] = i[49];
  assign o[25501] = i[49];
  assign o[25502] = i[49];
  assign o[25503] = i[49];
  assign o[25504] = i[49];
  assign o[25505] = i[49];
  assign o[25506] = i[49];
  assign o[25507] = i[49];
  assign o[25508] = i[49];
  assign o[25509] = i[49];
  assign o[25510] = i[49];
  assign o[25511] = i[49];
  assign o[25512] = i[49];
  assign o[25513] = i[49];
  assign o[25514] = i[49];
  assign o[25515] = i[49];
  assign o[25516] = i[49];
  assign o[25517] = i[49];
  assign o[25518] = i[49];
  assign o[25519] = i[49];
  assign o[25520] = i[49];
  assign o[25521] = i[49];
  assign o[25522] = i[49];
  assign o[25523] = i[49];
  assign o[25524] = i[49];
  assign o[25525] = i[49];
  assign o[25526] = i[49];
  assign o[25527] = i[49];
  assign o[25528] = i[49];
  assign o[25529] = i[49];
  assign o[25530] = i[49];
  assign o[25531] = i[49];
  assign o[25532] = i[49];
  assign o[25533] = i[49];
  assign o[25534] = i[49];
  assign o[25535] = i[49];
  assign o[25536] = i[49];
  assign o[25537] = i[49];
  assign o[25538] = i[49];
  assign o[25539] = i[49];
  assign o[25540] = i[49];
  assign o[25541] = i[49];
  assign o[25542] = i[49];
  assign o[25543] = i[49];
  assign o[25544] = i[49];
  assign o[25545] = i[49];
  assign o[25546] = i[49];
  assign o[25547] = i[49];
  assign o[25548] = i[49];
  assign o[25549] = i[49];
  assign o[25550] = i[49];
  assign o[25551] = i[49];
  assign o[25552] = i[49];
  assign o[25553] = i[49];
  assign o[25554] = i[49];
  assign o[25555] = i[49];
  assign o[25556] = i[49];
  assign o[25557] = i[49];
  assign o[25558] = i[49];
  assign o[25559] = i[49];
  assign o[25560] = i[49];
  assign o[25561] = i[49];
  assign o[25562] = i[49];
  assign o[25563] = i[49];
  assign o[25564] = i[49];
  assign o[25565] = i[49];
  assign o[25566] = i[49];
  assign o[25567] = i[49];
  assign o[25568] = i[49];
  assign o[25569] = i[49];
  assign o[25570] = i[49];
  assign o[25571] = i[49];
  assign o[25572] = i[49];
  assign o[25573] = i[49];
  assign o[25574] = i[49];
  assign o[25575] = i[49];
  assign o[25576] = i[49];
  assign o[25577] = i[49];
  assign o[25578] = i[49];
  assign o[25579] = i[49];
  assign o[25580] = i[49];
  assign o[25581] = i[49];
  assign o[25582] = i[49];
  assign o[25583] = i[49];
  assign o[25584] = i[49];
  assign o[25585] = i[49];
  assign o[25586] = i[49];
  assign o[25587] = i[49];
  assign o[25588] = i[49];
  assign o[25589] = i[49];
  assign o[25590] = i[49];
  assign o[25591] = i[49];
  assign o[25592] = i[49];
  assign o[25593] = i[49];
  assign o[25594] = i[49];
  assign o[25595] = i[49];
  assign o[25596] = i[49];
  assign o[25597] = i[49];
  assign o[25598] = i[49];
  assign o[25599] = i[49];
  assign o[24576] = i[48];
  assign o[24577] = i[48];
  assign o[24578] = i[48];
  assign o[24579] = i[48];
  assign o[24580] = i[48];
  assign o[24581] = i[48];
  assign o[24582] = i[48];
  assign o[24583] = i[48];
  assign o[24584] = i[48];
  assign o[24585] = i[48];
  assign o[24586] = i[48];
  assign o[24587] = i[48];
  assign o[24588] = i[48];
  assign o[24589] = i[48];
  assign o[24590] = i[48];
  assign o[24591] = i[48];
  assign o[24592] = i[48];
  assign o[24593] = i[48];
  assign o[24594] = i[48];
  assign o[24595] = i[48];
  assign o[24596] = i[48];
  assign o[24597] = i[48];
  assign o[24598] = i[48];
  assign o[24599] = i[48];
  assign o[24600] = i[48];
  assign o[24601] = i[48];
  assign o[24602] = i[48];
  assign o[24603] = i[48];
  assign o[24604] = i[48];
  assign o[24605] = i[48];
  assign o[24606] = i[48];
  assign o[24607] = i[48];
  assign o[24608] = i[48];
  assign o[24609] = i[48];
  assign o[24610] = i[48];
  assign o[24611] = i[48];
  assign o[24612] = i[48];
  assign o[24613] = i[48];
  assign o[24614] = i[48];
  assign o[24615] = i[48];
  assign o[24616] = i[48];
  assign o[24617] = i[48];
  assign o[24618] = i[48];
  assign o[24619] = i[48];
  assign o[24620] = i[48];
  assign o[24621] = i[48];
  assign o[24622] = i[48];
  assign o[24623] = i[48];
  assign o[24624] = i[48];
  assign o[24625] = i[48];
  assign o[24626] = i[48];
  assign o[24627] = i[48];
  assign o[24628] = i[48];
  assign o[24629] = i[48];
  assign o[24630] = i[48];
  assign o[24631] = i[48];
  assign o[24632] = i[48];
  assign o[24633] = i[48];
  assign o[24634] = i[48];
  assign o[24635] = i[48];
  assign o[24636] = i[48];
  assign o[24637] = i[48];
  assign o[24638] = i[48];
  assign o[24639] = i[48];
  assign o[24640] = i[48];
  assign o[24641] = i[48];
  assign o[24642] = i[48];
  assign o[24643] = i[48];
  assign o[24644] = i[48];
  assign o[24645] = i[48];
  assign o[24646] = i[48];
  assign o[24647] = i[48];
  assign o[24648] = i[48];
  assign o[24649] = i[48];
  assign o[24650] = i[48];
  assign o[24651] = i[48];
  assign o[24652] = i[48];
  assign o[24653] = i[48];
  assign o[24654] = i[48];
  assign o[24655] = i[48];
  assign o[24656] = i[48];
  assign o[24657] = i[48];
  assign o[24658] = i[48];
  assign o[24659] = i[48];
  assign o[24660] = i[48];
  assign o[24661] = i[48];
  assign o[24662] = i[48];
  assign o[24663] = i[48];
  assign o[24664] = i[48];
  assign o[24665] = i[48];
  assign o[24666] = i[48];
  assign o[24667] = i[48];
  assign o[24668] = i[48];
  assign o[24669] = i[48];
  assign o[24670] = i[48];
  assign o[24671] = i[48];
  assign o[24672] = i[48];
  assign o[24673] = i[48];
  assign o[24674] = i[48];
  assign o[24675] = i[48];
  assign o[24676] = i[48];
  assign o[24677] = i[48];
  assign o[24678] = i[48];
  assign o[24679] = i[48];
  assign o[24680] = i[48];
  assign o[24681] = i[48];
  assign o[24682] = i[48];
  assign o[24683] = i[48];
  assign o[24684] = i[48];
  assign o[24685] = i[48];
  assign o[24686] = i[48];
  assign o[24687] = i[48];
  assign o[24688] = i[48];
  assign o[24689] = i[48];
  assign o[24690] = i[48];
  assign o[24691] = i[48];
  assign o[24692] = i[48];
  assign o[24693] = i[48];
  assign o[24694] = i[48];
  assign o[24695] = i[48];
  assign o[24696] = i[48];
  assign o[24697] = i[48];
  assign o[24698] = i[48];
  assign o[24699] = i[48];
  assign o[24700] = i[48];
  assign o[24701] = i[48];
  assign o[24702] = i[48];
  assign o[24703] = i[48];
  assign o[24704] = i[48];
  assign o[24705] = i[48];
  assign o[24706] = i[48];
  assign o[24707] = i[48];
  assign o[24708] = i[48];
  assign o[24709] = i[48];
  assign o[24710] = i[48];
  assign o[24711] = i[48];
  assign o[24712] = i[48];
  assign o[24713] = i[48];
  assign o[24714] = i[48];
  assign o[24715] = i[48];
  assign o[24716] = i[48];
  assign o[24717] = i[48];
  assign o[24718] = i[48];
  assign o[24719] = i[48];
  assign o[24720] = i[48];
  assign o[24721] = i[48];
  assign o[24722] = i[48];
  assign o[24723] = i[48];
  assign o[24724] = i[48];
  assign o[24725] = i[48];
  assign o[24726] = i[48];
  assign o[24727] = i[48];
  assign o[24728] = i[48];
  assign o[24729] = i[48];
  assign o[24730] = i[48];
  assign o[24731] = i[48];
  assign o[24732] = i[48];
  assign o[24733] = i[48];
  assign o[24734] = i[48];
  assign o[24735] = i[48];
  assign o[24736] = i[48];
  assign o[24737] = i[48];
  assign o[24738] = i[48];
  assign o[24739] = i[48];
  assign o[24740] = i[48];
  assign o[24741] = i[48];
  assign o[24742] = i[48];
  assign o[24743] = i[48];
  assign o[24744] = i[48];
  assign o[24745] = i[48];
  assign o[24746] = i[48];
  assign o[24747] = i[48];
  assign o[24748] = i[48];
  assign o[24749] = i[48];
  assign o[24750] = i[48];
  assign o[24751] = i[48];
  assign o[24752] = i[48];
  assign o[24753] = i[48];
  assign o[24754] = i[48];
  assign o[24755] = i[48];
  assign o[24756] = i[48];
  assign o[24757] = i[48];
  assign o[24758] = i[48];
  assign o[24759] = i[48];
  assign o[24760] = i[48];
  assign o[24761] = i[48];
  assign o[24762] = i[48];
  assign o[24763] = i[48];
  assign o[24764] = i[48];
  assign o[24765] = i[48];
  assign o[24766] = i[48];
  assign o[24767] = i[48];
  assign o[24768] = i[48];
  assign o[24769] = i[48];
  assign o[24770] = i[48];
  assign o[24771] = i[48];
  assign o[24772] = i[48];
  assign o[24773] = i[48];
  assign o[24774] = i[48];
  assign o[24775] = i[48];
  assign o[24776] = i[48];
  assign o[24777] = i[48];
  assign o[24778] = i[48];
  assign o[24779] = i[48];
  assign o[24780] = i[48];
  assign o[24781] = i[48];
  assign o[24782] = i[48];
  assign o[24783] = i[48];
  assign o[24784] = i[48];
  assign o[24785] = i[48];
  assign o[24786] = i[48];
  assign o[24787] = i[48];
  assign o[24788] = i[48];
  assign o[24789] = i[48];
  assign o[24790] = i[48];
  assign o[24791] = i[48];
  assign o[24792] = i[48];
  assign o[24793] = i[48];
  assign o[24794] = i[48];
  assign o[24795] = i[48];
  assign o[24796] = i[48];
  assign o[24797] = i[48];
  assign o[24798] = i[48];
  assign o[24799] = i[48];
  assign o[24800] = i[48];
  assign o[24801] = i[48];
  assign o[24802] = i[48];
  assign o[24803] = i[48];
  assign o[24804] = i[48];
  assign o[24805] = i[48];
  assign o[24806] = i[48];
  assign o[24807] = i[48];
  assign o[24808] = i[48];
  assign o[24809] = i[48];
  assign o[24810] = i[48];
  assign o[24811] = i[48];
  assign o[24812] = i[48];
  assign o[24813] = i[48];
  assign o[24814] = i[48];
  assign o[24815] = i[48];
  assign o[24816] = i[48];
  assign o[24817] = i[48];
  assign o[24818] = i[48];
  assign o[24819] = i[48];
  assign o[24820] = i[48];
  assign o[24821] = i[48];
  assign o[24822] = i[48];
  assign o[24823] = i[48];
  assign o[24824] = i[48];
  assign o[24825] = i[48];
  assign o[24826] = i[48];
  assign o[24827] = i[48];
  assign o[24828] = i[48];
  assign o[24829] = i[48];
  assign o[24830] = i[48];
  assign o[24831] = i[48];
  assign o[24832] = i[48];
  assign o[24833] = i[48];
  assign o[24834] = i[48];
  assign o[24835] = i[48];
  assign o[24836] = i[48];
  assign o[24837] = i[48];
  assign o[24838] = i[48];
  assign o[24839] = i[48];
  assign o[24840] = i[48];
  assign o[24841] = i[48];
  assign o[24842] = i[48];
  assign o[24843] = i[48];
  assign o[24844] = i[48];
  assign o[24845] = i[48];
  assign o[24846] = i[48];
  assign o[24847] = i[48];
  assign o[24848] = i[48];
  assign o[24849] = i[48];
  assign o[24850] = i[48];
  assign o[24851] = i[48];
  assign o[24852] = i[48];
  assign o[24853] = i[48];
  assign o[24854] = i[48];
  assign o[24855] = i[48];
  assign o[24856] = i[48];
  assign o[24857] = i[48];
  assign o[24858] = i[48];
  assign o[24859] = i[48];
  assign o[24860] = i[48];
  assign o[24861] = i[48];
  assign o[24862] = i[48];
  assign o[24863] = i[48];
  assign o[24864] = i[48];
  assign o[24865] = i[48];
  assign o[24866] = i[48];
  assign o[24867] = i[48];
  assign o[24868] = i[48];
  assign o[24869] = i[48];
  assign o[24870] = i[48];
  assign o[24871] = i[48];
  assign o[24872] = i[48];
  assign o[24873] = i[48];
  assign o[24874] = i[48];
  assign o[24875] = i[48];
  assign o[24876] = i[48];
  assign o[24877] = i[48];
  assign o[24878] = i[48];
  assign o[24879] = i[48];
  assign o[24880] = i[48];
  assign o[24881] = i[48];
  assign o[24882] = i[48];
  assign o[24883] = i[48];
  assign o[24884] = i[48];
  assign o[24885] = i[48];
  assign o[24886] = i[48];
  assign o[24887] = i[48];
  assign o[24888] = i[48];
  assign o[24889] = i[48];
  assign o[24890] = i[48];
  assign o[24891] = i[48];
  assign o[24892] = i[48];
  assign o[24893] = i[48];
  assign o[24894] = i[48];
  assign o[24895] = i[48];
  assign o[24896] = i[48];
  assign o[24897] = i[48];
  assign o[24898] = i[48];
  assign o[24899] = i[48];
  assign o[24900] = i[48];
  assign o[24901] = i[48];
  assign o[24902] = i[48];
  assign o[24903] = i[48];
  assign o[24904] = i[48];
  assign o[24905] = i[48];
  assign o[24906] = i[48];
  assign o[24907] = i[48];
  assign o[24908] = i[48];
  assign o[24909] = i[48];
  assign o[24910] = i[48];
  assign o[24911] = i[48];
  assign o[24912] = i[48];
  assign o[24913] = i[48];
  assign o[24914] = i[48];
  assign o[24915] = i[48];
  assign o[24916] = i[48];
  assign o[24917] = i[48];
  assign o[24918] = i[48];
  assign o[24919] = i[48];
  assign o[24920] = i[48];
  assign o[24921] = i[48];
  assign o[24922] = i[48];
  assign o[24923] = i[48];
  assign o[24924] = i[48];
  assign o[24925] = i[48];
  assign o[24926] = i[48];
  assign o[24927] = i[48];
  assign o[24928] = i[48];
  assign o[24929] = i[48];
  assign o[24930] = i[48];
  assign o[24931] = i[48];
  assign o[24932] = i[48];
  assign o[24933] = i[48];
  assign o[24934] = i[48];
  assign o[24935] = i[48];
  assign o[24936] = i[48];
  assign o[24937] = i[48];
  assign o[24938] = i[48];
  assign o[24939] = i[48];
  assign o[24940] = i[48];
  assign o[24941] = i[48];
  assign o[24942] = i[48];
  assign o[24943] = i[48];
  assign o[24944] = i[48];
  assign o[24945] = i[48];
  assign o[24946] = i[48];
  assign o[24947] = i[48];
  assign o[24948] = i[48];
  assign o[24949] = i[48];
  assign o[24950] = i[48];
  assign o[24951] = i[48];
  assign o[24952] = i[48];
  assign o[24953] = i[48];
  assign o[24954] = i[48];
  assign o[24955] = i[48];
  assign o[24956] = i[48];
  assign o[24957] = i[48];
  assign o[24958] = i[48];
  assign o[24959] = i[48];
  assign o[24960] = i[48];
  assign o[24961] = i[48];
  assign o[24962] = i[48];
  assign o[24963] = i[48];
  assign o[24964] = i[48];
  assign o[24965] = i[48];
  assign o[24966] = i[48];
  assign o[24967] = i[48];
  assign o[24968] = i[48];
  assign o[24969] = i[48];
  assign o[24970] = i[48];
  assign o[24971] = i[48];
  assign o[24972] = i[48];
  assign o[24973] = i[48];
  assign o[24974] = i[48];
  assign o[24975] = i[48];
  assign o[24976] = i[48];
  assign o[24977] = i[48];
  assign o[24978] = i[48];
  assign o[24979] = i[48];
  assign o[24980] = i[48];
  assign o[24981] = i[48];
  assign o[24982] = i[48];
  assign o[24983] = i[48];
  assign o[24984] = i[48];
  assign o[24985] = i[48];
  assign o[24986] = i[48];
  assign o[24987] = i[48];
  assign o[24988] = i[48];
  assign o[24989] = i[48];
  assign o[24990] = i[48];
  assign o[24991] = i[48];
  assign o[24992] = i[48];
  assign o[24993] = i[48];
  assign o[24994] = i[48];
  assign o[24995] = i[48];
  assign o[24996] = i[48];
  assign o[24997] = i[48];
  assign o[24998] = i[48];
  assign o[24999] = i[48];
  assign o[25000] = i[48];
  assign o[25001] = i[48];
  assign o[25002] = i[48];
  assign o[25003] = i[48];
  assign o[25004] = i[48];
  assign o[25005] = i[48];
  assign o[25006] = i[48];
  assign o[25007] = i[48];
  assign o[25008] = i[48];
  assign o[25009] = i[48];
  assign o[25010] = i[48];
  assign o[25011] = i[48];
  assign o[25012] = i[48];
  assign o[25013] = i[48];
  assign o[25014] = i[48];
  assign o[25015] = i[48];
  assign o[25016] = i[48];
  assign o[25017] = i[48];
  assign o[25018] = i[48];
  assign o[25019] = i[48];
  assign o[25020] = i[48];
  assign o[25021] = i[48];
  assign o[25022] = i[48];
  assign o[25023] = i[48];
  assign o[25024] = i[48];
  assign o[25025] = i[48];
  assign o[25026] = i[48];
  assign o[25027] = i[48];
  assign o[25028] = i[48];
  assign o[25029] = i[48];
  assign o[25030] = i[48];
  assign o[25031] = i[48];
  assign o[25032] = i[48];
  assign o[25033] = i[48];
  assign o[25034] = i[48];
  assign o[25035] = i[48];
  assign o[25036] = i[48];
  assign o[25037] = i[48];
  assign o[25038] = i[48];
  assign o[25039] = i[48];
  assign o[25040] = i[48];
  assign o[25041] = i[48];
  assign o[25042] = i[48];
  assign o[25043] = i[48];
  assign o[25044] = i[48];
  assign o[25045] = i[48];
  assign o[25046] = i[48];
  assign o[25047] = i[48];
  assign o[25048] = i[48];
  assign o[25049] = i[48];
  assign o[25050] = i[48];
  assign o[25051] = i[48];
  assign o[25052] = i[48];
  assign o[25053] = i[48];
  assign o[25054] = i[48];
  assign o[25055] = i[48];
  assign o[25056] = i[48];
  assign o[25057] = i[48];
  assign o[25058] = i[48];
  assign o[25059] = i[48];
  assign o[25060] = i[48];
  assign o[25061] = i[48];
  assign o[25062] = i[48];
  assign o[25063] = i[48];
  assign o[25064] = i[48];
  assign o[25065] = i[48];
  assign o[25066] = i[48];
  assign o[25067] = i[48];
  assign o[25068] = i[48];
  assign o[25069] = i[48];
  assign o[25070] = i[48];
  assign o[25071] = i[48];
  assign o[25072] = i[48];
  assign o[25073] = i[48];
  assign o[25074] = i[48];
  assign o[25075] = i[48];
  assign o[25076] = i[48];
  assign o[25077] = i[48];
  assign o[25078] = i[48];
  assign o[25079] = i[48];
  assign o[25080] = i[48];
  assign o[25081] = i[48];
  assign o[25082] = i[48];
  assign o[25083] = i[48];
  assign o[25084] = i[48];
  assign o[25085] = i[48];
  assign o[25086] = i[48];
  assign o[25087] = i[48];
  assign o[24064] = i[47];
  assign o[24065] = i[47];
  assign o[24066] = i[47];
  assign o[24067] = i[47];
  assign o[24068] = i[47];
  assign o[24069] = i[47];
  assign o[24070] = i[47];
  assign o[24071] = i[47];
  assign o[24072] = i[47];
  assign o[24073] = i[47];
  assign o[24074] = i[47];
  assign o[24075] = i[47];
  assign o[24076] = i[47];
  assign o[24077] = i[47];
  assign o[24078] = i[47];
  assign o[24079] = i[47];
  assign o[24080] = i[47];
  assign o[24081] = i[47];
  assign o[24082] = i[47];
  assign o[24083] = i[47];
  assign o[24084] = i[47];
  assign o[24085] = i[47];
  assign o[24086] = i[47];
  assign o[24087] = i[47];
  assign o[24088] = i[47];
  assign o[24089] = i[47];
  assign o[24090] = i[47];
  assign o[24091] = i[47];
  assign o[24092] = i[47];
  assign o[24093] = i[47];
  assign o[24094] = i[47];
  assign o[24095] = i[47];
  assign o[24096] = i[47];
  assign o[24097] = i[47];
  assign o[24098] = i[47];
  assign o[24099] = i[47];
  assign o[24100] = i[47];
  assign o[24101] = i[47];
  assign o[24102] = i[47];
  assign o[24103] = i[47];
  assign o[24104] = i[47];
  assign o[24105] = i[47];
  assign o[24106] = i[47];
  assign o[24107] = i[47];
  assign o[24108] = i[47];
  assign o[24109] = i[47];
  assign o[24110] = i[47];
  assign o[24111] = i[47];
  assign o[24112] = i[47];
  assign o[24113] = i[47];
  assign o[24114] = i[47];
  assign o[24115] = i[47];
  assign o[24116] = i[47];
  assign o[24117] = i[47];
  assign o[24118] = i[47];
  assign o[24119] = i[47];
  assign o[24120] = i[47];
  assign o[24121] = i[47];
  assign o[24122] = i[47];
  assign o[24123] = i[47];
  assign o[24124] = i[47];
  assign o[24125] = i[47];
  assign o[24126] = i[47];
  assign o[24127] = i[47];
  assign o[24128] = i[47];
  assign o[24129] = i[47];
  assign o[24130] = i[47];
  assign o[24131] = i[47];
  assign o[24132] = i[47];
  assign o[24133] = i[47];
  assign o[24134] = i[47];
  assign o[24135] = i[47];
  assign o[24136] = i[47];
  assign o[24137] = i[47];
  assign o[24138] = i[47];
  assign o[24139] = i[47];
  assign o[24140] = i[47];
  assign o[24141] = i[47];
  assign o[24142] = i[47];
  assign o[24143] = i[47];
  assign o[24144] = i[47];
  assign o[24145] = i[47];
  assign o[24146] = i[47];
  assign o[24147] = i[47];
  assign o[24148] = i[47];
  assign o[24149] = i[47];
  assign o[24150] = i[47];
  assign o[24151] = i[47];
  assign o[24152] = i[47];
  assign o[24153] = i[47];
  assign o[24154] = i[47];
  assign o[24155] = i[47];
  assign o[24156] = i[47];
  assign o[24157] = i[47];
  assign o[24158] = i[47];
  assign o[24159] = i[47];
  assign o[24160] = i[47];
  assign o[24161] = i[47];
  assign o[24162] = i[47];
  assign o[24163] = i[47];
  assign o[24164] = i[47];
  assign o[24165] = i[47];
  assign o[24166] = i[47];
  assign o[24167] = i[47];
  assign o[24168] = i[47];
  assign o[24169] = i[47];
  assign o[24170] = i[47];
  assign o[24171] = i[47];
  assign o[24172] = i[47];
  assign o[24173] = i[47];
  assign o[24174] = i[47];
  assign o[24175] = i[47];
  assign o[24176] = i[47];
  assign o[24177] = i[47];
  assign o[24178] = i[47];
  assign o[24179] = i[47];
  assign o[24180] = i[47];
  assign o[24181] = i[47];
  assign o[24182] = i[47];
  assign o[24183] = i[47];
  assign o[24184] = i[47];
  assign o[24185] = i[47];
  assign o[24186] = i[47];
  assign o[24187] = i[47];
  assign o[24188] = i[47];
  assign o[24189] = i[47];
  assign o[24190] = i[47];
  assign o[24191] = i[47];
  assign o[24192] = i[47];
  assign o[24193] = i[47];
  assign o[24194] = i[47];
  assign o[24195] = i[47];
  assign o[24196] = i[47];
  assign o[24197] = i[47];
  assign o[24198] = i[47];
  assign o[24199] = i[47];
  assign o[24200] = i[47];
  assign o[24201] = i[47];
  assign o[24202] = i[47];
  assign o[24203] = i[47];
  assign o[24204] = i[47];
  assign o[24205] = i[47];
  assign o[24206] = i[47];
  assign o[24207] = i[47];
  assign o[24208] = i[47];
  assign o[24209] = i[47];
  assign o[24210] = i[47];
  assign o[24211] = i[47];
  assign o[24212] = i[47];
  assign o[24213] = i[47];
  assign o[24214] = i[47];
  assign o[24215] = i[47];
  assign o[24216] = i[47];
  assign o[24217] = i[47];
  assign o[24218] = i[47];
  assign o[24219] = i[47];
  assign o[24220] = i[47];
  assign o[24221] = i[47];
  assign o[24222] = i[47];
  assign o[24223] = i[47];
  assign o[24224] = i[47];
  assign o[24225] = i[47];
  assign o[24226] = i[47];
  assign o[24227] = i[47];
  assign o[24228] = i[47];
  assign o[24229] = i[47];
  assign o[24230] = i[47];
  assign o[24231] = i[47];
  assign o[24232] = i[47];
  assign o[24233] = i[47];
  assign o[24234] = i[47];
  assign o[24235] = i[47];
  assign o[24236] = i[47];
  assign o[24237] = i[47];
  assign o[24238] = i[47];
  assign o[24239] = i[47];
  assign o[24240] = i[47];
  assign o[24241] = i[47];
  assign o[24242] = i[47];
  assign o[24243] = i[47];
  assign o[24244] = i[47];
  assign o[24245] = i[47];
  assign o[24246] = i[47];
  assign o[24247] = i[47];
  assign o[24248] = i[47];
  assign o[24249] = i[47];
  assign o[24250] = i[47];
  assign o[24251] = i[47];
  assign o[24252] = i[47];
  assign o[24253] = i[47];
  assign o[24254] = i[47];
  assign o[24255] = i[47];
  assign o[24256] = i[47];
  assign o[24257] = i[47];
  assign o[24258] = i[47];
  assign o[24259] = i[47];
  assign o[24260] = i[47];
  assign o[24261] = i[47];
  assign o[24262] = i[47];
  assign o[24263] = i[47];
  assign o[24264] = i[47];
  assign o[24265] = i[47];
  assign o[24266] = i[47];
  assign o[24267] = i[47];
  assign o[24268] = i[47];
  assign o[24269] = i[47];
  assign o[24270] = i[47];
  assign o[24271] = i[47];
  assign o[24272] = i[47];
  assign o[24273] = i[47];
  assign o[24274] = i[47];
  assign o[24275] = i[47];
  assign o[24276] = i[47];
  assign o[24277] = i[47];
  assign o[24278] = i[47];
  assign o[24279] = i[47];
  assign o[24280] = i[47];
  assign o[24281] = i[47];
  assign o[24282] = i[47];
  assign o[24283] = i[47];
  assign o[24284] = i[47];
  assign o[24285] = i[47];
  assign o[24286] = i[47];
  assign o[24287] = i[47];
  assign o[24288] = i[47];
  assign o[24289] = i[47];
  assign o[24290] = i[47];
  assign o[24291] = i[47];
  assign o[24292] = i[47];
  assign o[24293] = i[47];
  assign o[24294] = i[47];
  assign o[24295] = i[47];
  assign o[24296] = i[47];
  assign o[24297] = i[47];
  assign o[24298] = i[47];
  assign o[24299] = i[47];
  assign o[24300] = i[47];
  assign o[24301] = i[47];
  assign o[24302] = i[47];
  assign o[24303] = i[47];
  assign o[24304] = i[47];
  assign o[24305] = i[47];
  assign o[24306] = i[47];
  assign o[24307] = i[47];
  assign o[24308] = i[47];
  assign o[24309] = i[47];
  assign o[24310] = i[47];
  assign o[24311] = i[47];
  assign o[24312] = i[47];
  assign o[24313] = i[47];
  assign o[24314] = i[47];
  assign o[24315] = i[47];
  assign o[24316] = i[47];
  assign o[24317] = i[47];
  assign o[24318] = i[47];
  assign o[24319] = i[47];
  assign o[24320] = i[47];
  assign o[24321] = i[47];
  assign o[24322] = i[47];
  assign o[24323] = i[47];
  assign o[24324] = i[47];
  assign o[24325] = i[47];
  assign o[24326] = i[47];
  assign o[24327] = i[47];
  assign o[24328] = i[47];
  assign o[24329] = i[47];
  assign o[24330] = i[47];
  assign o[24331] = i[47];
  assign o[24332] = i[47];
  assign o[24333] = i[47];
  assign o[24334] = i[47];
  assign o[24335] = i[47];
  assign o[24336] = i[47];
  assign o[24337] = i[47];
  assign o[24338] = i[47];
  assign o[24339] = i[47];
  assign o[24340] = i[47];
  assign o[24341] = i[47];
  assign o[24342] = i[47];
  assign o[24343] = i[47];
  assign o[24344] = i[47];
  assign o[24345] = i[47];
  assign o[24346] = i[47];
  assign o[24347] = i[47];
  assign o[24348] = i[47];
  assign o[24349] = i[47];
  assign o[24350] = i[47];
  assign o[24351] = i[47];
  assign o[24352] = i[47];
  assign o[24353] = i[47];
  assign o[24354] = i[47];
  assign o[24355] = i[47];
  assign o[24356] = i[47];
  assign o[24357] = i[47];
  assign o[24358] = i[47];
  assign o[24359] = i[47];
  assign o[24360] = i[47];
  assign o[24361] = i[47];
  assign o[24362] = i[47];
  assign o[24363] = i[47];
  assign o[24364] = i[47];
  assign o[24365] = i[47];
  assign o[24366] = i[47];
  assign o[24367] = i[47];
  assign o[24368] = i[47];
  assign o[24369] = i[47];
  assign o[24370] = i[47];
  assign o[24371] = i[47];
  assign o[24372] = i[47];
  assign o[24373] = i[47];
  assign o[24374] = i[47];
  assign o[24375] = i[47];
  assign o[24376] = i[47];
  assign o[24377] = i[47];
  assign o[24378] = i[47];
  assign o[24379] = i[47];
  assign o[24380] = i[47];
  assign o[24381] = i[47];
  assign o[24382] = i[47];
  assign o[24383] = i[47];
  assign o[24384] = i[47];
  assign o[24385] = i[47];
  assign o[24386] = i[47];
  assign o[24387] = i[47];
  assign o[24388] = i[47];
  assign o[24389] = i[47];
  assign o[24390] = i[47];
  assign o[24391] = i[47];
  assign o[24392] = i[47];
  assign o[24393] = i[47];
  assign o[24394] = i[47];
  assign o[24395] = i[47];
  assign o[24396] = i[47];
  assign o[24397] = i[47];
  assign o[24398] = i[47];
  assign o[24399] = i[47];
  assign o[24400] = i[47];
  assign o[24401] = i[47];
  assign o[24402] = i[47];
  assign o[24403] = i[47];
  assign o[24404] = i[47];
  assign o[24405] = i[47];
  assign o[24406] = i[47];
  assign o[24407] = i[47];
  assign o[24408] = i[47];
  assign o[24409] = i[47];
  assign o[24410] = i[47];
  assign o[24411] = i[47];
  assign o[24412] = i[47];
  assign o[24413] = i[47];
  assign o[24414] = i[47];
  assign o[24415] = i[47];
  assign o[24416] = i[47];
  assign o[24417] = i[47];
  assign o[24418] = i[47];
  assign o[24419] = i[47];
  assign o[24420] = i[47];
  assign o[24421] = i[47];
  assign o[24422] = i[47];
  assign o[24423] = i[47];
  assign o[24424] = i[47];
  assign o[24425] = i[47];
  assign o[24426] = i[47];
  assign o[24427] = i[47];
  assign o[24428] = i[47];
  assign o[24429] = i[47];
  assign o[24430] = i[47];
  assign o[24431] = i[47];
  assign o[24432] = i[47];
  assign o[24433] = i[47];
  assign o[24434] = i[47];
  assign o[24435] = i[47];
  assign o[24436] = i[47];
  assign o[24437] = i[47];
  assign o[24438] = i[47];
  assign o[24439] = i[47];
  assign o[24440] = i[47];
  assign o[24441] = i[47];
  assign o[24442] = i[47];
  assign o[24443] = i[47];
  assign o[24444] = i[47];
  assign o[24445] = i[47];
  assign o[24446] = i[47];
  assign o[24447] = i[47];
  assign o[24448] = i[47];
  assign o[24449] = i[47];
  assign o[24450] = i[47];
  assign o[24451] = i[47];
  assign o[24452] = i[47];
  assign o[24453] = i[47];
  assign o[24454] = i[47];
  assign o[24455] = i[47];
  assign o[24456] = i[47];
  assign o[24457] = i[47];
  assign o[24458] = i[47];
  assign o[24459] = i[47];
  assign o[24460] = i[47];
  assign o[24461] = i[47];
  assign o[24462] = i[47];
  assign o[24463] = i[47];
  assign o[24464] = i[47];
  assign o[24465] = i[47];
  assign o[24466] = i[47];
  assign o[24467] = i[47];
  assign o[24468] = i[47];
  assign o[24469] = i[47];
  assign o[24470] = i[47];
  assign o[24471] = i[47];
  assign o[24472] = i[47];
  assign o[24473] = i[47];
  assign o[24474] = i[47];
  assign o[24475] = i[47];
  assign o[24476] = i[47];
  assign o[24477] = i[47];
  assign o[24478] = i[47];
  assign o[24479] = i[47];
  assign o[24480] = i[47];
  assign o[24481] = i[47];
  assign o[24482] = i[47];
  assign o[24483] = i[47];
  assign o[24484] = i[47];
  assign o[24485] = i[47];
  assign o[24486] = i[47];
  assign o[24487] = i[47];
  assign o[24488] = i[47];
  assign o[24489] = i[47];
  assign o[24490] = i[47];
  assign o[24491] = i[47];
  assign o[24492] = i[47];
  assign o[24493] = i[47];
  assign o[24494] = i[47];
  assign o[24495] = i[47];
  assign o[24496] = i[47];
  assign o[24497] = i[47];
  assign o[24498] = i[47];
  assign o[24499] = i[47];
  assign o[24500] = i[47];
  assign o[24501] = i[47];
  assign o[24502] = i[47];
  assign o[24503] = i[47];
  assign o[24504] = i[47];
  assign o[24505] = i[47];
  assign o[24506] = i[47];
  assign o[24507] = i[47];
  assign o[24508] = i[47];
  assign o[24509] = i[47];
  assign o[24510] = i[47];
  assign o[24511] = i[47];
  assign o[24512] = i[47];
  assign o[24513] = i[47];
  assign o[24514] = i[47];
  assign o[24515] = i[47];
  assign o[24516] = i[47];
  assign o[24517] = i[47];
  assign o[24518] = i[47];
  assign o[24519] = i[47];
  assign o[24520] = i[47];
  assign o[24521] = i[47];
  assign o[24522] = i[47];
  assign o[24523] = i[47];
  assign o[24524] = i[47];
  assign o[24525] = i[47];
  assign o[24526] = i[47];
  assign o[24527] = i[47];
  assign o[24528] = i[47];
  assign o[24529] = i[47];
  assign o[24530] = i[47];
  assign o[24531] = i[47];
  assign o[24532] = i[47];
  assign o[24533] = i[47];
  assign o[24534] = i[47];
  assign o[24535] = i[47];
  assign o[24536] = i[47];
  assign o[24537] = i[47];
  assign o[24538] = i[47];
  assign o[24539] = i[47];
  assign o[24540] = i[47];
  assign o[24541] = i[47];
  assign o[24542] = i[47];
  assign o[24543] = i[47];
  assign o[24544] = i[47];
  assign o[24545] = i[47];
  assign o[24546] = i[47];
  assign o[24547] = i[47];
  assign o[24548] = i[47];
  assign o[24549] = i[47];
  assign o[24550] = i[47];
  assign o[24551] = i[47];
  assign o[24552] = i[47];
  assign o[24553] = i[47];
  assign o[24554] = i[47];
  assign o[24555] = i[47];
  assign o[24556] = i[47];
  assign o[24557] = i[47];
  assign o[24558] = i[47];
  assign o[24559] = i[47];
  assign o[24560] = i[47];
  assign o[24561] = i[47];
  assign o[24562] = i[47];
  assign o[24563] = i[47];
  assign o[24564] = i[47];
  assign o[24565] = i[47];
  assign o[24566] = i[47];
  assign o[24567] = i[47];
  assign o[24568] = i[47];
  assign o[24569] = i[47];
  assign o[24570] = i[47];
  assign o[24571] = i[47];
  assign o[24572] = i[47];
  assign o[24573] = i[47];
  assign o[24574] = i[47];
  assign o[24575] = i[47];
  assign o[23552] = i[46];
  assign o[23553] = i[46];
  assign o[23554] = i[46];
  assign o[23555] = i[46];
  assign o[23556] = i[46];
  assign o[23557] = i[46];
  assign o[23558] = i[46];
  assign o[23559] = i[46];
  assign o[23560] = i[46];
  assign o[23561] = i[46];
  assign o[23562] = i[46];
  assign o[23563] = i[46];
  assign o[23564] = i[46];
  assign o[23565] = i[46];
  assign o[23566] = i[46];
  assign o[23567] = i[46];
  assign o[23568] = i[46];
  assign o[23569] = i[46];
  assign o[23570] = i[46];
  assign o[23571] = i[46];
  assign o[23572] = i[46];
  assign o[23573] = i[46];
  assign o[23574] = i[46];
  assign o[23575] = i[46];
  assign o[23576] = i[46];
  assign o[23577] = i[46];
  assign o[23578] = i[46];
  assign o[23579] = i[46];
  assign o[23580] = i[46];
  assign o[23581] = i[46];
  assign o[23582] = i[46];
  assign o[23583] = i[46];
  assign o[23584] = i[46];
  assign o[23585] = i[46];
  assign o[23586] = i[46];
  assign o[23587] = i[46];
  assign o[23588] = i[46];
  assign o[23589] = i[46];
  assign o[23590] = i[46];
  assign o[23591] = i[46];
  assign o[23592] = i[46];
  assign o[23593] = i[46];
  assign o[23594] = i[46];
  assign o[23595] = i[46];
  assign o[23596] = i[46];
  assign o[23597] = i[46];
  assign o[23598] = i[46];
  assign o[23599] = i[46];
  assign o[23600] = i[46];
  assign o[23601] = i[46];
  assign o[23602] = i[46];
  assign o[23603] = i[46];
  assign o[23604] = i[46];
  assign o[23605] = i[46];
  assign o[23606] = i[46];
  assign o[23607] = i[46];
  assign o[23608] = i[46];
  assign o[23609] = i[46];
  assign o[23610] = i[46];
  assign o[23611] = i[46];
  assign o[23612] = i[46];
  assign o[23613] = i[46];
  assign o[23614] = i[46];
  assign o[23615] = i[46];
  assign o[23616] = i[46];
  assign o[23617] = i[46];
  assign o[23618] = i[46];
  assign o[23619] = i[46];
  assign o[23620] = i[46];
  assign o[23621] = i[46];
  assign o[23622] = i[46];
  assign o[23623] = i[46];
  assign o[23624] = i[46];
  assign o[23625] = i[46];
  assign o[23626] = i[46];
  assign o[23627] = i[46];
  assign o[23628] = i[46];
  assign o[23629] = i[46];
  assign o[23630] = i[46];
  assign o[23631] = i[46];
  assign o[23632] = i[46];
  assign o[23633] = i[46];
  assign o[23634] = i[46];
  assign o[23635] = i[46];
  assign o[23636] = i[46];
  assign o[23637] = i[46];
  assign o[23638] = i[46];
  assign o[23639] = i[46];
  assign o[23640] = i[46];
  assign o[23641] = i[46];
  assign o[23642] = i[46];
  assign o[23643] = i[46];
  assign o[23644] = i[46];
  assign o[23645] = i[46];
  assign o[23646] = i[46];
  assign o[23647] = i[46];
  assign o[23648] = i[46];
  assign o[23649] = i[46];
  assign o[23650] = i[46];
  assign o[23651] = i[46];
  assign o[23652] = i[46];
  assign o[23653] = i[46];
  assign o[23654] = i[46];
  assign o[23655] = i[46];
  assign o[23656] = i[46];
  assign o[23657] = i[46];
  assign o[23658] = i[46];
  assign o[23659] = i[46];
  assign o[23660] = i[46];
  assign o[23661] = i[46];
  assign o[23662] = i[46];
  assign o[23663] = i[46];
  assign o[23664] = i[46];
  assign o[23665] = i[46];
  assign o[23666] = i[46];
  assign o[23667] = i[46];
  assign o[23668] = i[46];
  assign o[23669] = i[46];
  assign o[23670] = i[46];
  assign o[23671] = i[46];
  assign o[23672] = i[46];
  assign o[23673] = i[46];
  assign o[23674] = i[46];
  assign o[23675] = i[46];
  assign o[23676] = i[46];
  assign o[23677] = i[46];
  assign o[23678] = i[46];
  assign o[23679] = i[46];
  assign o[23680] = i[46];
  assign o[23681] = i[46];
  assign o[23682] = i[46];
  assign o[23683] = i[46];
  assign o[23684] = i[46];
  assign o[23685] = i[46];
  assign o[23686] = i[46];
  assign o[23687] = i[46];
  assign o[23688] = i[46];
  assign o[23689] = i[46];
  assign o[23690] = i[46];
  assign o[23691] = i[46];
  assign o[23692] = i[46];
  assign o[23693] = i[46];
  assign o[23694] = i[46];
  assign o[23695] = i[46];
  assign o[23696] = i[46];
  assign o[23697] = i[46];
  assign o[23698] = i[46];
  assign o[23699] = i[46];
  assign o[23700] = i[46];
  assign o[23701] = i[46];
  assign o[23702] = i[46];
  assign o[23703] = i[46];
  assign o[23704] = i[46];
  assign o[23705] = i[46];
  assign o[23706] = i[46];
  assign o[23707] = i[46];
  assign o[23708] = i[46];
  assign o[23709] = i[46];
  assign o[23710] = i[46];
  assign o[23711] = i[46];
  assign o[23712] = i[46];
  assign o[23713] = i[46];
  assign o[23714] = i[46];
  assign o[23715] = i[46];
  assign o[23716] = i[46];
  assign o[23717] = i[46];
  assign o[23718] = i[46];
  assign o[23719] = i[46];
  assign o[23720] = i[46];
  assign o[23721] = i[46];
  assign o[23722] = i[46];
  assign o[23723] = i[46];
  assign o[23724] = i[46];
  assign o[23725] = i[46];
  assign o[23726] = i[46];
  assign o[23727] = i[46];
  assign o[23728] = i[46];
  assign o[23729] = i[46];
  assign o[23730] = i[46];
  assign o[23731] = i[46];
  assign o[23732] = i[46];
  assign o[23733] = i[46];
  assign o[23734] = i[46];
  assign o[23735] = i[46];
  assign o[23736] = i[46];
  assign o[23737] = i[46];
  assign o[23738] = i[46];
  assign o[23739] = i[46];
  assign o[23740] = i[46];
  assign o[23741] = i[46];
  assign o[23742] = i[46];
  assign o[23743] = i[46];
  assign o[23744] = i[46];
  assign o[23745] = i[46];
  assign o[23746] = i[46];
  assign o[23747] = i[46];
  assign o[23748] = i[46];
  assign o[23749] = i[46];
  assign o[23750] = i[46];
  assign o[23751] = i[46];
  assign o[23752] = i[46];
  assign o[23753] = i[46];
  assign o[23754] = i[46];
  assign o[23755] = i[46];
  assign o[23756] = i[46];
  assign o[23757] = i[46];
  assign o[23758] = i[46];
  assign o[23759] = i[46];
  assign o[23760] = i[46];
  assign o[23761] = i[46];
  assign o[23762] = i[46];
  assign o[23763] = i[46];
  assign o[23764] = i[46];
  assign o[23765] = i[46];
  assign o[23766] = i[46];
  assign o[23767] = i[46];
  assign o[23768] = i[46];
  assign o[23769] = i[46];
  assign o[23770] = i[46];
  assign o[23771] = i[46];
  assign o[23772] = i[46];
  assign o[23773] = i[46];
  assign o[23774] = i[46];
  assign o[23775] = i[46];
  assign o[23776] = i[46];
  assign o[23777] = i[46];
  assign o[23778] = i[46];
  assign o[23779] = i[46];
  assign o[23780] = i[46];
  assign o[23781] = i[46];
  assign o[23782] = i[46];
  assign o[23783] = i[46];
  assign o[23784] = i[46];
  assign o[23785] = i[46];
  assign o[23786] = i[46];
  assign o[23787] = i[46];
  assign o[23788] = i[46];
  assign o[23789] = i[46];
  assign o[23790] = i[46];
  assign o[23791] = i[46];
  assign o[23792] = i[46];
  assign o[23793] = i[46];
  assign o[23794] = i[46];
  assign o[23795] = i[46];
  assign o[23796] = i[46];
  assign o[23797] = i[46];
  assign o[23798] = i[46];
  assign o[23799] = i[46];
  assign o[23800] = i[46];
  assign o[23801] = i[46];
  assign o[23802] = i[46];
  assign o[23803] = i[46];
  assign o[23804] = i[46];
  assign o[23805] = i[46];
  assign o[23806] = i[46];
  assign o[23807] = i[46];
  assign o[23808] = i[46];
  assign o[23809] = i[46];
  assign o[23810] = i[46];
  assign o[23811] = i[46];
  assign o[23812] = i[46];
  assign o[23813] = i[46];
  assign o[23814] = i[46];
  assign o[23815] = i[46];
  assign o[23816] = i[46];
  assign o[23817] = i[46];
  assign o[23818] = i[46];
  assign o[23819] = i[46];
  assign o[23820] = i[46];
  assign o[23821] = i[46];
  assign o[23822] = i[46];
  assign o[23823] = i[46];
  assign o[23824] = i[46];
  assign o[23825] = i[46];
  assign o[23826] = i[46];
  assign o[23827] = i[46];
  assign o[23828] = i[46];
  assign o[23829] = i[46];
  assign o[23830] = i[46];
  assign o[23831] = i[46];
  assign o[23832] = i[46];
  assign o[23833] = i[46];
  assign o[23834] = i[46];
  assign o[23835] = i[46];
  assign o[23836] = i[46];
  assign o[23837] = i[46];
  assign o[23838] = i[46];
  assign o[23839] = i[46];
  assign o[23840] = i[46];
  assign o[23841] = i[46];
  assign o[23842] = i[46];
  assign o[23843] = i[46];
  assign o[23844] = i[46];
  assign o[23845] = i[46];
  assign o[23846] = i[46];
  assign o[23847] = i[46];
  assign o[23848] = i[46];
  assign o[23849] = i[46];
  assign o[23850] = i[46];
  assign o[23851] = i[46];
  assign o[23852] = i[46];
  assign o[23853] = i[46];
  assign o[23854] = i[46];
  assign o[23855] = i[46];
  assign o[23856] = i[46];
  assign o[23857] = i[46];
  assign o[23858] = i[46];
  assign o[23859] = i[46];
  assign o[23860] = i[46];
  assign o[23861] = i[46];
  assign o[23862] = i[46];
  assign o[23863] = i[46];
  assign o[23864] = i[46];
  assign o[23865] = i[46];
  assign o[23866] = i[46];
  assign o[23867] = i[46];
  assign o[23868] = i[46];
  assign o[23869] = i[46];
  assign o[23870] = i[46];
  assign o[23871] = i[46];
  assign o[23872] = i[46];
  assign o[23873] = i[46];
  assign o[23874] = i[46];
  assign o[23875] = i[46];
  assign o[23876] = i[46];
  assign o[23877] = i[46];
  assign o[23878] = i[46];
  assign o[23879] = i[46];
  assign o[23880] = i[46];
  assign o[23881] = i[46];
  assign o[23882] = i[46];
  assign o[23883] = i[46];
  assign o[23884] = i[46];
  assign o[23885] = i[46];
  assign o[23886] = i[46];
  assign o[23887] = i[46];
  assign o[23888] = i[46];
  assign o[23889] = i[46];
  assign o[23890] = i[46];
  assign o[23891] = i[46];
  assign o[23892] = i[46];
  assign o[23893] = i[46];
  assign o[23894] = i[46];
  assign o[23895] = i[46];
  assign o[23896] = i[46];
  assign o[23897] = i[46];
  assign o[23898] = i[46];
  assign o[23899] = i[46];
  assign o[23900] = i[46];
  assign o[23901] = i[46];
  assign o[23902] = i[46];
  assign o[23903] = i[46];
  assign o[23904] = i[46];
  assign o[23905] = i[46];
  assign o[23906] = i[46];
  assign o[23907] = i[46];
  assign o[23908] = i[46];
  assign o[23909] = i[46];
  assign o[23910] = i[46];
  assign o[23911] = i[46];
  assign o[23912] = i[46];
  assign o[23913] = i[46];
  assign o[23914] = i[46];
  assign o[23915] = i[46];
  assign o[23916] = i[46];
  assign o[23917] = i[46];
  assign o[23918] = i[46];
  assign o[23919] = i[46];
  assign o[23920] = i[46];
  assign o[23921] = i[46];
  assign o[23922] = i[46];
  assign o[23923] = i[46];
  assign o[23924] = i[46];
  assign o[23925] = i[46];
  assign o[23926] = i[46];
  assign o[23927] = i[46];
  assign o[23928] = i[46];
  assign o[23929] = i[46];
  assign o[23930] = i[46];
  assign o[23931] = i[46];
  assign o[23932] = i[46];
  assign o[23933] = i[46];
  assign o[23934] = i[46];
  assign o[23935] = i[46];
  assign o[23936] = i[46];
  assign o[23937] = i[46];
  assign o[23938] = i[46];
  assign o[23939] = i[46];
  assign o[23940] = i[46];
  assign o[23941] = i[46];
  assign o[23942] = i[46];
  assign o[23943] = i[46];
  assign o[23944] = i[46];
  assign o[23945] = i[46];
  assign o[23946] = i[46];
  assign o[23947] = i[46];
  assign o[23948] = i[46];
  assign o[23949] = i[46];
  assign o[23950] = i[46];
  assign o[23951] = i[46];
  assign o[23952] = i[46];
  assign o[23953] = i[46];
  assign o[23954] = i[46];
  assign o[23955] = i[46];
  assign o[23956] = i[46];
  assign o[23957] = i[46];
  assign o[23958] = i[46];
  assign o[23959] = i[46];
  assign o[23960] = i[46];
  assign o[23961] = i[46];
  assign o[23962] = i[46];
  assign o[23963] = i[46];
  assign o[23964] = i[46];
  assign o[23965] = i[46];
  assign o[23966] = i[46];
  assign o[23967] = i[46];
  assign o[23968] = i[46];
  assign o[23969] = i[46];
  assign o[23970] = i[46];
  assign o[23971] = i[46];
  assign o[23972] = i[46];
  assign o[23973] = i[46];
  assign o[23974] = i[46];
  assign o[23975] = i[46];
  assign o[23976] = i[46];
  assign o[23977] = i[46];
  assign o[23978] = i[46];
  assign o[23979] = i[46];
  assign o[23980] = i[46];
  assign o[23981] = i[46];
  assign o[23982] = i[46];
  assign o[23983] = i[46];
  assign o[23984] = i[46];
  assign o[23985] = i[46];
  assign o[23986] = i[46];
  assign o[23987] = i[46];
  assign o[23988] = i[46];
  assign o[23989] = i[46];
  assign o[23990] = i[46];
  assign o[23991] = i[46];
  assign o[23992] = i[46];
  assign o[23993] = i[46];
  assign o[23994] = i[46];
  assign o[23995] = i[46];
  assign o[23996] = i[46];
  assign o[23997] = i[46];
  assign o[23998] = i[46];
  assign o[23999] = i[46];
  assign o[24000] = i[46];
  assign o[24001] = i[46];
  assign o[24002] = i[46];
  assign o[24003] = i[46];
  assign o[24004] = i[46];
  assign o[24005] = i[46];
  assign o[24006] = i[46];
  assign o[24007] = i[46];
  assign o[24008] = i[46];
  assign o[24009] = i[46];
  assign o[24010] = i[46];
  assign o[24011] = i[46];
  assign o[24012] = i[46];
  assign o[24013] = i[46];
  assign o[24014] = i[46];
  assign o[24015] = i[46];
  assign o[24016] = i[46];
  assign o[24017] = i[46];
  assign o[24018] = i[46];
  assign o[24019] = i[46];
  assign o[24020] = i[46];
  assign o[24021] = i[46];
  assign o[24022] = i[46];
  assign o[24023] = i[46];
  assign o[24024] = i[46];
  assign o[24025] = i[46];
  assign o[24026] = i[46];
  assign o[24027] = i[46];
  assign o[24028] = i[46];
  assign o[24029] = i[46];
  assign o[24030] = i[46];
  assign o[24031] = i[46];
  assign o[24032] = i[46];
  assign o[24033] = i[46];
  assign o[24034] = i[46];
  assign o[24035] = i[46];
  assign o[24036] = i[46];
  assign o[24037] = i[46];
  assign o[24038] = i[46];
  assign o[24039] = i[46];
  assign o[24040] = i[46];
  assign o[24041] = i[46];
  assign o[24042] = i[46];
  assign o[24043] = i[46];
  assign o[24044] = i[46];
  assign o[24045] = i[46];
  assign o[24046] = i[46];
  assign o[24047] = i[46];
  assign o[24048] = i[46];
  assign o[24049] = i[46];
  assign o[24050] = i[46];
  assign o[24051] = i[46];
  assign o[24052] = i[46];
  assign o[24053] = i[46];
  assign o[24054] = i[46];
  assign o[24055] = i[46];
  assign o[24056] = i[46];
  assign o[24057] = i[46];
  assign o[24058] = i[46];
  assign o[24059] = i[46];
  assign o[24060] = i[46];
  assign o[24061] = i[46];
  assign o[24062] = i[46];
  assign o[24063] = i[46];
  assign o[23040] = i[45];
  assign o[23041] = i[45];
  assign o[23042] = i[45];
  assign o[23043] = i[45];
  assign o[23044] = i[45];
  assign o[23045] = i[45];
  assign o[23046] = i[45];
  assign o[23047] = i[45];
  assign o[23048] = i[45];
  assign o[23049] = i[45];
  assign o[23050] = i[45];
  assign o[23051] = i[45];
  assign o[23052] = i[45];
  assign o[23053] = i[45];
  assign o[23054] = i[45];
  assign o[23055] = i[45];
  assign o[23056] = i[45];
  assign o[23057] = i[45];
  assign o[23058] = i[45];
  assign o[23059] = i[45];
  assign o[23060] = i[45];
  assign o[23061] = i[45];
  assign o[23062] = i[45];
  assign o[23063] = i[45];
  assign o[23064] = i[45];
  assign o[23065] = i[45];
  assign o[23066] = i[45];
  assign o[23067] = i[45];
  assign o[23068] = i[45];
  assign o[23069] = i[45];
  assign o[23070] = i[45];
  assign o[23071] = i[45];
  assign o[23072] = i[45];
  assign o[23073] = i[45];
  assign o[23074] = i[45];
  assign o[23075] = i[45];
  assign o[23076] = i[45];
  assign o[23077] = i[45];
  assign o[23078] = i[45];
  assign o[23079] = i[45];
  assign o[23080] = i[45];
  assign o[23081] = i[45];
  assign o[23082] = i[45];
  assign o[23083] = i[45];
  assign o[23084] = i[45];
  assign o[23085] = i[45];
  assign o[23086] = i[45];
  assign o[23087] = i[45];
  assign o[23088] = i[45];
  assign o[23089] = i[45];
  assign o[23090] = i[45];
  assign o[23091] = i[45];
  assign o[23092] = i[45];
  assign o[23093] = i[45];
  assign o[23094] = i[45];
  assign o[23095] = i[45];
  assign o[23096] = i[45];
  assign o[23097] = i[45];
  assign o[23098] = i[45];
  assign o[23099] = i[45];
  assign o[23100] = i[45];
  assign o[23101] = i[45];
  assign o[23102] = i[45];
  assign o[23103] = i[45];
  assign o[23104] = i[45];
  assign o[23105] = i[45];
  assign o[23106] = i[45];
  assign o[23107] = i[45];
  assign o[23108] = i[45];
  assign o[23109] = i[45];
  assign o[23110] = i[45];
  assign o[23111] = i[45];
  assign o[23112] = i[45];
  assign o[23113] = i[45];
  assign o[23114] = i[45];
  assign o[23115] = i[45];
  assign o[23116] = i[45];
  assign o[23117] = i[45];
  assign o[23118] = i[45];
  assign o[23119] = i[45];
  assign o[23120] = i[45];
  assign o[23121] = i[45];
  assign o[23122] = i[45];
  assign o[23123] = i[45];
  assign o[23124] = i[45];
  assign o[23125] = i[45];
  assign o[23126] = i[45];
  assign o[23127] = i[45];
  assign o[23128] = i[45];
  assign o[23129] = i[45];
  assign o[23130] = i[45];
  assign o[23131] = i[45];
  assign o[23132] = i[45];
  assign o[23133] = i[45];
  assign o[23134] = i[45];
  assign o[23135] = i[45];
  assign o[23136] = i[45];
  assign o[23137] = i[45];
  assign o[23138] = i[45];
  assign o[23139] = i[45];
  assign o[23140] = i[45];
  assign o[23141] = i[45];
  assign o[23142] = i[45];
  assign o[23143] = i[45];
  assign o[23144] = i[45];
  assign o[23145] = i[45];
  assign o[23146] = i[45];
  assign o[23147] = i[45];
  assign o[23148] = i[45];
  assign o[23149] = i[45];
  assign o[23150] = i[45];
  assign o[23151] = i[45];
  assign o[23152] = i[45];
  assign o[23153] = i[45];
  assign o[23154] = i[45];
  assign o[23155] = i[45];
  assign o[23156] = i[45];
  assign o[23157] = i[45];
  assign o[23158] = i[45];
  assign o[23159] = i[45];
  assign o[23160] = i[45];
  assign o[23161] = i[45];
  assign o[23162] = i[45];
  assign o[23163] = i[45];
  assign o[23164] = i[45];
  assign o[23165] = i[45];
  assign o[23166] = i[45];
  assign o[23167] = i[45];
  assign o[23168] = i[45];
  assign o[23169] = i[45];
  assign o[23170] = i[45];
  assign o[23171] = i[45];
  assign o[23172] = i[45];
  assign o[23173] = i[45];
  assign o[23174] = i[45];
  assign o[23175] = i[45];
  assign o[23176] = i[45];
  assign o[23177] = i[45];
  assign o[23178] = i[45];
  assign o[23179] = i[45];
  assign o[23180] = i[45];
  assign o[23181] = i[45];
  assign o[23182] = i[45];
  assign o[23183] = i[45];
  assign o[23184] = i[45];
  assign o[23185] = i[45];
  assign o[23186] = i[45];
  assign o[23187] = i[45];
  assign o[23188] = i[45];
  assign o[23189] = i[45];
  assign o[23190] = i[45];
  assign o[23191] = i[45];
  assign o[23192] = i[45];
  assign o[23193] = i[45];
  assign o[23194] = i[45];
  assign o[23195] = i[45];
  assign o[23196] = i[45];
  assign o[23197] = i[45];
  assign o[23198] = i[45];
  assign o[23199] = i[45];
  assign o[23200] = i[45];
  assign o[23201] = i[45];
  assign o[23202] = i[45];
  assign o[23203] = i[45];
  assign o[23204] = i[45];
  assign o[23205] = i[45];
  assign o[23206] = i[45];
  assign o[23207] = i[45];
  assign o[23208] = i[45];
  assign o[23209] = i[45];
  assign o[23210] = i[45];
  assign o[23211] = i[45];
  assign o[23212] = i[45];
  assign o[23213] = i[45];
  assign o[23214] = i[45];
  assign o[23215] = i[45];
  assign o[23216] = i[45];
  assign o[23217] = i[45];
  assign o[23218] = i[45];
  assign o[23219] = i[45];
  assign o[23220] = i[45];
  assign o[23221] = i[45];
  assign o[23222] = i[45];
  assign o[23223] = i[45];
  assign o[23224] = i[45];
  assign o[23225] = i[45];
  assign o[23226] = i[45];
  assign o[23227] = i[45];
  assign o[23228] = i[45];
  assign o[23229] = i[45];
  assign o[23230] = i[45];
  assign o[23231] = i[45];
  assign o[23232] = i[45];
  assign o[23233] = i[45];
  assign o[23234] = i[45];
  assign o[23235] = i[45];
  assign o[23236] = i[45];
  assign o[23237] = i[45];
  assign o[23238] = i[45];
  assign o[23239] = i[45];
  assign o[23240] = i[45];
  assign o[23241] = i[45];
  assign o[23242] = i[45];
  assign o[23243] = i[45];
  assign o[23244] = i[45];
  assign o[23245] = i[45];
  assign o[23246] = i[45];
  assign o[23247] = i[45];
  assign o[23248] = i[45];
  assign o[23249] = i[45];
  assign o[23250] = i[45];
  assign o[23251] = i[45];
  assign o[23252] = i[45];
  assign o[23253] = i[45];
  assign o[23254] = i[45];
  assign o[23255] = i[45];
  assign o[23256] = i[45];
  assign o[23257] = i[45];
  assign o[23258] = i[45];
  assign o[23259] = i[45];
  assign o[23260] = i[45];
  assign o[23261] = i[45];
  assign o[23262] = i[45];
  assign o[23263] = i[45];
  assign o[23264] = i[45];
  assign o[23265] = i[45];
  assign o[23266] = i[45];
  assign o[23267] = i[45];
  assign o[23268] = i[45];
  assign o[23269] = i[45];
  assign o[23270] = i[45];
  assign o[23271] = i[45];
  assign o[23272] = i[45];
  assign o[23273] = i[45];
  assign o[23274] = i[45];
  assign o[23275] = i[45];
  assign o[23276] = i[45];
  assign o[23277] = i[45];
  assign o[23278] = i[45];
  assign o[23279] = i[45];
  assign o[23280] = i[45];
  assign o[23281] = i[45];
  assign o[23282] = i[45];
  assign o[23283] = i[45];
  assign o[23284] = i[45];
  assign o[23285] = i[45];
  assign o[23286] = i[45];
  assign o[23287] = i[45];
  assign o[23288] = i[45];
  assign o[23289] = i[45];
  assign o[23290] = i[45];
  assign o[23291] = i[45];
  assign o[23292] = i[45];
  assign o[23293] = i[45];
  assign o[23294] = i[45];
  assign o[23295] = i[45];
  assign o[23296] = i[45];
  assign o[23297] = i[45];
  assign o[23298] = i[45];
  assign o[23299] = i[45];
  assign o[23300] = i[45];
  assign o[23301] = i[45];
  assign o[23302] = i[45];
  assign o[23303] = i[45];
  assign o[23304] = i[45];
  assign o[23305] = i[45];
  assign o[23306] = i[45];
  assign o[23307] = i[45];
  assign o[23308] = i[45];
  assign o[23309] = i[45];
  assign o[23310] = i[45];
  assign o[23311] = i[45];
  assign o[23312] = i[45];
  assign o[23313] = i[45];
  assign o[23314] = i[45];
  assign o[23315] = i[45];
  assign o[23316] = i[45];
  assign o[23317] = i[45];
  assign o[23318] = i[45];
  assign o[23319] = i[45];
  assign o[23320] = i[45];
  assign o[23321] = i[45];
  assign o[23322] = i[45];
  assign o[23323] = i[45];
  assign o[23324] = i[45];
  assign o[23325] = i[45];
  assign o[23326] = i[45];
  assign o[23327] = i[45];
  assign o[23328] = i[45];
  assign o[23329] = i[45];
  assign o[23330] = i[45];
  assign o[23331] = i[45];
  assign o[23332] = i[45];
  assign o[23333] = i[45];
  assign o[23334] = i[45];
  assign o[23335] = i[45];
  assign o[23336] = i[45];
  assign o[23337] = i[45];
  assign o[23338] = i[45];
  assign o[23339] = i[45];
  assign o[23340] = i[45];
  assign o[23341] = i[45];
  assign o[23342] = i[45];
  assign o[23343] = i[45];
  assign o[23344] = i[45];
  assign o[23345] = i[45];
  assign o[23346] = i[45];
  assign o[23347] = i[45];
  assign o[23348] = i[45];
  assign o[23349] = i[45];
  assign o[23350] = i[45];
  assign o[23351] = i[45];
  assign o[23352] = i[45];
  assign o[23353] = i[45];
  assign o[23354] = i[45];
  assign o[23355] = i[45];
  assign o[23356] = i[45];
  assign o[23357] = i[45];
  assign o[23358] = i[45];
  assign o[23359] = i[45];
  assign o[23360] = i[45];
  assign o[23361] = i[45];
  assign o[23362] = i[45];
  assign o[23363] = i[45];
  assign o[23364] = i[45];
  assign o[23365] = i[45];
  assign o[23366] = i[45];
  assign o[23367] = i[45];
  assign o[23368] = i[45];
  assign o[23369] = i[45];
  assign o[23370] = i[45];
  assign o[23371] = i[45];
  assign o[23372] = i[45];
  assign o[23373] = i[45];
  assign o[23374] = i[45];
  assign o[23375] = i[45];
  assign o[23376] = i[45];
  assign o[23377] = i[45];
  assign o[23378] = i[45];
  assign o[23379] = i[45];
  assign o[23380] = i[45];
  assign o[23381] = i[45];
  assign o[23382] = i[45];
  assign o[23383] = i[45];
  assign o[23384] = i[45];
  assign o[23385] = i[45];
  assign o[23386] = i[45];
  assign o[23387] = i[45];
  assign o[23388] = i[45];
  assign o[23389] = i[45];
  assign o[23390] = i[45];
  assign o[23391] = i[45];
  assign o[23392] = i[45];
  assign o[23393] = i[45];
  assign o[23394] = i[45];
  assign o[23395] = i[45];
  assign o[23396] = i[45];
  assign o[23397] = i[45];
  assign o[23398] = i[45];
  assign o[23399] = i[45];
  assign o[23400] = i[45];
  assign o[23401] = i[45];
  assign o[23402] = i[45];
  assign o[23403] = i[45];
  assign o[23404] = i[45];
  assign o[23405] = i[45];
  assign o[23406] = i[45];
  assign o[23407] = i[45];
  assign o[23408] = i[45];
  assign o[23409] = i[45];
  assign o[23410] = i[45];
  assign o[23411] = i[45];
  assign o[23412] = i[45];
  assign o[23413] = i[45];
  assign o[23414] = i[45];
  assign o[23415] = i[45];
  assign o[23416] = i[45];
  assign o[23417] = i[45];
  assign o[23418] = i[45];
  assign o[23419] = i[45];
  assign o[23420] = i[45];
  assign o[23421] = i[45];
  assign o[23422] = i[45];
  assign o[23423] = i[45];
  assign o[23424] = i[45];
  assign o[23425] = i[45];
  assign o[23426] = i[45];
  assign o[23427] = i[45];
  assign o[23428] = i[45];
  assign o[23429] = i[45];
  assign o[23430] = i[45];
  assign o[23431] = i[45];
  assign o[23432] = i[45];
  assign o[23433] = i[45];
  assign o[23434] = i[45];
  assign o[23435] = i[45];
  assign o[23436] = i[45];
  assign o[23437] = i[45];
  assign o[23438] = i[45];
  assign o[23439] = i[45];
  assign o[23440] = i[45];
  assign o[23441] = i[45];
  assign o[23442] = i[45];
  assign o[23443] = i[45];
  assign o[23444] = i[45];
  assign o[23445] = i[45];
  assign o[23446] = i[45];
  assign o[23447] = i[45];
  assign o[23448] = i[45];
  assign o[23449] = i[45];
  assign o[23450] = i[45];
  assign o[23451] = i[45];
  assign o[23452] = i[45];
  assign o[23453] = i[45];
  assign o[23454] = i[45];
  assign o[23455] = i[45];
  assign o[23456] = i[45];
  assign o[23457] = i[45];
  assign o[23458] = i[45];
  assign o[23459] = i[45];
  assign o[23460] = i[45];
  assign o[23461] = i[45];
  assign o[23462] = i[45];
  assign o[23463] = i[45];
  assign o[23464] = i[45];
  assign o[23465] = i[45];
  assign o[23466] = i[45];
  assign o[23467] = i[45];
  assign o[23468] = i[45];
  assign o[23469] = i[45];
  assign o[23470] = i[45];
  assign o[23471] = i[45];
  assign o[23472] = i[45];
  assign o[23473] = i[45];
  assign o[23474] = i[45];
  assign o[23475] = i[45];
  assign o[23476] = i[45];
  assign o[23477] = i[45];
  assign o[23478] = i[45];
  assign o[23479] = i[45];
  assign o[23480] = i[45];
  assign o[23481] = i[45];
  assign o[23482] = i[45];
  assign o[23483] = i[45];
  assign o[23484] = i[45];
  assign o[23485] = i[45];
  assign o[23486] = i[45];
  assign o[23487] = i[45];
  assign o[23488] = i[45];
  assign o[23489] = i[45];
  assign o[23490] = i[45];
  assign o[23491] = i[45];
  assign o[23492] = i[45];
  assign o[23493] = i[45];
  assign o[23494] = i[45];
  assign o[23495] = i[45];
  assign o[23496] = i[45];
  assign o[23497] = i[45];
  assign o[23498] = i[45];
  assign o[23499] = i[45];
  assign o[23500] = i[45];
  assign o[23501] = i[45];
  assign o[23502] = i[45];
  assign o[23503] = i[45];
  assign o[23504] = i[45];
  assign o[23505] = i[45];
  assign o[23506] = i[45];
  assign o[23507] = i[45];
  assign o[23508] = i[45];
  assign o[23509] = i[45];
  assign o[23510] = i[45];
  assign o[23511] = i[45];
  assign o[23512] = i[45];
  assign o[23513] = i[45];
  assign o[23514] = i[45];
  assign o[23515] = i[45];
  assign o[23516] = i[45];
  assign o[23517] = i[45];
  assign o[23518] = i[45];
  assign o[23519] = i[45];
  assign o[23520] = i[45];
  assign o[23521] = i[45];
  assign o[23522] = i[45];
  assign o[23523] = i[45];
  assign o[23524] = i[45];
  assign o[23525] = i[45];
  assign o[23526] = i[45];
  assign o[23527] = i[45];
  assign o[23528] = i[45];
  assign o[23529] = i[45];
  assign o[23530] = i[45];
  assign o[23531] = i[45];
  assign o[23532] = i[45];
  assign o[23533] = i[45];
  assign o[23534] = i[45];
  assign o[23535] = i[45];
  assign o[23536] = i[45];
  assign o[23537] = i[45];
  assign o[23538] = i[45];
  assign o[23539] = i[45];
  assign o[23540] = i[45];
  assign o[23541] = i[45];
  assign o[23542] = i[45];
  assign o[23543] = i[45];
  assign o[23544] = i[45];
  assign o[23545] = i[45];
  assign o[23546] = i[45];
  assign o[23547] = i[45];
  assign o[23548] = i[45];
  assign o[23549] = i[45];
  assign o[23550] = i[45];
  assign o[23551] = i[45];
  assign o[22528] = i[44];
  assign o[22529] = i[44];
  assign o[22530] = i[44];
  assign o[22531] = i[44];
  assign o[22532] = i[44];
  assign o[22533] = i[44];
  assign o[22534] = i[44];
  assign o[22535] = i[44];
  assign o[22536] = i[44];
  assign o[22537] = i[44];
  assign o[22538] = i[44];
  assign o[22539] = i[44];
  assign o[22540] = i[44];
  assign o[22541] = i[44];
  assign o[22542] = i[44];
  assign o[22543] = i[44];
  assign o[22544] = i[44];
  assign o[22545] = i[44];
  assign o[22546] = i[44];
  assign o[22547] = i[44];
  assign o[22548] = i[44];
  assign o[22549] = i[44];
  assign o[22550] = i[44];
  assign o[22551] = i[44];
  assign o[22552] = i[44];
  assign o[22553] = i[44];
  assign o[22554] = i[44];
  assign o[22555] = i[44];
  assign o[22556] = i[44];
  assign o[22557] = i[44];
  assign o[22558] = i[44];
  assign o[22559] = i[44];
  assign o[22560] = i[44];
  assign o[22561] = i[44];
  assign o[22562] = i[44];
  assign o[22563] = i[44];
  assign o[22564] = i[44];
  assign o[22565] = i[44];
  assign o[22566] = i[44];
  assign o[22567] = i[44];
  assign o[22568] = i[44];
  assign o[22569] = i[44];
  assign o[22570] = i[44];
  assign o[22571] = i[44];
  assign o[22572] = i[44];
  assign o[22573] = i[44];
  assign o[22574] = i[44];
  assign o[22575] = i[44];
  assign o[22576] = i[44];
  assign o[22577] = i[44];
  assign o[22578] = i[44];
  assign o[22579] = i[44];
  assign o[22580] = i[44];
  assign o[22581] = i[44];
  assign o[22582] = i[44];
  assign o[22583] = i[44];
  assign o[22584] = i[44];
  assign o[22585] = i[44];
  assign o[22586] = i[44];
  assign o[22587] = i[44];
  assign o[22588] = i[44];
  assign o[22589] = i[44];
  assign o[22590] = i[44];
  assign o[22591] = i[44];
  assign o[22592] = i[44];
  assign o[22593] = i[44];
  assign o[22594] = i[44];
  assign o[22595] = i[44];
  assign o[22596] = i[44];
  assign o[22597] = i[44];
  assign o[22598] = i[44];
  assign o[22599] = i[44];
  assign o[22600] = i[44];
  assign o[22601] = i[44];
  assign o[22602] = i[44];
  assign o[22603] = i[44];
  assign o[22604] = i[44];
  assign o[22605] = i[44];
  assign o[22606] = i[44];
  assign o[22607] = i[44];
  assign o[22608] = i[44];
  assign o[22609] = i[44];
  assign o[22610] = i[44];
  assign o[22611] = i[44];
  assign o[22612] = i[44];
  assign o[22613] = i[44];
  assign o[22614] = i[44];
  assign o[22615] = i[44];
  assign o[22616] = i[44];
  assign o[22617] = i[44];
  assign o[22618] = i[44];
  assign o[22619] = i[44];
  assign o[22620] = i[44];
  assign o[22621] = i[44];
  assign o[22622] = i[44];
  assign o[22623] = i[44];
  assign o[22624] = i[44];
  assign o[22625] = i[44];
  assign o[22626] = i[44];
  assign o[22627] = i[44];
  assign o[22628] = i[44];
  assign o[22629] = i[44];
  assign o[22630] = i[44];
  assign o[22631] = i[44];
  assign o[22632] = i[44];
  assign o[22633] = i[44];
  assign o[22634] = i[44];
  assign o[22635] = i[44];
  assign o[22636] = i[44];
  assign o[22637] = i[44];
  assign o[22638] = i[44];
  assign o[22639] = i[44];
  assign o[22640] = i[44];
  assign o[22641] = i[44];
  assign o[22642] = i[44];
  assign o[22643] = i[44];
  assign o[22644] = i[44];
  assign o[22645] = i[44];
  assign o[22646] = i[44];
  assign o[22647] = i[44];
  assign o[22648] = i[44];
  assign o[22649] = i[44];
  assign o[22650] = i[44];
  assign o[22651] = i[44];
  assign o[22652] = i[44];
  assign o[22653] = i[44];
  assign o[22654] = i[44];
  assign o[22655] = i[44];
  assign o[22656] = i[44];
  assign o[22657] = i[44];
  assign o[22658] = i[44];
  assign o[22659] = i[44];
  assign o[22660] = i[44];
  assign o[22661] = i[44];
  assign o[22662] = i[44];
  assign o[22663] = i[44];
  assign o[22664] = i[44];
  assign o[22665] = i[44];
  assign o[22666] = i[44];
  assign o[22667] = i[44];
  assign o[22668] = i[44];
  assign o[22669] = i[44];
  assign o[22670] = i[44];
  assign o[22671] = i[44];
  assign o[22672] = i[44];
  assign o[22673] = i[44];
  assign o[22674] = i[44];
  assign o[22675] = i[44];
  assign o[22676] = i[44];
  assign o[22677] = i[44];
  assign o[22678] = i[44];
  assign o[22679] = i[44];
  assign o[22680] = i[44];
  assign o[22681] = i[44];
  assign o[22682] = i[44];
  assign o[22683] = i[44];
  assign o[22684] = i[44];
  assign o[22685] = i[44];
  assign o[22686] = i[44];
  assign o[22687] = i[44];
  assign o[22688] = i[44];
  assign o[22689] = i[44];
  assign o[22690] = i[44];
  assign o[22691] = i[44];
  assign o[22692] = i[44];
  assign o[22693] = i[44];
  assign o[22694] = i[44];
  assign o[22695] = i[44];
  assign o[22696] = i[44];
  assign o[22697] = i[44];
  assign o[22698] = i[44];
  assign o[22699] = i[44];
  assign o[22700] = i[44];
  assign o[22701] = i[44];
  assign o[22702] = i[44];
  assign o[22703] = i[44];
  assign o[22704] = i[44];
  assign o[22705] = i[44];
  assign o[22706] = i[44];
  assign o[22707] = i[44];
  assign o[22708] = i[44];
  assign o[22709] = i[44];
  assign o[22710] = i[44];
  assign o[22711] = i[44];
  assign o[22712] = i[44];
  assign o[22713] = i[44];
  assign o[22714] = i[44];
  assign o[22715] = i[44];
  assign o[22716] = i[44];
  assign o[22717] = i[44];
  assign o[22718] = i[44];
  assign o[22719] = i[44];
  assign o[22720] = i[44];
  assign o[22721] = i[44];
  assign o[22722] = i[44];
  assign o[22723] = i[44];
  assign o[22724] = i[44];
  assign o[22725] = i[44];
  assign o[22726] = i[44];
  assign o[22727] = i[44];
  assign o[22728] = i[44];
  assign o[22729] = i[44];
  assign o[22730] = i[44];
  assign o[22731] = i[44];
  assign o[22732] = i[44];
  assign o[22733] = i[44];
  assign o[22734] = i[44];
  assign o[22735] = i[44];
  assign o[22736] = i[44];
  assign o[22737] = i[44];
  assign o[22738] = i[44];
  assign o[22739] = i[44];
  assign o[22740] = i[44];
  assign o[22741] = i[44];
  assign o[22742] = i[44];
  assign o[22743] = i[44];
  assign o[22744] = i[44];
  assign o[22745] = i[44];
  assign o[22746] = i[44];
  assign o[22747] = i[44];
  assign o[22748] = i[44];
  assign o[22749] = i[44];
  assign o[22750] = i[44];
  assign o[22751] = i[44];
  assign o[22752] = i[44];
  assign o[22753] = i[44];
  assign o[22754] = i[44];
  assign o[22755] = i[44];
  assign o[22756] = i[44];
  assign o[22757] = i[44];
  assign o[22758] = i[44];
  assign o[22759] = i[44];
  assign o[22760] = i[44];
  assign o[22761] = i[44];
  assign o[22762] = i[44];
  assign o[22763] = i[44];
  assign o[22764] = i[44];
  assign o[22765] = i[44];
  assign o[22766] = i[44];
  assign o[22767] = i[44];
  assign o[22768] = i[44];
  assign o[22769] = i[44];
  assign o[22770] = i[44];
  assign o[22771] = i[44];
  assign o[22772] = i[44];
  assign o[22773] = i[44];
  assign o[22774] = i[44];
  assign o[22775] = i[44];
  assign o[22776] = i[44];
  assign o[22777] = i[44];
  assign o[22778] = i[44];
  assign o[22779] = i[44];
  assign o[22780] = i[44];
  assign o[22781] = i[44];
  assign o[22782] = i[44];
  assign o[22783] = i[44];
  assign o[22784] = i[44];
  assign o[22785] = i[44];
  assign o[22786] = i[44];
  assign o[22787] = i[44];
  assign o[22788] = i[44];
  assign o[22789] = i[44];
  assign o[22790] = i[44];
  assign o[22791] = i[44];
  assign o[22792] = i[44];
  assign o[22793] = i[44];
  assign o[22794] = i[44];
  assign o[22795] = i[44];
  assign o[22796] = i[44];
  assign o[22797] = i[44];
  assign o[22798] = i[44];
  assign o[22799] = i[44];
  assign o[22800] = i[44];
  assign o[22801] = i[44];
  assign o[22802] = i[44];
  assign o[22803] = i[44];
  assign o[22804] = i[44];
  assign o[22805] = i[44];
  assign o[22806] = i[44];
  assign o[22807] = i[44];
  assign o[22808] = i[44];
  assign o[22809] = i[44];
  assign o[22810] = i[44];
  assign o[22811] = i[44];
  assign o[22812] = i[44];
  assign o[22813] = i[44];
  assign o[22814] = i[44];
  assign o[22815] = i[44];
  assign o[22816] = i[44];
  assign o[22817] = i[44];
  assign o[22818] = i[44];
  assign o[22819] = i[44];
  assign o[22820] = i[44];
  assign o[22821] = i[44];
  assign o[22822] = i[44];
  assign o[22823] = i[44];
  assign o[22824] = i[44];
  assign o[22825] = i[44];
  assign o[22826] = i[44];
  assign o[22827] = i[44];
  assign o[22828] = i[44];
  assign o[22829] = i[44];
  assign o[22830] = i[44];
  assign o[22831] = i[44];
  assign o[22832] = i[44];
  assign o[22833] = i[44];
  assign o[22834] = i[44];
  assign o[22835] = i[44];
  assign o[22836] = i[44];
  assign o[22837] = i[44];
  assign o[22838] = i[44];
  assign o[22839] = i[44];
  assign o[22840] = i[44];
  assign o[22841] = i[44];
  assign o[22842] = i[44];
  assign o[22843] = i[44];
  assign o[22844] = i[44];
  assign o[22845] = i[44];
  assign o[22846] = i[44];
  assign o[22847] = i[44];
  assign o[22848] = i[44];
  assign o[22849] = i[44];
  assign o[22850] = i[44];
  assign o[22851] = i[44];
  assign o[22852] = i[44];
  assign o[22853] = i[44];
  assign o[22854] = i[44];
  assign o[22855] = i[44];
  assign o[22856] = i[44];
  assign o[22857] = i[44];
  assign o[22858] = i[44];
  assign o[22859] = i[44];
  assign o[22860] = i[44];
  assign o[22861] = i[44];
  assign o[22862] = i[44];
  assign o[22863] = i[44];
  assign o[22864] = i[44];
  assign o[22865] = i[44];
  assign o[22866] = i[44];
  assign o[22867] = i[44];
  assign o[22868] = i[44];
  assign o[22869] = i[44];
  assign o[22870] = i[44];
  assign o[22871] = i[44];
  assign o[22872] = i[44];
  assign o[22873] = i[44];
  assign o[22874] = i[44];
  assign o[22875] = i[44];
  assign o[22876] = i[44];
  assign o[22877] = i[44];
  assign o[22878] = i[44];
  assign o[22879] = i[44];
  assign o[22880] = i[44];
  assign o[22881] = i[44];
  assign o[22882] = i[44];
  assign o[22883] = i[44];
  assign o[22884] = i[44];
  assign o[22885] = i[44];
  assign o[22886] = i[44];
  assign o[22887] = i[44];
  assign o[22888] = i[44];
  assign o[22889] = i[44];
  assign o[22890] = i[44];
  assign o[22891] = i[44];
  assign o[22892] = i[44];
  assign o[22893] = i[44];
  assign o[22894] = i[44];
  assign o[22895] = i[44];
  assign o[22896] = i[44];
  assign o[22897] = i[44];
  assign o[22898] = i[44];
  assign o[22899] = i[44];
  assign o[22900] = i[44];
  assign o[22901] = i[44];
  assign o[22902] = i[44];
  assign o[22903] = i[44];
  assign o[22904] = i[44];
  assign o[22905] = i[44];
  assign o[22906] = i[44];
  assign o[22907] = i[44];
  assign o[22908] = i[44];
  assign o[22909] = i[44];
  assign o[22910] = i[44];
  assign o[22911] = i[44];
  assign o[22912] = i[44];
  assign o[22913] = i[44];
  assign o[22914] = i[44];
  assign o[22915] = i[44];
  assign o[22916] = i[44];
  assign o[22917] = i[44];
  assign o[22918] = i[44];
  assign o[22919] = i[44];
  assign o[22920] = i[44];
  assign o[22921] = i[44];
  assign o[22922] = i[44];
  assign o[22923] = i[44];
  assign o[22924] = i[44];
  assign o[22925] = i[44];
  assign o[22926] = i[44];
  assign o[22927] = i[44];
  assign o[22928] = i[44];
  assign o[22929] = i[44];
  assign o[22930] = i[44];
  assign o[22931] = i[44];
  assign o[22932] = i[44];
  assign o[22933] = i[44];
  assign o[22934] = i[44];
  assign o[22935] = i[44];
  assign o[22936] = i[44];
  assign o[22937] = i[44];
  assign o[22938] = i[44];
  assign o[22939] = i[44];
  assign o[22940] = i[44];
  assign o[22941] = i[44];
  assign o[22942] = i[44];
  assign o[22943] = i[44];
  assign o[22944] = i[44];
  assign o[22945] = i[44];
  assign o[22946] = i[44];
  assign o[22947] = i[44];
  assign o[22948] = i[44];
  assign o[22949] = i[44];
  assign o[22950] = i[44];
  assign o[22951] = i[44];
  assign o[22952] = i[44];
  assign o[22953] = i[44];
  assign o[22954] = i[44];
  assign o[22955] = i[44];
  assign o[22956] = i[44];
  assign o[22957] = i[44];
  assign o[22958] = i[44];
  assign o[22959] = i[44];
  assign o[22960] = i[44];
  assign o[22961] = i[44];
  assign o[22962] = i[44];
  assign o[22963] = i[44];
  assign o[22964] = i[44];
  assign o[22965] = i[44];
  assign o[22966] = i[44];
  assign o[22967] = i[44];
  assign o[22968] = i[44];
  assign o[22969] = i[44];
  assign o[22970] = i[44];
  assign o[22971] = i[44];
  assign o[22972] = i[44];
  assign o[22973] = i[44];
  assign o[22974] = i[44];
  assign o[22975] = i[44];
  assign o[22976] = i[44];
  assign o[22977] = i[44];
  assign o[22978] = i[44];
  assign o[22979] = i[44];
  assign o[22980] = i[44];
  assign o[22981] = i[44];
  assign o[22982] = i[44];
  assign o[22983] = i[44];
  assign o[22984] = i[44];
  assign o[22985] = i[44];
  assign o[22986] = i[44];
  assign o[22987] = i[44];
  assign o[22988] = i[44];
  assign o[22989] = i[44];
  assign o[22990] = i[44];
  assign o[22991] = i[44];
  assign o[22992] = i[44];
  assign o[22993] = i[44];
  assign o[22994] = i[44];
  assign o[22995] = i[44];
  assign o[22996] = i[44];
  assign o[22997] = i[44];
  assign o[22998] = i[44];
  assign o[22999] = i[44];
  assign o[23000] = i[44];
  assign o[23001] = i[44];
  assign o[23002] = i[44];
  assign o[23003] = i[44];
  assign o[23004] = i[44];
  assign o[23005] = i[44];
  assign o[23006] = i[44];
  assign o[23007] = i[44];
  assign o[23008] = i[44];
  assign o[23009] = i[44];
  assign o[23010] = i[44];
  assign o[23011] = i[44];
  assign o[23012] = i[44];
  assign o[23013] = i[44];
  assign o[23014] = i[44];
  assign o[23015] = i[44];
  assign o[23016] = i[44];
  assign o[23017] = i[44];
  assign o[23018] = i[44];
  assign o[23019] = i[44];
  assign o[23020] = i[44];
  assign o[23021] = i[44];
  assign o[23022] = i[44];
  assign o[23023] = i[44];
  assign o[23024] = i[44];
  assign o[23025] = i[44];
  assign o[23026] = i[44];
  assign o[23027] = i[44];
  assign o[23028] = i[44];
  assign o[23029] = i[44];
  assign o[23030] = i[44];
  assign o[23031] = i[44];
  assign o[23032] = i[44];
  assign o[23033] = i[44];
  assign o[23034] = i[44];
  assign o[23035] = i[44];
  assign o[23036] = i[44];
  assign o[23037] = i[44];
  assign o[23038] = i[44];
  assign o[23039] = i[44];
  assign o[22016] = i[43];
  assign o[22017] = i[43];
  assign o[22018] = i[43];
  assign o[22019] = i[43];
  assign o[22020] = i[43];
  assign o[22021] = i[43];
  assign o[22022] = i[43];
  assign o[22023] = i[43];
  assign o[22024] = i[43];
  assign o[22025] = i[43];
  assign o[22026] = i[43];
  assign o[22027] = i[43];
  assign o[22028] = i[43];
  assign o[22029] = i[43];
  assign o[22030] = i[43];
  assign o[22031] = i[43];
  assign o[22032] = i[43];
  assign o[22033] = i[43];
  assign o[22034] = i[43];
  assign o[22035] = i[43];
  assign o[22036] = i[43];
  assign o[22037] = i[43];
  assign o[22038] = i[43];
  assign o[22039] = i[43];
  assign o[22040] = i[43];
  assign o[22041] = i[43];
  assign o[22042] = i[43];
  assign o[22043] = i[43];
  assign o[22044] = i[43];
  assign o[22045] = i[43];
  assign o[22046] = i[43];
  assign o[22047] = i[43];
  assign o[22048] = i[43];
  assign o[22049] = i[43];
  assign o[22050] = i[43];
  assign o[22051] = i[43];
  assign o[22052] = i[43];
  assign o[22053] = i[43];
  assign o[22054] = i[43];
  assign o[22055] = i[43];
  assign o[22056] = i[43];
  assign o[22057] = i[43];
  assign o[22058] = i[43];
  assign o[22059] = i[43];
  assign o[22060] = i[43];
  assign o[22061] = i[43];
  assign o[22062] = i[43];
  assign o[22063] = i[43];
  assign o[22064] = i[43];
  assign o[22065] = i[43];
  assign o[22066] = i[43];
  assign o[22067] = i[43];
  assign o[22068] = i[43];
  assign o[22069] = i[43];
  assign o[22070] = i[43];
  assign o[22071] = i[43];
  assign o[22072] = i[43];
  assign o[22073] = i[43];
  assign o[22074] = i[43];
  assign o[22075] = i[43];
  assign o[22076] = i[43];
  assign o[22077] = i[43];
  assign o[22078] = i[43];
  assign o[22079] = i[43];
  assign o[22080] = i[43];
  assign o[22081] = i[43];
  assign o[22082] = i[43];
  assign o[22083] = i[43];
  assign o[22084] = i[43];
  assign o[22085] = i[43];
  assign o[22086] = i[43];
  assign o[22087] = i[43];
  assign o[22088] = i[43];
  assign o[22089] = i[43];
  assign o[22090] = i[43];
  assign o[22091] = i[43];
  assign o[22092] = i[43];
  assign o[22093] = i[43];
  assign o[22094] = i[43];
  assign o[22095] = i[43];
  assign o[22096] = i[43];
  assign o[22097] = i[43];
  assign o[22098] = i[43];
  assign o[22099] = i[43];
  assign o[22100] = i[43];
  assign o[22101] = i[43];
  assign o[22102] = i[43];
  assign o[22103] = i[43];
  assign o[22104] = i[43];
  assign o[22105] = i[43];
  assign o[22106] = i[43];
  assign o[22107] = i[43];
  assign o[22108] = i[43];
  assign o[22109] = i[43];
  assign o[22110] = i[43];
  assign o[22111] = i[43];
  assign o[22112] = i[43];
  assign o[22113] = i[43];
  assign o[22114] = i[43];
  assign o[22115] = i[43];
  assign o[22116] = i[43];
  assign o[22117] = i[43];
  assign o[22118] = i[43];
  assign o[22119] = i[43];
  assign o[22120] = i[43];
  assign o[22121] = i[43];
  assign o[22122] = i[43];
  assign o[22123] = i[43];
  assign o[22124] = i[43];
  assign o[22125] = i[43];
  assign o[22126] = i[43];
  assign o[22127] = i[43];
  assign o[22128] = i[43];
  assign o[22129] = i[43];
  assign o[22130] = i[43];
  assign o[22131] = i[43];
  assign o[22132] = i[43];
  assign o[22133] = i[43];
  assign o[22134] = i[43];
  assign o[22135] = i[43];
  assign o[22136] = i[43];
  assign o[22137] = i[43];
  assign o[22138] = i[43];
  assign o[22139] = i[43];
  assign o[22140] = i[43];
  assign o[22141] = i[43];
  assign o[22142] = i[43];
  assign o[22143] = i[43];
  assign o[22144] = i[43];
  assign o[22145] = i[43];
  assign o[22146] = i[43];
  assign o[22147] = i[43];
  assign o[22148] = i[43];
  assign o[22149] = i[43];
  assign o[22150] = i[43];
  assign o[22151] = i[43];
  assign o[22152] = i[43];
  assign o[22153] = i[43];
  assign o[22154] = i[43];
  assign o[22155] = i[43];
  assign o[22156] = i[43];
  assign o[22157] = i[43];
  assign o[22158] = i[43];
  assign o[22159] = i[43];
  assign o[22160] = i[43];
  assign o[22161] = i[43];
  assign o[22162] = i[43];
  assign o[22163] = i[43];
  assign o[22164] = i[43];
  assign o[22165] = i[43];
  assign o[22166] = i[43];
  assign o[22167] = i[43];
  assign o[22168] = i[43];
  assign o[22169] = i[43];
  assign o[22170] = i[43];
  assign o[22171] = i[43];
  assign o[22172] = i[43];
  assign o[22173] = i[43];
  assign o[22174] = i[43];
  assign o[22175] = i[43];
  assign o[22176] = i[43];
  assign o[22177] = i[43];
  assign o[22178] = i[43];
  assign o[22179] = i[43];
  assign o[22180] = i[43];
  assign o[22181] = i[43];
  assign o[22182] = i[43];
  assign o[22183] = i[43];
  assign o[22184] = i[43];
  assign o[22185] = i[43];
  assign o[22186] = i[43];
  assign o[22187] = i[43];
  assign o[22188] = i[43];
  assign o[22189] = i[43];
  assign o[22190] = i[43];
  assign o[22191] = i[43];
  assign o[22192] = i[43];
  assign o[22193] = i[43];
  assign o[22194] = i[43];
  assign o[22195] = i[43];
  assign o[22196] = i[43];
  assign o[22197] = i[43];
  assign o[22198] = i[43];
  assign o[22199] = i[43];
  assign o[22200] = i[43];
  assign o[22201] = i[43];
  assign o[22202] = i[43];
  assign o[22203] = i[43];
  assign o[22204] = i[43];
  assign o[22205] = i[43];
  assign o[22206] = i[43];
  assign o[22207] = i[43];
  assign o[22208] = i[43];
  assign o[22209] = i[43];
  assign o[22210] = i[43];
  assign o[22211] = i[43];
  assign o[22212] = i[43];
  assign o[22213] = i[43];
  assign o[22214] = i[43];
  assign o[22215] = i[43];
  assign o[22216] = i[43];
  assign o[22217] = i[43];
  assign o[22218] = i[43];
  assign o[22219] = i[43];
  assign o[22220] = i[43];
  assign o[22221] = i[43];
  assign o[22222] = i[43];
  assign o[22223] = i[43];
  assign o[22224] = i[43];
  assign o[22225] = i[43];
  assign o[22226] = i[43];
  assign o[22227] = i[43];
  assign o[22228] = i[43];
  assign o[22229] = i[43];
  assign o[22230] = i[43];
  assign o[22231] = i[43];
  assign o[22232] = i[43];
  assign o[22233] = i[43];
  assign o[22234] = i[43];
  assign o[22235] = i[43];
  assign o[22236] = i[43];
  assign o[22237] = i[43];
  assign o[22238] = i[43];
  assign o[22239] = i[43];
  assign o[22240] = i[43];
  assign o[22241] = i[43];
  assign o[22242] = i[43];
  assign o[22243] = i[43];
  assign o[22244] = i[43];
  assign o[22245] = i[43];
  assign o[22246] = i[43];
  assign o[22247] = i[43];
  assign o[22248] = i[43];
  assign o[22249] = i[43];
  assign o[22250] = i[43];
  assign o[22251] = i[43];
  assign o[22252] = i[43];
  assign o[22253] = i[43];
  assign o[22254] = i[43];
  assign o[22255] = i[43];
  assign o[22256] = i[43];
  assign o[22257] = i[43];
  assign o[22258] = i[43];
  assign o[22259] = i[43];
  assign o[22260] = i[43];
  assign o[22261] = i[43];
  assign o[22262] = i[43];
  assign o[22263] = i[43];
  assign o[22264] = i[43];
  assign o[22265] = i[43];
  assign o[22266] = i[43];
  assign o[22267] = i[43];
  assign o[22268] = i[43];
  assign o[22269] = i[43];
  assign o[22270] = i[43];
  assign o[22271] = i[43];
  assign o[22272] = i[43];
  assign o[22273] = i[43];
  assign o[22274] = i[43];
  assign o[22275] = i[43];
  assign o[22276] = i[43];
  assign o[22277] = i[43];
  assign o[22278] = i[43];
  assign o[22279] = i[43];
  assign o[22280] = i[43];
  assign o[22281] = i[43];
  assign o[22282] = i[43];
  assign o[22283] = i[43];
  assign o[22284] = i[43];
  assign o[22285] = i[43];
  assign o[22286] = i[43];
  assign o[22287] = i[43];
  assign o[22288] = i[43];
  assign o[22289] = i[43];
  assign o[22290] = i[43];
  assign o[22291] = i[43];
  assign o[22292] = i[43];
  assign o[22293] = i[43];
  assign o[22294] = i[43];
  assign o[22295] = i[43];
  assign o[22296] = i[43];
  assign o[22297] = i[43];
  assign o[22298] = i[43];
  assign o[22299] = i[43];
  assign o[22300] = i[43];
  assign o[22301] = i[43];
  assign o[22302] = i[43];
  assign o[22303] = i[43];
  assign o[22304] = i[43];
  assign o[22305] = i[43];
  assign o[22306] = i[43];
  assign o[22307] = i[43];
  assign o[22308] = i[43];
  assign o[22309] = i[43];
  assign o[22310] = i[43];
  assign o[22311] = i[43];
  assign o[22312] = i[43];
  assign o[22313] = i[43];
  assign o[22314] = i[43];
  assign o[22315] = i[43];
  assign o[22316] = i[43];
  assign o[22317] = i[43];
  assign o[22318] = i[43];
  assign o[22319] = i[43];
  assign o[22320] = i[43];
  assign o[22321] = i[43];
  assign o[22322] = i[43];
  assign o[22323] = i[43];
  assign o[22324] = i[43];
  assign o[22325] = i[43];
  assign o[22326] = i[43];
  assign o[22327] = i[43];
  assign o[22328] = i[43];
  assign o[22329] = i[43];
  assign o[22330] = i[43];
  assign o[22331] = i[43];
  assign o[22332] = i[43];
  assign o[22333] = i[43];
  assign o[22334] = i[43];
  assign o[22335] = i[43];
  assign o[22336] = i[43];
  assign o[22337] = i[43];
  assign o[22338] = i[43];
  assign o[22339] = i[43];
  assign o[22340] = i[43];
  assign o[22341] = i[43];
  assign o[22342] = i[43];
  assign o[22343] = i[43];
  assign o[22344] = i[43];
  assign o[22345] = i[43];
  assign o[22346] = i[43];
  assign o[22347] = i[43];
  assign o[22348] = i[43];
  assign o[22349] = i[43];
  assign o[22350] = i[43];
  assign o[22351] = i[43];
  assign o[22352] = i[43];
  assign o[22353] = i[43];
  assign o[22354] = i[43];
  assign o[22355] = i[43];
  assign o[22356] = i[43];
  assign o[22357] = i[43];
  assign o[22358] = i[43];
  assign o[22359] = i[43];
  assign o[22360] = i[43];
  assign o[22361] = i[43];
  assign o[22362] = i[43];
  assign o[22363] = i[43];
  assign o[22364] = i[43];
  assign o[22365] = i[43];
  assign o[22366] = i[43];
  assign o[22367] = i[43];
  assign o[22368] = i[43];
  assign o[22369] = i[43];
  assign o[22370] = i[43];
  assign o[22371] = i[43];
  assign o[22372] = i[43];
  assign o[22373] = i[43];
  assign o[22374] = i[43];
  assign o[22375] = i[43];
  assign o[22376] = i[43];
  assign o[22377] = i[43];
  assign o[22378] = i[43];
  assign o[22379] = i[43];
  assign o[22380] = i[43];
  assign o[22381] = i[43];
  assign o[22382] = i[43];
  assign o[22383] = i[43];
  assign o[22384] = i[43];
  assign o[22385] = i[43];
  assign o[22386] = i[43];
  assign o[22387] = i[43];
  assign o[22388] = i[43];
  assign o[22389] = i[43];
  assign o[22390] = i[43];
  assign o[22391] = i[43];
  assign o[22392] = i[43];
  assign o[22393] = i[43];
  assign o[22394] = i[43];
  assign o[22395] = i[43];
  assign o[22396] = i[43];
  assign o[22397] = i[43];
  assign o[22398] = i[43];
  assign o[22399] = i[43];
  assign o[22400] = i[43];
  assign o[22401] = i[43];
  assign o[22402] = i[43];
  assign o[22403] = i[43];
  assign o[22404] = i[43];
  assign o[22405] = i[43];
  assign o[22406] = i[43];
  assign o[22407] = i[43];
  assign o[22408] = i[43];
  assign o[22409] = i[43];
  assign o[22410] = i[43];
  assign o[22411] = i[43];
  assign o[22412] = i[43];
  assign o[22413] = i[43];
  assign o[22414] = i[43];
  assign o[22415] = i[43];
  assign o[22416] = i[43];
  assign o[22417] = i[43];
  assign o[22418] = i[43];
  assign o[22419] = i[43];
  assign o[22420] = i[43];
  assign o[22421] = i[43];
  assign o[22422] = i[43];
  assign o[22423] = i[43];
  assign o[22424] = i[43];
  assign o[22425] = i[43];
  assign o[22426] = i[43];
  assign o[22427] = i[43];
  assign o[22428] = i[43];
  assign o[22429] = i[43];
  assign o[22430] = i[43];
  assign o[22431] = i[43];
  assign o[22432] = i[43];
  assign o[22433] = i[43];
  assign o[22434] = i[43];
  assign o[22435] = i[43];
  assign o[22436] = i[43];
  assign o[22437] = i[43];
  assign o[22438] = i[43];
  assign o[22439] = i[43];
  assign o[22440] = i[43];
  assign o[22441] = i[43];
  assign o[22442] = i[43];
  assign o[22443] = i[43];
  assign o[22444] = i[43];
  assign o[22445] = i[43];
  assign o[22446] = i[43];
  assign o[22447] = i[43];
  assign o[22448] = i[43];
  assign o[22449] = i[43];
  assign o[22450] = i[43];
  assign o[22451] = i[43];
  assign o[22452] = i[43];
  assign o[22453] = i[43];
  assign o[22454] = i[43];
  assign o[22455] = i[43];
  assign o[22456] = i[43];
  assign o[22457] = i[43];
  assign o[22458] = i[43];
  assign o[22459] = i[43];
  assign o[22460] = i[43];
  assign o[22461] = i[43];
  assign o[22462] = i[43];
  assign o[22463] = i[43];
  assign o[22464] = i[43];
  assign o[22465] = i[43];
  assign o[22466] = i[43];
  assign o[22467] = i[43];
  assign o[22468] = i[43];
  assign o[22469] = i[43];
  assign o[22470] = i[43];
  assign o[22471] = i[43];
  assign o[22472] = i[43];
  assign o[22473] = i[43];
  assign o[22474] = i[43];
  assign o[22475] = i[43];
  assign o[22476] = i[43];
  assign o[22477] = i[43];
  assign o[22478] = i[43];
  assign o[22479] = i[43];
  assign o[22480] = i[43];
  assign o[22481] = i[43];
  assign o[22482] = i[43];
  assign o[22483] = i[43];
  assign o[22484] = i[43];
  assign o[22485] = i[43];
  assign o[22486] = i[43];
  assign o[22487] = i[43];
  assign o[22488] = i[43];
  assign o[22489] = i[43];
  assign o[22490] = i[43];
  assign o[22491] = i[43];
  assign o[22492] = i[43];
  assign o[22493] = i[43];
  assign o[22494] = i[43];
  assign o[22495] = i[43];
  assign o[22496] = i[43];
  assign o[22497] = i[43];
  assign o[22498] = i[43];
  assign o[22499] = i[43];
  assign o[22500] = i[43];
  assign o[22501] = i[43];
  assign o[22502] = i[43];
  assign o[22503] = i[43];
  assign o[22504] = i[43];
  assign o[22505] = i[43];
  assign o[22506] = i[43];
  assign o[22507] = i[43];
  assign o[22508] = i[43];
  assign o[22509] = i[43];
  assign o[22510] = i[43];
  assign o[22511] = i[43];
  assign o[22512] = i[43];
  assign o[22513] = i[43];
  assign o[22514] = i[43];
  assign o[22515] = i[43];
  assign o[22516] = i[43];
  assign o[22517] = i[43];
  assign o[22518] = i[43];
  assign o[22519] = i[43];
  assign o[22520] = i[43];
  assign o[22521] = i[43];
  assign o[22522] = i[43];
  assign o[22523] = i[43];
  assign o[22524] = i[43];
  assign o[22525] = i[43];
  assign o[22526] = i[43];
  assign o[22527] = i[43];
  assign o[21504] = i[42];
  assign o[21505] = i[42];
  assign o[21506] = i[42];
  assign o[21507] = i[42];
  assign o[21508] = i[42];
  assign o[21509] = i[42];
  assign o[21510] = i[42];
  assign o[21511] = i[42];
  assign o[21512] = i[42];
  assign o[21513] = i[42];
  assign o[21514] = i[42];
  assign o[21515] = i[42];
  assign o[21516] = i[42];
  assign o[21517] = i[42];
  assign o[21518] = i[42];
  assign o[21519] = i[42];
  assign o[21520] = i[42];
  assign o[21521] = i[42];
  assign o[21522] = i[42];
  assign o[21523] = i[42];
  assign o[21524] = i[42];
  assign o[21525] = i[42];
  assign o[21526] = i[42];
  assign o[21527] = i[42];
  assign o[21528] = i[42];
  assign o[21529] = i[42];
  assign o[21530] = i[42];
  assign o[21531] = i[42];
  assign o[21532] = i[42];
  assign o[21533] = i[42];
  assign o[21534] = i[42];
  assign o[21535] = i[42];
  assign o[21536] = i[42];
  assign o[21537] = i[42];
  assign o[21538] = i[42];
  assign o[21539] = i[42];
  assign o[21540] = i[42];
  assign o[21541] = i[42];
  assign o[21542] = i[42];
  assign o[21543] = i[42];
  assign o[21544] = i[42];
  assign o[21545] = i[42];
  assign o[21546] = i[42];
  assign o[21547] = i[42];
  assign o[21548] = i[42];
  assign o[21549] = i[42];
  assign o[21550] = i[42];
  assign o[21551] = i[42];
  assign o[21552] = i[42];
  assign o[21553] = i[42];
  assign o[21554] = i[42];
  assign o[21555] = i[42];
  assign o[21556] = i[42];
  assign o[21557] = i[42];
  assign o[21558] = i[42];
  assign o[21559] = i[42];
  assign o[21560] = i[42];
  assign o[21561] = i[42];
  assign o[21562] = i[42];
  assign o[21563] = i[42];
  assign o[21564] = i[42];
  assign o[21565] = i[42];
  assign o[21566] = i[42];
  assign o[21567] = i[42];
  assign o[21568] = i[42];
  assign o[21569] = i[42];
  assign o[21570] = i[42];
  assign o[21571] = i[42];
  assign o[21572] = i[42];
  assign o[21573] = i[42];
  assign o[21574] = i[42];
  assign o[21575] = i[42];
  assign o[21576] = i[42];
  assign o[21577] = i[42];
  assign o[21578] = i[42];
  assign o[21579] = i[42];
  assign o[21580] = i[42];
  assign o[21581] = i[42];
  assign o[21582] = i[42];
  assign o[21583] = i[42];
  assign o[21584] = i[42];
  assign o[21585] = i[42];
  assign o[21586] = i[42];
  assign o[21587] = i[42];
  assign o[21588] = i[42];
  assign o[21589] = i[42];
  assign o[21590] = i[42];
  assign o[21591] = i[42];
  assign o[21592] = i[42];
  assign o[21593] = i[42];
  assign o[21594] = i[42];
  assign o[21595] = i[42];
  assign o[21596] = i[42];
  assign o[21597] = i[42];
  assign o[21598] = i[42];
  assign o[21599] = i[42];
  assign o[21600] = i[42];
  assign o[21601] = i[42];
  assign o[21602] = i[42];
  assign o[21603] = i[42];
  assign o[21604] = i[42];
  assign o[21605] = i[42];
  assign o[21606] = i[42];
  assign o[21607] = i[42];
  assign o[21608] = i[42];
  assign o[21609] = i[42];
  assign o[21610] = i[42];
  assign o[21611] = i[42];
  assign o[21612] = i[42];
  assign o[21613] = i[42];
  assign o[21614] = i[42];
  assign o[21615] = i[42];
  assign o[21616] = i[42];
  assign o[21617] = i[42];
  assign o[21618] = i[42];
  assign o[21619] = i[42];
  assign o[21620] = i[42];
  assign o[21621] = i[42];
  assign o[21622] = i[42];
  assign o[21623] = i[42];
  assign o[21624] = i[42];
  assign o[21625] = i[42];
  assign o[21626] = i[42];
  assign o[21627] = i[42];
  assign o[21628] = i[42];
  assign o[21629] = i[42];
  assign o[21630] = i[42];
  assign o[21631] = i[42];
  assign o[21632] = i[42];
  assign o[21633] = i[42];
  assign o[21634] = i[42];
  assign o[21635] = i[42];
  assign o[21636] = i[42];
  assign o[21637] = i[42];
  assign o[21638] = i[42];
  assign o[21639] = i[42];
  assign o[21640] = i[42];
  assign o[21641] = i[42];
  assign o[21642] = i[42];
  assign o[21643] = i[42];
  assign o[21644] = i[42];
  assign o[21645] = i[42];
  assign o[21646] = i[42];
  assign o[21647] = i[42];
  assign o[21648] = i[42];
  assign o[21649] = i[42];
  assign o[21650] = i[42];
  assign o[21651] = i[42];
  assign o[21652] = i[42];
  assign o[21653] = i[42];
  assign o[21654] = i[42];
  assign o[21655] = i[42];
  assign o[21656] = i[42];
  assign o[21657] = i[42];
  assign o[21658] = i[42];
  assign o[21659] = i[42];
  assign o[21660] = i[42];
  assign o[21661] = i[42];
  assign o[21662] = i[42];
  assign o[21663] = i[42];
  assign o[21664] = i[42];
  assign o[21665] = i[42];
  assign o[21666] = i[42];
  assign o[21667] = i[42];
  assign o[21668] = i[42];
  assign o[21669] = i[42];
  assign o[21670] = i[42];
  assign o[21671] = i[42];
  assign o[21672] = i[42];
  assign o[21673] = i[42];
  assign o[21674] = i[42];
  assign o[21675] = i[42];
  assign o[21676] = i[42];
  assign o[21677] = i[42];
  assign o[21678] = i[42];
  assign o[21679] = i[42];
  assign o[21680] = i[42];
  assign o[21681] = i[42];
  assign o[21682] = i[42];
  assign o[21683] = i[42];
  assign o[21684] = i[42];
  assign o[21685] = i[42];
  assign o[21686] = i[42];
  assign o[21687] = i[42];
  assign o[21688] = i[42];
  assign o[21689] = i[42];
  assign o[21690] = i[42];
  assign o[21691] = i[42];
  assign o[21692] = i[42];
  assign o[21693] = i[42];
  assign o[21694] = i[42];
  assign o[21695] = i[42];
  assign o[21696] = i[42];
  assign o[21697] = i[42];
  assign o[21698] = i[42];
  assign o[21699] = i[42];
  assign o[21700] = i[42];
  assign o[21701] = i[42];
  assign o[21702] = i[42];
  assign o[21703] = i[42];
  assign o[21704] = i[42];
  assign o[21705] = i[42];
  assign o[21706] = i[42];
  assign o[21707] = i[42];
  assign o[21708] = i[42];
  assign o[21709] = i[42];
  assign o[21710] = i[42];
  assign o[21711] = i[42];
  assign o[21712] = i[42];
  assign o[21713] = i[42];
  assign o[21714] = i[42];
  assign o[21715] = i[42];
  assign o[21716] = i[42];
  assign o[21717] = i[42];
  assign o[21718] = i[42];
  assign o[21719] = i[42];
  assign o[21720] = i[42];
  assign o[21721] = i[42];
  assign o[21722] = i[42];
  assign o[21723] = i[42];
  assign o[21724] = i[42];
  assign o[21725] = i[42];
  assign o[21726] = i[42];
  assign o[21727] = i[42];
  assign o[21728] = i[42];
  assign o[21729] = i[42];
  assign o[21730] = i[42];
  assign o[21731] = i[42];
  assign o[21732] = i[42];
  assign o[21733] = i[42];
  assign o[21734] = i[42];
  assign o[21735] = i[42];
  assign o[21736] = i[42];
  assign o[21737] = i[42];
  assign o[21738] = i[42];
  assign o[21739] = i[42];
  assign o[21740] = i[42];
  assign o[21741] = i[42];
  assign o[21742] = i[42];
  assign o[21743] = i[42];
  assign o[21744] = i[42];
  assign o[21745] = i[42];
  assign o[21746] = i[42];
  assign o[21747] = i[42];
  assign o[21748] = i[42];
  assign o[21749] = i[42];
  assign o[21750] = i[42];
  assign o[21751] = i[42];
  assign o[21752] = i[42];
  assign o[21753] = i[42];
  assign o[21754] = i[42];
  assign o[21755] = i[42];
  assign o[21756] = i[42];
  assign o[21757] = i[42];
  assign o[21758] = i[42];
  assign o[21759] = i[42];
  assign o[21760] = i[42];
  assign o[21761] = i[42];
  assign o[21762] = i[42];
  assign o[21763] = i[42];
  assign o[21764] = i[42];
  assign o[21765] = i[42];
  assign o[21766] = i[42];
  assign o[21767] = i[42];
  assign o[21768] = i[42];
  assign o[21769] = i[42];
  assign o[21770] = i[42];
  assign o[21771] = i[42];
  assign o[21772] = i[42];
  assign o[21773] = i[42];
  assign o[21774] = i[42];
  assign o[21775] = i[42];
  assign o[21776] = i[42];
  assign o[21777] = i[42];
  assign o[21778] = i[42];
  assign o[21779] = i[42];
  assign o[21780] = i[42];
  assign o[21781] = i[42];
  assign o[21782] = i[42];
  assign o[21783] = i[42];
  assign o[21784] = i[42];
  assign o[21785] = i[42];
  assign o[21786] = i[42];
  assign o[21787] = i[42];
  assign o[21788] = i[42];
  assign o[21789] = i[42];
  assign o[21790] = i[42];
  assign o[21791] = i[42];
  assign o[21792] = i[42];
  assign o[21793] = i[42];
  assign o[21794] = i[42];
  assign o[21795] = i[42];
  assign o[21796] = i[42];
  assign o[21797] = i[42];
  assign o[21798] = i[42];
  assign o[21799] = i[42];
  assign o[21800] = i[42];
  assign o[21801] = i[42];
  assign o[21802] = i[42];
  assign o[21803] = i[42];
  assign o[21804] = i[42];
  assign o[21805] = i[42];
  assign o[21806] = i[42];
  assign o[21807] = i[42];
  assign o[21808] = i[42];
  assign o[21809] = i[42];
  assign o[21810] = i[42];
  assign o[21811] = i[42];
  assign o[21812] = i[42];
  assign o[21813] = i[42];
  assign o[21814] = i[42];
  assign o[21815] = i[42];
  assign o[21816] = i[42];
  assign o[21817] = i[42];
  assign o[21818] = i[42];
  assign o[21819] = i[42];
  assign o[21820] = i[42];
  assign o[21821] = i[42];
  assign o[21822] = i[42];
  assign o[21823] = i[42];
  assign o[21824] = i[42];
  assign o[21825] = i[42];
  assign o[21826] = i[42];
  assign o[21827] = i[42];
  assign o[21828] = i[42];
  assign o[21829] = i[42];
  assign o[21830] = i[42];
  assign o[21831] = i[42];
  assign o[21832] = i[42];
  assign o[21833] = i[42];
  assign o[21834] = i[42];
  assign o[21835] = i[42];
  assign o[21836] = i[42];
  assign o[21837] = i[42];
  assign o[21838] = i[42];
  assign o[21839] = i[42];
  assign o[21840] = i[42];
  assign o[21841] = i[42];
  assign o[21842] = i[42];
  assign o[21843] = i[42];
  assign o[21844] = i[42];
  assign o[21845] = i[42];
  assign o[21846] = i[42];
  assign o[21847] = i[42];
  assign o[21848] = i[42];
  assign o[21849] = i[42];
  assign o[21850] = i[42];
  assign o[21851] = i[42];
  assign o[21852] = i[42];
  assign o[21853] = i[42];
  assign o[21854] = i[42];
  assign o[21855] = i[42];
  assign o[21856] = i[42];
  assign o[21857] = i[42];
  assign o[21858] = i[42];
  assign o[21859] = i[42];
  assign o[21860] = i[42];
  assign o[21861] = i[42];
  assign o[21862] = i[42];
  assign o[21863] = i[42];
  assign o[21864] = i[42];
  assign o[21865] = i[42];
  assign o[21866] = i[42];
  assign o[21867] = i[42];
  assign o[21868] = i[42];
  assign o[21869] = i[42];
  assign o[21870] = i[42];
  assign o[21871] = i[42];
  assign o[21872] = i[42];
  assign o[21873] = i[42];
  assign o[21874] = i[42];
  assign o[21875] = i[42];
  assign o[21876] = i[42];
  assign o[21877] = i[42];
  assign o[21878] = i[42];
  assign o[21879] = i[42];
  assign o[21880] = i[42];
  assign o[21881] = i[42];
  assign o[21882] = i[42];
  assign o[21883] = i[42];
  assign o[21884] = i[42];
  assign o[21885] = i[42];
  assign o[21886] = i[42];
  assign o[21887] = i[42];
  assign o[21888] = i[42];
  assign o[21889] = i[42];
  assign o[21890] = i[42];
  assign o[21891] = i[42];
  assign o[21892] = i[42];
  assign o[21893] = i[42];
  assign o[21894] = i[42];
  assign o[21895] = i[42];
  assign o[21896] = i[42];
  assign o[21897] = i[42];
  assign o[21898] = i[42];
  assign o[21899] = i[42];
  assign o[21900] = i[42];
  assign o[21901] = i[42];
  assign o[21902] = i[42];
  assign o[21903] = i[42];
  assign o[21904] = i[42];
  assign o[21905] = i[42];
  assign o[21906] = i[42];
  assign o[21907] = i[42];
  assign o[21908] = i[42];
  assign o[21909] = i[42];
  assign o[21910] = i[42];
  assign o[21911] = i[42];
  assign o[21912] = i[42];
  assign o[21913] = i[42];
  assign o[21914] = i[42];
  assign o[21915] = i[42];
  assign o[21916] = i[42];
  assign o[21917] = i[42];
  assign o[21918] = i[42];
  assign o[21919] = i[42];
  assign o[21920] = i[42];
  assign o[21921] = i[42];
  assign o[21922] = i[42];
  assign o[21923] = i[42];
  assign o[21924] = i[42];
  assign o[21925] = i[42];
  assign o[21926] = i[42];
  assign o[21927] = i[42];
  assign o[21928] = i[42];
  assign o[21929] = i[42];
  assign o[21930] = i[42];
  assign o[21931] = i[42];
  assign o[21932] = i[42];
  assign o[21933] = i[42];
  assign o[21934] = i[42];
  assign o[21935] = i[42];
  assign o[21936] = i[42];
  assign o[21937] = i[42];
  assign o[21938] = i[42];
  assign o[21939] = i[42];
  assign o[21940] = i[42];
  assign o[21941] = i[42];
  assign o[21942] = i[42];
  assign o[21943] = i[42];
  assign o[21944] = i[42];
  assign o[21945] = i[42];
  assign o[21946] = i[42];
  assign o[21947] = i[42];
  assign o[21948] = i[42];
  assign o[21949] = i[42];
  assign o[21950] = i[42];
  assign o[21951] = i[42];
  assign o[21952] = i[42];
  assign o[21953] = i[42];
  assign o[21954] = i[42];
  assign o[21955] = i[42];
  assign o[21956] = i[42];
  assign o[21957] = i[42];
  assign o[21958] = i[42];
  assign o[21959] = i[42];
  assign o[21960] = i[42];
  assign o[21961] = i[42];
  assign o[21962] = i[42];
  assign o[21963] = i[42];
  assign o[21964] = i[42];
  assign o[21965] = i[42];
  assign o[21966] = i[42];
  assign o[21967] = i[42];
  assign o[21968] = i[42];
  assign o[21969] = i[42];
  assign o[21970] = i[42];
  assign o[21971] = i[42];
  assign o[21972] = i[42];
  assign o[21973] = i[42];
  assign o[21974] = i[42];
  assign o[21975] = i[42];
  assign o[21976] = i[42];
  assign o[21977] = i[42];
  assign o[21978] = i[42];
  assign o[21979] = i[42];
  assign o[21980] = i[42];
  assign o[21981] = i[42];
  assign o[21982] = i[42];
  assign o[21983] = i[42];
  assign o[21984] = i[42];
  assign o[21985] = i[42];
  assign o[21986] = i[42];
  assign o[21987] = i[42];
  assign o[21988] = i[42];
  assign o[21989] = i[42];
  assign o[21990] = i[42];
  assign o[21991] = i[42];
  assign o[21992] = i[42];
  assign o[21993] = i[42];
  assign o[21994] = i[42];
  assign o[21995] = i[42];
  assign o[21996] = i[42];
  assign o[21997] = i[42];
  assign o[21998] = i[42];
  assign o[21999] = i[42];
  assign o[22000] = i[42];
  assign o[22001] = i[42];
  assign o[22002] = i[42];
  assign o[22003] = i[42];
  assign o[22004] = i[42];
  assign o[22005] = i[42];
  assign o[22006] = i[42];
  assign o[22007] = i[42];
  assign o[22008] = i[42];
  assign o[22009] = i[42];
  assign o[22010] = i[42];
  assign o[22011] = i[42];
  assign o[22012] = i[42];
  assign o[22013] = i[42];
  assign o[22014] = i[42];
  assign o[22015] = i[42];
  assign o[20992] = i[41];
  assign o[20993] = i[41];
  assign o[20994] = i[41];
  assign o[20995] = i[41];
  assign o[20996] = i[41];
  assign o[20997] = i[41];
  assign o[20998] = i[41];
  assign o[20999] = i[41];
  assign o[21000] = i[41];
  assign o[21001] = i[41];
  assign o[21002] = i[41];
  assign o[21003] = i[41];
  assign o[21004] = i[41];
  assign o[21005] = i[41];
  assign o[21006] = i[41];
  assign o[21007] = i[41];
  assign o[21008] = i[41];
  assign o[21009] = i[41];
  assign o[21010] = i[41];
  assign o[21011] = i[41];
  assign o[21012] = i[41];
  assign o[21013] = i[41];
  assign o[21014] = i[41];
  assign o[21015] = i[41];
  assign o[21016] = i[41];
  assign o[21017] = i[41];
  assign o[21018] = i[41];
  assign o[21019] = i[41];
  assign o[21020] = i[41];
  assign o[21021] = i[41];
  assign o[21022] = i[41];
  assign o[21023] = i[41];
  assign o[21024] = i[41];
  assign o[21025] = i[41];
  assign o[21026] = i[41];
  assign o[21027] = i[41];
  assign o[21028] = i[41];
  assign o[21029] = i[41];
  assign o[21030] = i[41];
  assign o[21031] = i[41];
  assign o[21032] = i[41];
  assign o[21033] = i[41];
  assign o[21034] = i[41];
  assign o[21035] = i[41];
  assign o[21036] = i[41];
  assign o[21037] = i[41];
  assign o[21038] = i[41];
  assign o[21039] = i[41];
  assign o[21040] = i[41];
  assign o[21041] = i[41];
  assign o[21042] = i[41];
  assign o[21043] = i[41];
  assign o[21044] = i[41];
  assign o[21045] = i[41];
  assign o[21046] = i[41];
  assign o[21047] = i[41];
  assign o[21048] = i[41];
  assign o[21049] = i[41];
  assign o[21050] = i[41];
  assign o[21051] = i[41];
  assign o[21052] = i[41];
  assign o[21053] = i[41];
  assign o[21054] = i[41];
  assign o[21055] = i[41];
  assign o[21056] = i[41];
  assign o[21057] = i[41];
  assign o[21058] = i[41];
  assign o[21059] = i[41];
  assign o[21060] = i[41];
  assign o[21061] = i[41];
  assign o[21062] = i[41];
  assign o[21063] = i[41];
  assign o[21064] = i[41];
  assign o[21065] = i[41];
  assign o[21066] = i[41];
  assign o[21067] = i[41];
  assign o[21068] = i[41];
  assign o[21069] = i[41];
  assign o[21070] = i[41];
  assign o[21071] = i[41];
  assign o[21072] = i[41];
  assign o[21073] = i[41];
  assign o[21074] = i[41];
  assign o[21075] = i[41];
  assign o[21076] = i[41];
  assign o[21077] = i[41];
  assign o[21078] = i[41];
  assign o[21079] = i[41];
  assign o[21080] = i[41];
  assign o[21081] = i[41];
  assign o[21082] = i[41];
  assign o[21083] = i[41];
  assign o[21084] = i[41];
  assign o[21085] = i[41];
  assign o[21086] = i[41];
  assign o[21087] = i[41];
  assign o[21088] = i[41];
  assign o[21089] = i[41];
  assign o[21090] = i[41];
  assign o[21091] = i[41];
  assign o[21092] = i[41];
  assign o[21093] = i[41];
  assign o[21094] = i[41];
  assign o[21095] = i[41];
  assign o[21096] = i[41];
  assign o[21097] = i[41];
  assign o[21098] = i[41];
  assign o[21099] = i[41];
  assign o[21100] = i[41];
  assign o[21101] = i[41];
  assign o[21102] = i[41];
  assign o[21103] = i[41];
  assign o[21104] = i[41];
  assign o[21105] = i[41];
  assign o[21106] = i[41];
  assign o[21107] = i[41];
  assign o[21108] = i[41];
  assign o[21109] = i[41];
  assign o[21110] = i[41];
  assign o[21111] = i[41];
  assign o[21112] = i[41];
  assign o[21113] = i[41];
  assign o[21114] = i[41];
  assign o[21115] = i[41];
  assign o[21116] = i[41];
  assign o[21117] = i[41];
  assign o[21118] = i[41];
  assign o[21119] = i[41];
  assign o[21120] = i[41];
  assign o[21121] = i[41];
  assign o[21122] = i[41];
  assign o[21123] = i[41];
  assign o[21124] = i[41];
  assign o[21125] = i[41];
  assign o[21126] = i[41];
  assign o[21127] = i[41];
  assign o[21128] = i[41];
  assign o[21129] = i[41];
  assign o[21130] = i[41];
  assign o[21131] = i[41];
  assign o[21132] = i[41];
  assign o[21133] = i[41];
  assign o[21134] = i[41];
  assign o[21135] = i[41];
  assign o[21136] = i[41];
  assign o[21137] = i[41];
  assign o[21138] = i[41];
  assign o[21139] = i[41];
  assign o[21140] = i[41];
  assign o[21141] = i[41];
  assign o[21142] = i[41];
  assign o[21143] = i[41];
  assign o[21144] = i[41];
  assign o[21145] = i[41];
  assign o[21146] = i[41];
  assign o[21147] = i[41];
  assign o[21148] = i[41];
  assign o[21149] = i[41];
  assign o[21150] = i[41];
  assign o[21151] = i[41];
  assign o[21152] = i[41];
  assign o[21153] = i[41];
  assign o[21154] = i[41];
  assign o[21155] = i[41];
  assign o[21156] = i[41];
  assign o[21157] = i[41];
  assign o[21158] = i[41];
  assign o[21159] = i[41];
  assign o[21160] = i[41];
  assign o[21161] = i[41];
  assign o[21162] = i[41];
  assign o[21163] = i[41];
  assign o[21164] = i[41];
  assign o[21165] = i[41];
  assign o[21166] = i[41];
  assign o[21167] = i[41];
  assign o[21168] = i[41];
  assign o[21169] = i[41];
  assign o[21170] = i[41];
  assign o[21171] = i[41];
  assign o[21172] = i[41];
  assign o[21173] = i[41];
  assign o[21174] = i[41];
  assign o[21175] = i[41];
  assign o[21176] = i[41];
  assign o[21177] = i[41];
  assign o[21178] = i[41];
  assign o[21179] = i[41];
  assign o[21180] = i[41];
  assign o[21181] = i[41];
  assign o[21182] = i[41];
  assign o[21183] = i[41];
  assign o[21184] = i[41];
  assign o[21185] = i[41];
  assign o[21186] = i[41];
  assign o[21187] = i[41];
  assign o[21188] = i[41];
  assign o[21189] = i[41];
  assign o[21190] = i[41];
  assign o[21191] = i[41];
  assign o[21192] = i[41];
  assign o[21193] = i[41];
  assign o[21194] = i[41];
  assign o[21195] = i[41];
  assign o[21196] = i[41];
  assign o[21197] = i[41];
  assign o[21198] = i[41];
  assign o[21199] = i[41];
  assign o[21200] = i[41];
  assign o[21201] = i[41];
  assign o[21202] = i[41];
  assign o[21203] = i[41];
  assign o[21204] = i[41];
  assign o[21205] = i[41];
  assign o[21206] = i[41];
  assign o[21207] = i[41];
  assign o[21208] = i[41];
  assign o[21209] = i[41];
  assign o[21210] = i[41];
  assign o[21211] = i[41];
  assign o[21212] = i[41];
  assign o[21213] = i[41];
  assign o[21214] = i[41];
  assign o[21215] = i[41];
  assign o[21216] = i[41];
  assign o[21217] = i[41];
  assign o[21218] = i[41];
  assign o[21219] = i[41];
  assign o[21220] = i[41];
  assign o[21221] = i[41];
  assign o[21222] = i[41];
  assign o[21223] = i[41];
  assign o[21224] = i[41];
  assign o[21225] = i[41];
  assign o[21226] = i[41];
  assign o[21227] = i[41];
  assign o[21228] = i[41];
  assign o[21229] = i[41];
  assign o[21230] = i[41];
  assign o[21231] = i[41];
  assign o[21232] = i[41];
  assign o[21233] = i[41];
  assign o[21234] = i[41];
  assign o[21235] = i[41];
  assign o[21236] = i[41];
  assign o[21237] = i[41];
  assign o[21238] = i[41];
  assign o[21239] = i[41];
  assign o[21240] = i[41];
  assign o[21241] = i[41];
  assign o[21242] = i[41];
  assign o[21243] = i[41];
  assign o[21244] = i[41];
  assign o[21245] = i[41];
  assign o[21246] = i[41];
  assign o[21247] = i[41];
  assign o[21248] = i[41];
  assign o[21249] = i[41];
  assign o[21250] = i[41];
  assign o[21251] = i[41];
  assign o[21252] = i[41];
  assign o[21253] = i[41];
  assign o[21254] = i[41];
  assign o[21255] = i[41];
  assign o[21256] = i[41];
  assign o[21257] = i[41];
  assign o[21258] = i[41];
  assign o[21259] = i[41];
  assign o[21260] = i[41];
  assign o[21261] = i[41];
  assign o[21262] = i[41];
  assign o[21263] = i[41];
  assign o[21264] = i[41];
  assign o[21265] = i[41];
  assign o[21266] = i[41];
  assign o[21267] = i[41];
  assign o[21268] = i[41];
  assign o[21269] = i[41];
  assign o[21270] = i[41];
  assign o[21271] = i[41];
  assign o[21272] = i[41];
  assign o[21273] = i[41];
  assign o[21274] = i[41];
  assign o[21275] = i[41];
  assign o[21276] = i[41];
  assign o[21277] = i[41];
  assign o[21278] = i[41];
  assign o[21279] = i[41];
  assign o[21280] = i[41];
  assign o[21281] = i[41];
  assign o[21282] = i[41];
  assign o[21283] = i[41];
  assign o[21284] = i[41];
  assign o[21285] = i[41];
  assign o[21286] = i[41];
  assign o[21287] = i[41];
  assign o[21288] = i[41];
  assign o[21289] = i[41];
  assign o[21290] = i[41];
  assign o[21291] = i[41];
  assign o[21292] = i[41];
  assign o[21293] = i[41];
  assign o[21294] = i[41];
  assign o[21295] = i[41];
  assign o[21296] = i[41];
  assign o[21297] = i[41];
  assign o[21298] = i[41];
  assign o[21299] = i[41];
  assign o[21300] = i[41];
  assign o[21301] = i[41];
  assign o[21302] = i[41];
  assign o[21303] = i[41];
  assign o[21304] = i[41];
  assign o[21305] = i[41];
  assign o[21306] = i[41];
  assign o[21307] = i[41];
  assign o[21308] = i[41];
  assign o[21309] = i[41];
  assign o[21310] = i[41];
  assign o[21311] = i[41];
  assign o[21312] = i[41];
  assign o[21313] = i[41];
  assign o[21314] = i[41];
  assign o[21315] = i[41];
  assign o[21316] = i[41];
  assign o[21317] = i[41];
  assign o[21318] = i[41];
  assign o[21319] = i[41];
  assign o[21320] = i[41];
  assign o[21321] = i[41];
  assign o[21322] = i[41];
  assign o[21323] = i[41];
  assign o[21324] = i[41];
  assign o[21325] = i[41];
  assign o[21326] = i[41];
  assign o[21327] = i[41];
  assign o[21328] = i[41];
  assign o[21329] = i[41];
  assign o[21330] = i[41];
  assign o[21331] = i[41];
  assign o[21332] = i[41];
  assign o[21333] = i[41];
  assign o[21334] = i[41];
  assign o[21335] = i[41];
  assign o[21336] = i[41];
  assign o[21337] = i[41];
  assign o[21338] = i[41];
  assign o[21339] = i[41];
  assign o[21340] = i[41];
  assign o[21341] = i[41];
  assign o[21342] = i[41];
  assign o[21343] = i[41];
  assign o[21344] = i[41];
  assign o[21345] = i[41];
  assign o[21346] = i[41];
  assign o[21347] = i[41];
  assign o[21348] = i[41];
  assign o[21349] = i[41];
  assign o[21350] = i[41];
  assign o[21351] = i[41];
  assign o[21352] = i[41];
  assign o[21353] = i[41];
  assign o[21354] = i[41];
  assign o[21355] = i[41];
  assign o[21356] = i[41];
  assign o[21357] = i[41];
  assign o[21358] = i[41];
  assign o[21359] = i[41];
  assign o[21360] = i[41];
  assign o[21361] = i[41];
  assign o[21362] = i[41];
  assign o[21363] = i[41];
  assign o[21364] = i[41];
  assign o[21365] = i[41];
  assign o[21366] = i[41];
  assign o[21367] = i[41];
  assign o[21368] = i[41];
  assign o[21369] = i[41];
  assign o[21370] = i[41];
  assign o[21371] = i[41];
  assign o[21372] = i[41];
  assign o[21373] = i[41];
  assign o[21374] = i[41];
  assign o[21375] = i[41];
  assign o[21376] = i[41];
  assign o[21377] = i[41];
  assign o[21378] = i[41];
  assign o[21379] = i[41];
  assign o[21380] = i[41];
  assign o[21381] = i[41];
  assign o[21382] = i[41];
  assign o[21383] = i[41];
  assign o[21384] = i[41];
  assign o[21385] = i[41];
  assign o[21386] = i[41];
  assign o[21387] = i[41];
  assign o[21388] = i[41];
  assign o[21389] = i[41];
  assign o[21390] = i[41];
  assign o[21391] = i[41];
  assign o[21392] = i[41];
  assign o[21393] = i[41];
  assign o[21394] = i[41];
  assign o[21395] = i[41];
  assign o[21396] = i[41];
  assign o[21397] = i[41];
  assign o[21398] = i[41];
  assign o[21399] = i[41];
  assign o[21400] = i[41];
  assign o[21401] = i[41];
  assign o[21402] = i[41];
  assign o[21403] = i[41];
  assign o[21404] = i[41];
  assign o[21405] = i[41];
  assign o[21406] = i[41];
  assign o[21407] = i[41];
  assign o[21408] = i[41];
  assign o[21409] = i[41];
  assign o[21410] = i[41];
  assign o[21411] = i[41];
  assign o[21412] = i[41];
  assign o[21413] = i[41];
  assign o[21414] = i[41];
  assign o[21415] = i[41];
  assign o[21416] = i[41];
  assign o[21417] = i[41];
  assign o[21418] = i[41];
  assign o[21419] = i[41];
  assign o[21420] = i[41];
  assign o[21421] = i[41];
  assign o[21422] = i[41];
  assign o[21423] = i[41];
  assign o[21424] = i[41];
  assign o[21425] = i[41];
  assign o[21426] = i[41];
  assign o[21427] = i[41];
  assign o[21428] = i[41];
  assign o[21429] = i[41];
  assign o[21430] = i[41];
  assign o[21431] = i[41];
  assign o[21432] = i[41];
  assign o[21433] = i[41];
  assign o[21434] = i[41];
  assign o[21435] = i[41];
  assign o[21436] = i[41];
  assign o[21437] = i[41];
  assign o[21438] = i[41];
  assign o[21439] = i[41];
  assign o[21440] = i[41];
  assign o[21441] = i[41];
  assign o[21442] = i[41];
  assign o[21443] = i[41];
  assign o[21444] = i[41];
  assign o[21445] = i[41];
  assign o[21446] = i[41];
  assign o[21447] = i[41];
  assign o[21448] = i[41];
  assign o[21449] = i[41];
  assign o[21450] = i[41];
  assign o[21451] = i[41];
  assign o[21452] = i[41];
  assign o[21453] = i[41];
  assign o[21454] = i[41];
  assign o[21455] = i[41];
  assign o[21456] = i[41];
  assign o[21457] = i[41];
  assign o[21458] = i[41];
  assign o[21459] = i[41];
  assign o[21460] = i[41];
  assign o[21461] = i[41];
  assign o[21462] = i[41];
  assign o[21463] = i[41];
  assign o[21464] = i[41];
  assign o[21465] = i[41];
  assign o[21466] = i[41];
  assign o[21467] = i[41];
  assign o[21468] = i[41];
  assign o[21469] = i[41];
  assign o[21470] = i[41];
  assign o[21471] = i[41];
  assign o[21472] = i[41];
  assign o[21473] = i[41];
  assign o[21474] = i[41];
  assign o[21475] = i[41];
  assign o[21476] = i[41];
  assign o[21477] = i[41];
  assign o[21478] = i[41];
  assign o[21479] = i[41];
  assign o[21480] = i[41];
  assign o[21481] = i[41];
  assign o[21482] = i[41];
  assign o[21483] = i[41];
  assign o[21484] = i[41];
  assign o[21485] = i[41];
  assign o[21486] = i[41];
  assign o[21487] = i[41];
  assign o[21488] = i[41];
  assign o[21489] = i[41];
  assign o[21490] = i[41];
  assign o[21491] = i[41];
  assign o[21492] = i[41];
  assign o[21493] = i[41];
  assign o[21494] = i[41];
  assign o[21495] = i[41];
  assign o[21496] = i[41];
  assign o[21497] = i[41];
  assign o[21498] = i[41];
  assign o[21499] = i[41];
  assign o[21500] = i[41];
  assign o[21501] = i[41];
  assign o[21502] = i[41];
  assign o[21503] = i[41];
  assign o[20480] = i[40];
  assign o[20481] = i[40];
  assign o[20482] = i[40];
  assign o[20483] = i[40];
  assign o[20484] = i[40];
  assign o[20485] = i[40];
  assign o[20486] = i[40];
  assign o[20487] = i[40];
  assign o[20488] = i[40];
  assign o[20489] = i[40];
  assign o[20490] = i[40];
  assign o[20491] = i[40];
  assign o[20492] = i[40];
  assign o[20493] = i[40];
  assign o[20494] = i[40];
  assign o[20495] = i[40];
  assign o[20496] = i[40];
  assign o[20497] = i[40];
  assign o[20498] = i[40];
  assign o[20499] = i[40];
  assign o[20500] = i[40];
  assign o[20501] = i[40];
  assign o[20502] = i[40];
  assign o[20503] = i[40];
  assign o[20504] = i[40];
  assign o[20505] = i[40];
  assign o[20506] = i[40];
  assign o[20507] = i[40];
  assign o[20508] = i[40];
  assign o[20509] = i[40];
  assign o[20510] = i[40];
  assign o[20511] = i[40];
  assign o[20512] = i[40];
  assign o[20513] = i[40];
  assign o[20514] = i[40];
  assign o[20515] = i[40];
  assign o[20516] = i[40];
  assign o[20517] = i[40];
  assign o[20518] = i[40];
  assign o[20519] = i[40];
  assign o[20520] = i[40];
  assign o[20521] = i[40];
  assign o[20522] = i[40];
  assign o[20523] = i[40];
  assign o[20524] = i[40];
  assign o[20525] = i[40];
  assign o[20526] = i[40];
  assign o[20527] = i[40];
  assign o[20528] = i[40];
  assign o[20529] = i[40];
  assign o[20530] = i[40];
  assign o[20531] = i[40];
  assign o[20532] = i[40];
  assign o[20533] = i[40];
  assign o[20534] = i[40];
  assign o[20535] = i[40];
  assign o[20536] = i[40];
  assign o[20537] = i[40];
  assign o[20538] = i[40];
  assign o[20539] = i[40];
  assign o[20540] = i[40];
  assign o[20541] = i[40];
  assign o[20542] = i[40];
  assign o[20543] = i[40];
  assign o[20544] = i[40];
  assign o[20545] = i[40];
  assign o[20546] = i[40];
  assign o[20547] = i[40];
  assign o[20548] = i[40];
  assign o[20549] = i[40];
  assign o[20550] = i[40];
  assign o[20551] = i[40];
  assign o[20552] = i[40];
  assign o[20553] = i[40];
  assign o[20554] = i[40];
  assign o[20555] = i[40];
  assign o[20556] = i[40];
  assign o[20557] = i[40];
  assign o[20558] = i[40];
  assign o[20559] = i[40];
  assign o[20560] = i[40];
  assign o[20561] = i[40];
  assign o[20562] = i[40];
  assign o[20563] = i[40];
  assign o[20564] = i[40];
  assign o[20565] = i[40];
  assign o[20566] = i[40];
  assign o[20567] = i[40];
  assign o[20568] = i[40];
  assign o[20569] = i[40];
  assign o[20570] = i[40];
  assign o[20571] = i[40];
  assign o[20572] = i[40];
  assign o[20573] = i[40];
  assign o[20574] = i[40];
  assign o[20575] = i[40];
  assign o[20576] = i[40];
  assign o[20577] = i[40];
  assign o[20578] = i[40];
  assign o[20579] = i[40];
  assign o[20580] = i[40];
  assign o[20581] = i[40];
  assign o[20582] = i[40];
  assign o[20583] = i[40];
  assign o[20584] = i[40];
  assign o[20585] = i[40];
  assign o[20586] = i[40];
  assign o[20587] = i[40];
  assign o[20588] = i[40];
  assign o[20589] = i[40];
  assign o[20590] = i[40];
  assign o[20591] = i[40];
  assign o[20592] = i[40];
  assign o[20593] = i[40];
  assign o[20594] = i[40];
  assign o[20595] = i[40];
  assign o[20596] = i[40];
  assign o[20597] = i[40];
  assign o[20598] = i[40];
  assign o[20599] = i[40];
  assign o[20600] = i[40];
  assign o[20601] = i[40];
  assign o[20602] = i[40];
  assign o[20603] = i[40];
  assign o[20604] = i[40];
  assign o[20605] = i[40];
  assign o[20606] = i[40];
  assign o[20607] = i[40];
  assign o[20608] = i[40];
  assign o[20609] = i[40];
  assign o[20610] = i[40];
  assign o[20611] = i[40];
  assign o[20612] = i[40];
  assign o[20613] = i[40];
  assign o[20614] = i[40];
  assign o[20615] = i[40];
  assign o[20616] = i[40];
  assign o[20617] = i[40];
  assign o[20618] = i[40];
  assign o[20619] = i[40];
  assign o[20620] = i[40];
  assign o[20621] = i[40];
  assign o[20622] = i[40];
  assign o[20623] = i[40];
  assign o[20624] = i[40];
  assign o[20625] = i[40];
  assign o[20626] = i[40];
  assign o[20627] = i[40];
  assign o[20628] = i[40];
  assign o[20629] = i[40];
  assign o[20630] = i[40];
  assign o[20631] = i[40];
  assign o[20632] = i[40];
  assign o[20633] = i[40];
  assign o[20634] = i[40];
  assign o[20635] = i[40];
  assign o[20636] = i[40];
  assign o[20637] = i[40];
  assign o[20638] = i[40];
  assign o[20639] = i[40];
  assign o[20640] = i[40];
  assign o[20641] = i[40];
  assign o[20642] = i[40];
  assign o[20643] = i[40];
  assign o[20644] = i[40];
  assign o[20645] = i[40];
  assign o[20646] = i[40];
  assign o[20647] = i[40];
  assign o[20648] = i[40];
  assign o[20649] = i[40];
  assign o[20650] = i[40];
  assign o[20651] = i[40];
  assign o[20652] = i[40];
  assign o[20653] = i[40];
  assign o[20654] = i[40];
  assign o[20655] = i[40];
  assign o[20656] = i[40];
  assign o[20657] = i[40];
  assign o[20658] = i[40];
  assign o[20659] = i[40];
  assign o[20660] = i[40];
  assign o[20661] = i[40];
  assign o[20662] = i[40];
  assign o[20663] = i[40];
  assign o[20664] = i[40];
  assign o[20665] = i[40];
  assign o[20666] = i[40];
  assign o[20667] = i[40];
  assign o[20668] = i[40];
  assign o[20669] = i[40];
  assign o[20670] = i[40];
  assign o[20671] = i[40];
  assign o[20672] = i[40];
  assign o[20673] = i[40];
  assign o[20674] = i[40];
  assign o[20675] = i[40];
  assign o[20676] = i[40];
  assign o[20677] = i[40];
  assign o[20678] = i[40];
  assign o[20679] = i[40];
  assign o[20680] = i[40];
  assign o[20681] = i[40];
  assign o[20682] = i[40];
  assign o[20683] = i[40];
  assign o[20684] = i[40];
  assign o[20685] = i[40];
  assign o[20686] = i[40];
  assign o[20687] = i[40];
  assign o[20688] = i[40];
  assign o[20689] = i[40];
  assign o[20690] = i[40];
  assign o[20691] = i[40];
  assign o[20692] = i[40];
  assign o[20693] = i[40];
  assign o[20694] = i[40];
  assign o[20695] = i[40];
  assign o[20696] = i[40];
  assign o[20697] = i[40];
  assign o[20698] = i[40];
  assign o[20699] = i[40];
  assign o[20700] = i[40];
  assign o[20701] = i[40];
  assign o[20702] = i[40];
  assign o[20703] = i[40];
  assign o[20704] = i[40];
  assign o[20705] = i[40];
  assign o[20706] = i[40];
  assign o[20707] = i[40];
  assign o[20708] = i[40];
  assign o[20709] = i[40];
  assign o[20710] = i[40];
  assign o[20711] = i[40];
  assign o[20712] = i[40];
  assign o[20713] = i[40];
  assign o[20714] = i[40];
  assign o[20715] = i[40];
  assign o[20716] = i[40];
  assign o[20717] = i[40];
  assign o[20718] = i[40];
  assign o[20719] = i[40];
  assign o[20720] = i[40];
  assign o[20721] = i[40];
  assign o[20722] = i[40];
  assign o[20723] = i[40];
  assign o[20724] = i[40];
  assign o[20725] = i[40];
  assign o[20726] = i[40];
  assign o[20727] = i[40];
  assign o[20728] = i[40];
  assign o[20729] = i[40];
  assign o[20730] = i[40];
  assign o[20731] = i[40];
  assign o[20732] = i[40];
  assign o[20733] = i[40];
  assign o[20734] = i[40];
  assign o[20735] = i[40];
  assign o[20736] = i[40];
  assign o[20737] = i[40];
  assign o[20738] = i[40];
  assign o[20739] = i[40];
  assign o[20740] = i[40];
  assign o[20741] = i[40];
  assign o[20742] = i[40];
  assign o[20743] = i[40];
  assign o[20744] = i[40];
  assign o[20745] = i[40];
  assign o[20746] = i[40];
  assign o[20747] = i[40];
  assign o[20748] = i[40];
  assign o[20749] = i[40];
  assign o[20750] = i[40];
  assign o[20751] = i[40];
  assign o[20752] = i[40];
  assign o[20753] = i[40];
  assign o[20754] = i[40];
  assign o[20755] = i[40];
  assign o[20756] = i[40];
  assign o[20757] = i[40];
  assign o[20758] = i[40];
  assign o[20759] = i[40];
  assign o[20760] = i[40];
  assign o[20761] = i[40];
  assign o[20762] = i[40];
  assign o[20763] = i[40];
  assign o[20764] = i[40];
  assign o[20765] = i[40];
  assign o[20766] = i[40];
  assign o[20767] = i[40];
  assign o[20768] = i[40];
  assign o[20769] = i[40];
  assign o[20770] = i[40];
  assign o[20771] = i[40];
  assign o[20772] = i[40];
  assign o[20773] = i[40];
  assign o[20774] = i[40];
  assign o[20775] = i[40];
  assign o[20776] = i[40];
  assign o[20777] = i[40];
  assign o[20778] = i[40];
  assign o[20779] = i[40];
  assign o[20780] = i[40];
  assign o[20781] = i[40];
  assign o[20782] = i[40];
  assign o[20783] = i[40];
  assign o[20784] = i[40];
  assign o[20785] = i[40];
  assign o[20786] = i[40];
  assign o[20787] = i[40];
  assign o[20788] = i[40];
  assign o[20789] = i[40];
  assign o[20790] = i[40];
  assign o[20791] = i[40];
  assign o[20792] = i[40];
  assign o[20793] = i[40];
  assign o[20794] = i[40];
  assign o[20795] = i[40];
  assign o[20796] = i[40];
  assign o[20797] = i[40];
  assign o[20798] = i[40];
  assign o[20799] = i[40];
  assign o[20800] = i[40];
  assign o[20801] = i[40];
  assign o[20802] = i[40];
  assign o[20803] = i[40];
  assign o[20804] = i[40];
  assign o[20805] = i[40];
  assign o[20806] = i[40];
  assign o[20807] = i[40];
  assign o[20808] = i[40];
  assign o[20809] = i[40];
  assign o[20810] = i[40];
  assign o[20811] = i[40];
  assign o[20812] = i[40];
  assign o[20813] = i[40];
  assign o[20814] = i[40];
  assign o[20815] = i[40];
  assign o[20816] = i[40];
  assign o[20817] = i[40];
  assign o[20818] = i[40];
  assign o[20819] = i[40];
  assign o[20820] = i[40];
  assign o[20821] = i[40];
  assign o[20822] = i[40];
  assign o[20823] = i[40];
  assign o[20824] = i[40];
  assign o[20825] = i[40];
  assign o[20826] = i[40];
  assign o[20827] = i[40];
  assign o[20828] = i[40];
  assign o[20829] = i[40];
  assign o[20830] = i[40];
  assign o[20831] = i[40];
  assign o[20832] = i[40];
  assign o[20833] = i[40];
  assign o[20834] = i[40];
  assign o[20835] = i[40];
  assign o[20836] = i[40];
  assign o[20837] = i[40];
  assign o[20838] = i[40];
  assign o[20839] = i[40];
  assign o[20840] = i[40];
  assign o[20841] = i[40];
  assign o[20842] = i[40];
  assign o[20843] = i[40];
  assign o[20844] = i[40];
  assign o[20845] = i[40];
  assign o[20846] = i[40];
  assign o[20847] = i[40];
  assign o[20848] = i[40];
  assign o[20849] = i[40];
  assign o[20850] = i[40];
  assign o[20851] = i[40];
  assign o[20852] = i[40];
  assign o[20853] = i[40];
  assign o[20854] = i[40];
  assign o[20855] = i[40];
  assign o[20856] = i[40];
  assign o[20857] = i[40];
  assign o[20858] = i[40];
  assign o[20859] = i[40];
  assign o[20860] = i[40];
  assign o[20861] = i[40];
  assign o[20862] = i[40];
  assign o[20863] = i[40];
  assign o[20864] = i[40];
  assign o[20865] = i[40];
  assign o[20866] = i[40];
  assign o[20867] = i[40];
  assign o[20868] = i[40];
  assign o[20869] = i[40];
  assign o[20870] = i[40];
  assign o[20871] = i[40];
  assign o[20872] = i[40];
  assign o[20873] = i[40];
  assign o[20874] = i[40];
  assign o[20875] = i[40];
  assign o[20876] = i[40];
  assign o[20877] = i[40];
  assign o[20878] = i[40];
  assign o[20879] = i[40];
  assign o[20880] = i[40];
  assign o[20881] = i[40];
  assign o[20882] = i[40];
  assign o[20883] = i[40];
  assign o[20884] = i[40];
  assign o[20885] = i[40];
  assign o[20886] = i[40];
  assign o[20887] = i[40];
  assign o[20888] = i[40];
  assign o[20889] = i[40];
  assign o[20890] = i[40];
  assign o[20891] = i[40];
  assign o[20892] = i[40];
  assign o[20893] = i[40];
  assign o[20894] = i[40];
  assign o[20895] = i[40];
  assign o[20896] = i[40];
  assign o[20897] = i[40];
  assign o[20898] = i[40];
  assign o[20899] = i[40];
  assign o[20900] = i[40];
  assign o[20901] = i[40];
  assign o[20902] = i[40];
  assign o[20903] = i[40];
  assign o[20904] = i[40];
  assign o[20905] = i[40];
  assign o[20906] = i[40];
  assign o[20907] = i[40];
  assign o[20908] = i[40];
  assign o[20909] = i[40];
  assign o[20910] = i[40];
  assign o[20911] = i[40];
  assign o[20912] = i[40];
  assign o[20913] = i[40];
  assign o[20914] = i[40];
  assign o[20915] = i[40];
  assign o[20916] = i[40];
  assign o[20917] = i[40];
  assign o[20918] = i[40];
  assign o[20919] = i[40];
  assign o[20920] = i[40];
  assign o[20921] = i[40];
  assign o[20922] = i[40];
  assign o[20923] = i[40];
  assign o[20924] = i[40];
  assign o[20925] = i[40];
  assign o[20926] = i[40];
  assign o[20927] = i[40];
  assign o[20928] = i[40];
  assign o[20929] = i[40];
  assign o[20930] = i[40];
  assign o[20931] = i[40];
  assign o[20932] = i[40];
  assign o[20933] = i[40];
  assign o[20934] = i[40];
  assign o[20935] = i[40];
  assign o[20936] = i[40];
  assign o[20937] = i[40];
  assign o[20938] = i[40];
  assign o[20939] = i[40];
  assign o[20940] = i[40];
  assign o[20941] = i[40];
  assign o[20942] = i[40];
  assign o[20943] = i[40];
  assign o[20944] = i[40];
  assign o[20945] = i[40];
  assign o[20946] = i[40];
  assign o[20947] = i[40];
  assign o[20948] = i[40];
  assign o[20949] = i[40];
  assign o[20950] = i[40];
  assign o[20951] = i[40];
  assign o[20952] = i[40];
  assign o[20953] = i[40];
  assign o[20954] = i[40];
  assign o[20955] = i[40];
  assign o[20956] = i[40];
  assign o[20957] = i[40];
  assign o[20958] = i[40];
  assign o[20959] = i[40];
  assign o[20960] = i[40];
  assign o[20961] = i[40];
  assign o[20962] = i[40];
  assign o[20963] = i[40];
  assign o[20964] = i[40];
  assign o[20965] = i[40];
  assign o[20966] = i[40];
  assign o[20967] = i[40];
  assign o[20968] = i[40];
  assign o[20969] = i[40];
  assign o[20970] = i[40];
  assign o[20971] = i[40];
  assign o[20972] = i[40];
  assign o[20973] = i[40];
  assign o[20974] = i[40];
  assign o[20975] = i[40];
  assign o[20976] = i[40];
  assign o[20977] = i[40];
  assign o[20978] = i[40];
  assign o[20979] = i[40];
  assign o[20980] = i[40];
  assign o[20981] = i[40];
  assign o[20982] = i[40];
  assign o[20983] = i[40];
  assign o[20984] = i[40];
  assign o[20985] = i[40];
  assign o[20986] = i[40];
  assign o[20987] = i[40];
  assign o[20988] = i[40];
  assign o[20989] = i[40];
  assign o[20990] = i[40];
  assign o[20991] = i[40];
  assign o[19968] = i[39];
  assign o[19969] = i[39];
  assign o[19970] = i[39];
  assign o[19971] = i[39];
  assign o[19972] = i[39];
  assign o[19973] = i[39];
  assign o[19974] = i[39];
  assign o[19975] = i[39];
  assign o[19976] = i[39];
  assign o[19977] = i[39];
  assign o[19978] = i[39];
  assign o[19979] = i[39];
  assign o[19980] = i[39];
  assign o[19981] = i[39];
  assign o[19982] = i[39];
  assign o[19983] = i[39];
  assign o[19984] = i[39];
  assign o[19985] = i[39];
  assign o[19986] = i[39];
  assign o[19987] = i[39];
  assign o[19988] = i[39];
  assign o[19989] = i[39];
  assign o[19990] = i[39];
  assign o[19991] = i[39];
  assign o[19992] = i[39];
  assign o[19993] = i[39];
  assign o[19994] = i[39];
  assign o[19995] = i[39];
  assign o[19996] = i[39];
  assign o[19997] = i[39];
  assign o[19998] = i[39];
  assign o[19999] = i[39];
  assign o[20000] = i[39];
  assign o[20001] = i[39];
  assign o[20002] = i[39];
  assign o[20003] = i[39];
  assign o[20004] = i[39];
  assign o[20005] = i[39];
  assign o[20006] = i[39];
  assign o[20007] = i[39];
  assign o[20008] = i[39];
  assign o[20009] = i[39];
  assign o[20010] = i[39];
  assign o[20011] = i[39];
  assign o[20012] = i[39];
  assign o[20013] = i[39];
  assign o[20014] = i[39];
  assign o[20015] = i[39];
  assign o[20016] = i[39];
  assign o[20017] = i[39];
  assign o[20018] = i[39];
  assign o[20019] = i[39];
  assign o[20020] = i[39];
  assign o[20021] = i[39];
  assign o[20022] = i[39];
  assign o[20023] = i[39];
  assign o[20024] = i[39];
  assign o[20025] = i[39];
  assign o[20026] = i[39];
  assign o[20027] = i[39];
  assign o[20028] = i[39];
  assign o[20029] = i[39];
  assign o[20030] = i[39];
  assign o[20031] = i[39];
  assign o[20032] = i[39];
  assign o[20033] = i[39];
  assign o[20034] = i[39];
  assign o[20035] = i[39];
  assign o[20036] = i[39];
  assign o[20037] = i[39];
  assign o[20038] = i[39];
  assign o[20039] = i[39];
  assign o[20040] = i[39];
  assign o[20041] = i[39];
  assign o[20042] = i[39];
  assign o[20043] = i[39];
  assign o[20044] = i[39];
  assign o[20045] = i[39];
  assign o[20046] = i[39];
  assign o[20047] = i[39];
  assign o[20048] = i[39];
  assign o[20049] = i[39];
  assign o[20050] = i[39];
  assign o[20051] = i[39];
  assign o[20052] = i[39];
  assign o[20053] = i[39];
  assign o[20054] = i[39];
  assign o[20055] = i[39];
  assign o[20056] = i[39];
  assign o[20057] = i[39];
  assign o[20058] = i[39];
  assign o[20059] = i[39];
  assign o[20060] = i[39];
  assign o[20061] = i[39];
  assign o[20062] = i[39];
  assign o[20063] = i[39];
  assign o[20064] = i[39];
  assign o[20065] = i[39];
  assign o[20066] = i[39];
  assign o[20067] = i[39];
  assign o[20068] = i[39];
  assign o[20069] = i[39];
  assign o[20070] = i[39];
  assign o[20071] = i[39];
  assign o[20072] = i[39];
  assign o[20073] = i[39];
  assign o[20074] = i[39];
  assign o[20075] = i[39];
  assign o[20076] = i[39];
  assign o[20077] = i[39];
  assign o[20078] = i[39];
  assign o[20079] = i[39];
  assign o[20080] = i[39];
  assign o[20081] = i[39];
  assign o[20082] = i[39];
  assign o[20083] = i[39];
  assign o[20084] = i[39];
  assign o[20085] = i[39];
  assign o[20086] = i[39];
  assign o[20087] = i[39];
  assign o[20088] = i[39];
  assign o[20089] = i[39];
  assign o[20090] = i[39];
  assign o[20091] = i[39];
  assign o[20092] = i[39];
  assign o[20093] = i[39];
  assign o[20094] = i[39];
  assign o[20095] = i[39];
  assign o[20096] = i[39];
  assign o[20097] = i[39];
  assign o[20098] = i[39];
  assign o[20099] = i[39];
  assign o[20100] = i[39];
  assign o[20101] = i[39];
  assign o[20102] = i[39];
  assign o[20103] = i[39];
  assign o[20104] = i[39];
  assign o[20105] = i[39];
  assign o[20106] = i[39];
  assign o[20107] = i[39];
  assign o[20108] = i[39];
  assign o[20109] = i[39];
  assign o[20110] = i[39];
  assign o[20111] = i[39];
  assign o[20112] = i[39];
  assign o[20113] = i[39];
  assign o[20114] = i[39];
  assign o[20115] = i[39];
  assign o[20116] = i[39];
  assign o[20117] = i[39];
  assign o[20118] = i[39];
  assign o[20119] = i[39];
  assign o[20120] = i[39];
  assign o[20121] = i[39];
  assign o[20122] = i[39];
  assign o[20123] = i[39];
  assign o[20124] = i[39];
  assign o[20125] = i[39];
  assign o[20126] = i[39];
  assign o[20127] = i[39];
  assign o[20128] = i[39];
  assign o[20129] = i[39];
  assign o[20130] = i[39];
  assign o[20131] = i[39];
  assign o[20132] = i[39];
  assign o[20133] = i[39];
  assign o[20134] = i[39];
  assign o[20135] = i[39];
  assign o[20136] = i[39];
  assign o[20137] = i[39];
  assign o[20138] = i[39];
  assign o[20139] = i[39];
  assign o[20140] = i[39];
  assign o[20141] = i[39];
  assign o[20142] = i[39];
  assign o[20143] = i[39];
  assign o[20144] = i[39];
  assign o[20145] = i[39];
  assign o[20146] = i[39];
  assign o[20147] = i[39];
  assign o[20148] = i[39];
  assign o[20149] = i[39];
  assign o[20150] = i[39];
  assign o[20151] = i[39];
  assign o[20152] = i[39];
  assign o[20153] = i[39];
  assign o[20154] = i[39];
  assign o[20155] = i[39];
  assign o[20156] = i[39];
  assign o[20157] = i[39];
  assign o[20158] = i[39];
  assign o[20159] = i[39];
  assign o[20160] = i[39];
  assign o[20161] = i[39];
  assign o[20162] = i[39];
  assign o[20163] = i[39];
  assign o[20164] = i[39];
  assign o[20165] = i[39];
  assign o[20166] = i[39];
  assign o[20167] = i[39];
  assign o[20168] = i[39];
  assign o[20169] = i[39];
  assign o[20170] = i[39];
  assign o[20171] = i[39];
  assign o[20172] = i[39];
  assign o[20173] = i[39];
  assign o[20174] = i[39];
  assign o[20175] = i[39];
  assign o[20176] = i[39];
  assign o[20177] = i[39];
  assign o[20178] = i[39];
  assign o[20179] = i[39];
  assign o[20180] = i[39];
  assign o[20181] = i[39];
  assign o[20182] = i[39];
  assign o[20183] = i[39];
  assign o[20184] = i[39];
  assign o[20185] = i[39];
  assign o[20186] = i[39];
  assign o[20187] = i[39];
  assign o[20188] = i[39];
  assign o[20189] = i[39];
  assign o[20190] = i[39];
  assign o[20191] = i[39];
  assign o[20192] = i[39];
  assign o[20193] = i[39];
  assign o[20194] = i[39];
  assign o[20195] = i[39];
  assign o[20196] = i[39];
  assign o[20197] = i[39];
  assign o[20198] = i[39];
  assign o[20199] = i[39];
  assign o[20200] = i[39];
  assign o[20201] = i[39];
  assign o[20202] = i[39];
  assign o[20203] = i[39];
  assign o[20204] = i[39];
  assign o[20205] = i[39];
  assign o[20206] = i[39];
  assign o[20207] = i[39];
  assign o[20208] = i[39];
  assign o[20209] = i[39];
  assign o[20210] = i[39];
  assign o[20211] = i[39];
  assign o[20212] = i[39];
  assign o[20213] = i[39];
  assign o[20214] = i[39];
  assign o[20215] = i[39];
  assign o[20216] = i[39];
  assign o[20217] = i[39];
  assign o[20218] = i[39];
  assign o[20219] = i[39];
  assign o[20220] = i[39];
  assign o[20221] = i[39];
  assign o[20222] = i[39];
  assign o[20223] = i[39];
  assign o[20224] = i[39];
  assign o[20225] = i[39];
  assign o[20226] = i[39];
  assign o[20227] = i[39];
  assign o[20228] = i[39];
  assign o[20229] = i[39];
  assign o[20230] = i[39];
  assign o[20231] = i[39];
  assign o[20232] = i[39];
  assign o[20233] = i[39];
  assign o[20234] = i[39];
  assign o[20235] = i[39];
  assign o[20236] = i[39];
  assign o[20237] = i[39];
  assign o[20238] = i[39];
  assign o[20239] = i[39];
  assign o[20240] = i[39];
  assign o[20241] = i[39];
  assign o[20242] = i[39];
  assign o[20243] = i[39];
  assign o[20244] = i[39];
  assign o[20245] = i[39];
  assign o[20246] = i[39];
  assign o[20247] = i[39];
  assign o[20248] = i[39];
  assign o[20249] = i[39];
  assign o[20250] = i[39];
  assign o[20251] = i[39];
  assign o[20252] = i[39];
  assign o[20253] = i[39];
  assign o[20254] = i[39];
  assign o[20255] = i[39];
  assign o[20256] = i[39];
  assign o[20257] = i[39];
  assign o[20258] = i[39];
  assign o[20259] = i[39];
  assign o[20260] = i[39];
  assign o[20261] = i[39];
  assign o[20262] = i[39];
  assign o[20263] = i[39];
  assign o[20264] = i[39];
  assign o[20265] = i[39];
  assign o[20266] = i[39];
  assign o[20267] = i[39];
  assign o[20268] = i[39];
  assign o[20269] = i[39];
  assign o[20270] = i[39];
  assign o[20271] = i[39];
  assign o[20272] = i[39];
  assign o[20273] = i[39];
  assign o[20274] = i[39];
  assign o[20275] = i[39];
  assign o[20276] = i[39];
  assign o[20277] = i[39];
  assign o[20278] = i[39];
  assign o[20279] = i[39];
  assign o[20280] = i[39];
  assign o[20281] = i[39];
  assign o[20282] = i[39];
  assign o[20283] = i[39];
  assign o[20284] = i[39];
  assign o[20285] = i[39];
  assign o[20286] = i[39];
  assign o[20287] = i[39];
  assign o[20288] = i[39];
  assign o[20289] = i[39];
  assign o[20290] = i[39];
  assign o[20291] = i[39];
  assign o[20292] = i[39];
  assign o[20293] = i[39];
  assign o[20294] = i[39];
  assign o[20295] = i[39];
  assign o[20296] = i[39];
  assign o[20297] = i[39];
  assign o[20298] = i[39];
  assign o[20299] = i[39];
  assign o[20300] = i[39];
  assign o[20301] = i[39];
  assign o[20302] = i[39];
  assign o[20303] = i[39];
  assign o[20304] = i[39];
  assign o[20305] = i[39];
  assign o[20306] = i[39];
  assign o[20307] = i[39];
  assign o[20308] = i[39];
  assign o[20309] = i[39];
  assign o[20310] = i[39];
  assign o[20311] = i[39];
  assign o[20312] = i[39];
  assign o[20313] = i[39];
  assign o[20314] = i[39];
  assign o[20315] = i[39];
  assign o[20316] = i[39];
  assign o[20317] = i[39];
  assign o[20318] = i[39];
  assign o[20319] = i[39];
  assign o[20320] = i[39];
  assign o[20321] = i[39];
  assign o[20322] = i[39];
  assign o[20323] = i[39];
  assign o[20324] = i[39];
  assign o[20325] = i[39];
  assign o[20326] = i[39];
  assign o[20327] = i[39];
  assign o[20328] = i[39];
  assign o[20329] = i[39];
  assign o[20330] = i[39];
  assign o[20331] = i[39];
  assign o[20332] = i[39];
  assign o[20333] = i[39];
  assign o[20334] = i[39];
  assign o[20335] = i[39];
  assign o[20336] = i[39];
  assign o[20337] = i[39];
  assign o[20338] = i[39];
  assign o[20339] = i[39];
  assign o[20340] = i[39];
  assign o[20341] = i[39];
  assign o[20342] = i[39];
  assign o[20343] = i[39];
  assign o[20344] = i[39];
  assign o[20345] = i[39];
  assign o[20346] = i[39];
  assign o[20347] = i[39];
  assign o[20348] = i[39];
  assign o[20349] = i[39];
  assign o[20350] = i[39];
  assign o[20351] = i[39];
  assign o[20352] = i[39];
  assign o[20353] = i[39];
  assign o[20354] = i[39];
  assign o[20355] = i[39];
  assign o[20356] = i[39];
  assign o[20357] = i[39];
  assign o[20358] = i[39];
  assign o[20359] = i[39];
  assign o[20360] = i[39];
  assign o[20361] = i[39];
  assign o[20362] = i[39];
  assign o[20363] = i[39];
  assign o[20364] = i[39];
  assign o[20365] = i[39];
  assign o[20366] = i[39];
  assign o[20367] = i[39];
  assign o[20368] = i[39];
  assign o[20369] = i[39];
  assign o[20370] = i[39];
  assign o[20371] = i[39];
  assign o[20372] = i[39];
  assign o[20373] = i[39];
  assign o[20374] = i[39];
  assign o[20375] = i[39];
  assign o[20376] = i[39];
  assign o[20377] = i[39];
  assign o[20378] = i[39];
  assign o[20379] = i[39];
  assign o[20380] = i[39];
  assign o[20381] = i[39];
  assign o[20382] = i[39];
  assign o[20383] = i[39];
  assign o[20384] = i[39];
  assign o[20385] = i[39];
  assign o[20386] = i[39];
  assign o[20387] = i[39];
  assign o[20388] = i[39];
  assign o[20389] = i[39];
  assign o[20390] = i[39];
  assign o[20391] = i[39];
  assign o[20392] = i[39];
  assign o[20393] = i[39];
  assign o[20394] = i[39];
  assign o[20395] = i[39];
  assign o[20396] = i[39];
  assign o[20397] = i[39];
  assign o[20398] = i[39];
  assign o[20399] = i[39];
  assign o[20400] = i[39];
  assign o[20401] = i[39];
  assign o[20402] = i[39];
  assign o[20403] = i[39];
  assign o[20404] = i[39];
  assign o[20405] = i[39];
  assign o[20406] = i[39];
  assign o[20407] = i[39];
  assign o[20408] = i[39];
  assign o[20409] = i[39];
  assign o[20410] = i[39];
  assign o[20411] = i[39];
  assign o[20412] = i[39];
  assign o[20413] = i[39];
  assign o[20414] = i[39];
  assign o[20415] = i[39];
  assign o[20416] = i[39];
  assign o[20417] = i[39];
  assign o[20418] = i[39];
  assign o[20419] = i[39];
  assign o[20420] = i[39];
  assign o[20421] = i[39];
  assign o[20422] = i[39];
  assign o[20423] = i[39];
  assign o[20424] = i[39];
  assign o[20425] = i[39];
  assign o[20426] = i[39];
  assign o[20427] = i[39];
  assign o[20428] = i[39];
  assign o[20429] = i[39];
  assign o[20430] = i[39];
  assign o[20431] = i[39];
  assign o[20432] = i[39];
  assign o[20433] = i[39];
  assign o[20434] = i[39];
  assign o[20435] = i[39];
  assign o[20436] = i[39];
  assign o[20437] = i[39];
  assign o[20438] = i[39];
  assign o[20439] = i[39];
  assign o[20440] = i[39];
  assign o[20441] = i[39];
  assign o[20442] = i[39];
  assign o[20443] = i[39];
  assign o[20444] = i[39];
  assign o[20445] = i[39];
  assign o[20446] = i[39];
  assign o[20447] = i[39];
  assign o[20448] = i[39];
  assign o[20449] = i[39];
  assign o[20450] = i[39];
  assign o[20451] = i[39];
  assign o[20452] = i[39];
  assign o[20453] = i[39];
  assign o[20454] = i[39];
  assign o[20455] = i[39];
  assign o[20456] = i[39];
  assign o[20457] = i[39];
  assign o[20458] = i[39];
  assign o[20459] = i[39];
  assign o[20460] = i[39];
  assign o[20461] = i[39];
  assign o[20462] = i[39];
  assign o[20463] = i[39];
  assign o[20464] = i[39];
  assign o[20465] = i[39];
  assign o[20466] = i[39];
  assign o[20467] = i[39];
  assign o[20468] = i[39];
  assign o[20469] = i[39];
  assign o[20470] = i[39];
  assign o[20471] = i[39];
  assign o[20472] = i[39];
  assign o[20473] = i[39];
  assign o[20474] = i[39];
  assign o[20475] = i[39];
  assign o[20476] = i[39];
  assign o[20477] = i[39];
  assign o[20478] = i[39];
  assign o[20479] = i[39];
  assign o[19456] = i[38];
  assign o[19457] = i[38];
  assign o[19458] = i[38];
  assign o[19459] = i[38];
  assign o[19460] = i[38];
  assign o[19461] = i[38];
  assign o[19462] = i[38];
  assign o[19463] = i[38];
  assign o[19464] = i[38];
  assign o[19465] = i[38];
  assign o[19466] = i[38];
  assign o[19467] = i[38];
  assign o[19468] = i[38];
  assign o[19469] = i[38];
  assign o[19470] = i[38];
  assign o[19471] = i[38];
  assign o[19472] = i[38];
  assign o[19473] = i[38];
  assign o[19474] = i[38];
  assign o[19475] = i[38];
  assign o[19476] = i[38];
  assign o[19477] = i[38];
  assign o[19478] = i[38];
  assign o[19479] = i[38];
  assign o[19480] = i[38];
  assign o[19481] = i[38];
  assign o[19482] = i[38];
  assign o[19483] = i[38];
  assign o[19484] = i[38];
  assign o[19485] = i[38];
  assign o[19486] = i[38];
  assign o[19487] = i[38];
  assign o[19488] = i[38];
  assign o[19489] = i[38];
  assign o[19490] = i[38];
  assign o[19491] = i[38];
  assign o[19492] = i[38];
  assign o[19493] = i[38];
  assign o[19494] = i[38];
  assign o[19495] = i[38];
  assign o[19496] = i[38];
  assign o[19497] = i[38];
  assign o[19498] = i[38];
  assign o[19499] = i[38];
  assign o[19500] = i[38];
  assign o[19501] = i[38];
  assign o[19502] = i[38];
  assign o[19503] = i[38];
  assign o[19504] = i[38];
  assign o[19505] = i[38];
  assign o[19506] = i[38];
  assign o[19507] = i[38];
  assign o[19508] = i[38];
  assign o[19509] = i[38];
  assign o[19510] = i[38];
  assign o[19511] = i[38];
  assign o[19512] = i[38];
  assign o[19513] = i[38];
  assign o[19514] = i[38];
  assign o[19515] = i[38];
  assign o[19516] = i[38];
  assign o[19517] = i[38];
  assign o[19518] = i[38];
  assign o[19519] = i[38];
  assign o[19520] = i[38];
  assign o[19521] = i[38];
  assign o[19522] = i[38];
  assign o[19523] = i[38];
  assign o[19524] = i[38];
  assign o[19525] = i[38];
  assign o[19526] = i[38];
  assign o[19527] = i[38];
  assign o[19528] = i[38];
  assign o[19529] = i[38];
  assign o[19530] = i[38];
  assign o[19531] = i[38];
  assign o[19532] = i[38];
  assign o[19533] = i[38];
  assign o[19534] = i[38];
  assign o[19535] = i[38];
  assign o[19536] = i[38];
  assign o[19537] = i[38];
  assign o[19538] = i[38];
  assign o[19539] = i[38];
  assign o[19540] = i[38];
  assign o[19541] = i[38];
  assign o[19542] = i[38];
  assign o[19543] = i[38];
  assign o[19544] = i[38];
  assign o[19545] = i[38];
  assign o[19546] = i[38];
  assign o[19547] = i[38];
  assign o[19548] = i[38];
  assign o[19549] = i[38];
  assign o[19550] = i[38];
  assign o[19551] = i[38];
  assign o[19552] = i[38];
  assign o[19553] = i[38];
  assign o[19554] = i[38];
  assign o[19555] = i[38];
  assign o[19556] = i[38];
  assign o[19557] = i[38];
  assign o[19558] = i[38];
  assign o[19559] = i[38];
  assign o[19560] = i[38];
  assign o[19561] = i[38];
  assign o[19562] = i[38];
  assign o[19563] = i[38];
  assign o[19564] = i[38];
  assign o[19565] = i[38];
  assign o[19566] = i[38];
  assign o[19567] = i[38];
  assign o[19568] = i[38];
  assign o[19569] = i[38];
  assign o[19570] = i[38];
  assign o[19571] = i[38];
  assign o[19572] = i[38];
  assign o[19573] = i[38];
  assign o[19574] = i[38];
  assign o[19575] = i[38];
  assign o[19576] = i[38];
  assign o[19577] = i[38];
  assign o[19578] = i[38];
  assign o[19579] = i[38];
  assign o[19580] = i[38];
  assign o[19581] = i[38];
  assign o[19582] = i[38];
  assign o[19583] = i[38];
  assign o[19584] = i[38];
  assign o[19585] = i[38];
  assign o[19586] = i[38];
  assign o[19587] = i[38];
  assign o[19588] = i[38];
  assign o[19589] = i[38];
  assign o[19590] = i[38];
  assign o[19591] = i[38];
  assign o[19592] = i[38];
  assign o[19593] = i[38];
  assign o[19594] = i[38];
  assign o[19595] = i[38];
  assign o[19596] = i[38];
  assign o[19597] = i[38];
  assign o[19598] = i[38];
  assign o[19599] = i[38];
  assign o[19600] = i[38];
  assign o[19601] = i[38];
  assign o[19602] = i[38];
  assign o[19603] = i[38];
  assign o[19604] = i[38];
  assign o[19605] = i[38];
  assign o[19606] = i[38];
  assign o[19607] = i[38];
  assign o[19608] = i[38];
  assign o[19609] = i[38];
  assign o[19610] = i[38];
  assign o[19611] = i[38];
  assign o[19612] = i[38];
  assign o[19613] = i[38];
  assign o[19614] = i[38];
  assign o[19615] = i[38];
  assign o[19616] = i[38];
  assign o[19617] = i[38];
  assign o[19618] = i[38];
  assign o[19619] = i[38];
  assign o[19620] = i[38];
  assign o[19621] = i[38];
  assign o[19622] = i[38];
  assign o[19623] = i[38];
  assign o[19624] = i[38];
  assign o[19625] = i[38];
  assign o[19626] = i[38];
  assign o[19627] = i[38];
  assign o[19628] = i[38];
  assign o[19629] = i[38];
  assign o[19630] = i[38];
  assign o[19631] = i[38];
  assign o[19632] = i[38];
  assign o[19633] = i[38];
  assign o[19634] = i[38];
  assign o[19635] = i[38];
  assign o[19636] = i[38];
  assign o[19637] = i[38];
  assign o[19638] = i[38];
  assign o[19639] = i[38];
  assign o[19640] = i[38];
  assign o[19641] = i[38];
  assign o[19642] = i[38];
  assign o[19643] = i[38];
  assign o[19644] = i[38];
  assign o[19645] = i[38];
  assign o[19646] = i[38];
  assign o[19647] = i[38];
  assign o[19648] = i[38];
  assign o[19649] = i[38];
  assign o[19650] = i[38];
  assign o[19651] = i[38];
  assign o[19652] = i[38];
  assign o[19653] = i[38];
  assign o[19654] = i[38];
  assign o[19655] = i[38];
  assign o[19656] = i[38];
  assign o[19657] = i[38];
  assign o[19658] = i[38];
  assign o[19659] = i[38];
  assign o[19660] = i[38];
  assign o[19661] = i[38];
  assign o[19662] = i[38];
  assign o[19663] = i[38];
  assign o[19664] = i[38];
  assign o[19665] = i[38];
  assign o[19666] = i[38];
  assign o[19667] = i[38];
  assign o[19668] = i[38];
  assign o[19669] = i[38];
  assign o[19670] = i[38];
  assign o[19671] = i[38];
  assign o[19672] = i[38];
  assign o[19673] = i[38];
  assign o[19674] = i[38];
  assign o[19675] = i[38];
  assign o[19676] = i[38];
  assign o[19677] = i[38];
  assign o[19678] = i[38];
  assign o[19679] = i[38];
  assign o[19680] = i[38];
  assign o[19681] = i[38];
  assign o[19682] = i[38];
  assign o[19683] = i[38];
  assign o[19684] = i[38];
  assign o[19685] = i[38];
  assign o[19686] = i[38];
  assign o[19687] = i[38];
  assign o[19688] = i[38];
  assign o[19689] = i[38];
  assign o[19690] = i[38];
  assign o[19691] = i[38];
  assign o[19692] = i[38];
  assign o[19693] = i[38];
  assign o[19694] = i[38];
  assign o[19695] = i[38];
  assign o[19696] = i[38];
  assign o[19697] = i[38];
  assign o[19698] = i[38];
  assign o[19699] = i[38];
  assign o[19700] = i[38];
  assign o[19701] = i[38];
  assign o[19702] = i[38];
  assign o[19703] = i[38];
  assign o[19704] = i[38];
  assign o[19705] = i[38];
  assign o[19706] = i[38];
  assign o[19707] = i[38];
  assign o[19708] = i[38];
  assign o[19709] = i[38];
  assign o[19710] = i[38];
  assign o[19711] = i[38];
  assign o[19712] = i[38];
  assign o[19713] = i[38];
  assign o[19714] = i[38];
  assign o[19715] = i[38];
  assign o[19716] = i[38];
  assign o[19717] = i[38];
  assign o[19718] = i[38];
  assign o[19719] = i[38];
  assign o[19720] = i[38];
  assign o[19721] = i[38];
  assign o[19722] = i[38];
  assign o[19723] = i[38];
  assign o[19724] = i[38];
  assign o[19725] = i[38];
  assign o[19726] = i[38];
  assign o[19727] = i[38];
  assign o[19728] = i[38];
  assign o[19729] = i[38];
  assign o[19730] = i[38];
  assign o[19731] = i[38];
  assign o[19732] = i[38];
  assign o[19733] = i[38];
  assign o[19734] = i[38];
  assign o[19735] = i[38];
  assign o[19736] = i[38];
  assign o[19737] = i[38];
  assign o[19738] = i[38];
  assign o[19739] = i[38];
  assign o[19740] = i[38];
  assign o[19741] = i[38];
  assign o[19742] = i[38];
  assign o[19743] = i[38];
  assign o[19744] = i[38];
  assign o[19745] = i[38];
  assign o[19746] = i[38];
  assign o[19747] = i[38];
  assign o[19748] = i[38];
  assign o[19749] = i[38];
  assign o[19750] = i[38];
  assign o[19751] = i[38];
  assign o[19752] = i[38];
  assign o[19753] = i[38];
  assign o[19754] = i[38];
  assign o[19755] = i[38];
  assign o[19756] = i[38];
  assign o[19757] = i[38];
  assign o[19758] = i[38];
  assign o[19759] = i[38];
  assign o[19760] = i[38];
  assign o[19761] = i[38];
  assign o[19762] = i[38];
  assign o[19763] = i[38];
  assign o[19764] = i[38];
  assign o[19765] = i[38];
  assign o[19766] = i[38];
  assign o[19767] = i[38];
  assign o[19768] = i[38];
  assign o[19769] = i[38];
  assign o[19770] = i[38];
  assign o[19771] = i[38];
  assign o[19772] = i[38];
  assign o[19773] = i[38];
  assign o[19774] = i[38];
  assign o[19775] = i[38];
  assign o[19776] = i[38];
  assign o[19777] = i[38];
  assign o[19778] = i[38];
  assign o[19779] = i[38];
  assign o[19780] = i[38];
  assign o[19781] = i[38];
  assign o[19782] = i[38];
  assign o[19783] = i[38];
  assign o[19784] = i[38];
  assign o[19785] = i[38];
  assign o[19786] = i[38];
  assign o[19787] = i[38];
  assign o[19788] = i[38];
  assign o[19789] = i[38];
  assign o[19790] = i[38];
  assign o[19791] = i[38];
  assign o[19792] = i[38];
  assign o[19793] = i[38];
  assign o[19794] = i[38];
  assign o[19795] = i[38];
  assign o[19796] = i[38];
  assign o[19797] = i[38];
  assign o[19798] = i[38];
  assign o[19799] = i[38];
  assign o[19800] = i[38];
  assign o[19801] = i[38];
  assign o[19802] = i[38];
  assign o[19803] = i[38];
  assign o[19804] = i[38];
  assign o[19805] = i[38];
  assign o[19806] = i[38];
  assign o[19807] = i[38];
  assign o[19808] = i[38];
  assign o[19809] = i[38];
  assign o[19810] = i[38];
  assign o[19811] = i[38];
  assign o[19812] = i[38];
  assign o[19813] = i[38];
  assign o[19814] = i[38];
  assign o[19815] = i[38];
  assign o[19816] = i[38];
  assign o[19817] = i[38];
  assign o[19818] = i[38];
  assign o[19819] = i[38];
  assign o[19820] = i[38];
  assign o[19821] = i[38];
  assign o[19822] = i[38];
  assign o[19823] = i[38];
  assign o[19824] = i[38];
  assign o[19825] = i[38];
  assign o[19826] = i[38];
  assign o[19827] = i[38];
  assign o[19828] = i[38];
  assign o[19829] = i[38];
  assign o[19830] = i[38];
  assign o[19831] = i[38];
  assign o[19832] = i[38];
  assign o[19833] = i[38];
  assign o[19834] = i[38];
  assign o[19835] = i[38];
  assign o[19836] = i[38];
  assign o[19837] = i[38];
  assign o[19838] = i[38];
  assign o[19839] = i[38];
  assign o[19840] = i[38];
  assign o[19841] = i[38];
  assign o[19842] = i[38];
  assign o[19843] = i[38];
  assign o[19844] = i[38];
  assign o[19845] = i[38];
  assign o[19846] = i[38];
  assign o[19847] = i[38];
  assign o[19848] = i[38];
  assign o[19849] = i[38];
  assign o[19850] = i[38];
  assign o[19851] = i[38];
  assign o[19852] = i[38];
  assign o[19853] = i[38];
  assign o[19854] = i[38];
  assign o[19855] = i[38];
  assign o[19856] = i[38];
  assign o[19857] = i[38];
  assign o[19858] = i[38];
  assign o[19859] = i[38];
  assign o[19860] = i[38];
  assign o[19861] = i[38];
  assign o[19862] = i[38];
  assign o[19863] = i[38];
  assign o[19864] = i[38];
  assign o[19865] = i[38];
  assign o[19866] = i[38];
  assign o[19867] = i[38];
  assign o[19868] = i[38];
  assign o[19869] = i[38];
  assign o[19870] = i[38];
  assign o[19871] = i[38];
  assign o[19872] = i[38];
  assign o[19873] = i[38];
  assign o[19874] = i[38];
  assign o[19875] = i[38];
  assign o[19876] = i[38];
  assign o[19877] = i[38];
  assign o[19878] = i[38];
  assign o[19879] = i[38];
  assign o[19880] = i[38];
  assign o[19881] = i[38];
  assign o[19882] = i[38];
  assign o[19883] = i[38];
  assign o[19884] = i[38];
  assign o[19885] = i[38];
  assign o[19886] = i[38];
  assign o[19887] = i[38];
  assign o[19888] = i[38];
  assign o[19889] = i[38];
  assign o[19890] = i[38];
  assign o[19891] = i[38];
  assign o[19892] = i[38];
  assign o[19893] = i[38];
  assign o[19894] = i[38];
  assign o[19895] = i[38];
  assign o[19896] = i[38];
  assign o[19897] = i[38];
  assign o[19898] = i[38];
  assign o[19899] = i[38];
  assign o[19900] = i[38];
  assign o[19901] = i[38];
  assign o[19902] = i[38];
  assign o[19903] = i[38];
  assign o[19904] = i[38];
  assign o[19905] = i[38];
  assign o[19906] = i[38];
  assign o[19907] = i[38];
  assign o[19908] = i[38];
  assign o[19909] = i[38];
  assign o[19910] = i[38];
  assign o[19911] = i[38];
  assign o[19912] = i[38];
  assign o[19913] = i[38];
  assign o[19914] = i[38];
  assign o[19915] = i[38];
  assign o[19916] = i[38];
  assign o[19917] = i[38];
  assign o[19918] = i[38];
  assign o[19919] = i[38];
  assign o[19920] = i[38];
  assign o[19921] = i[38];
  assign o[19922] = i[38];
  assign o[19923] = i[38];
  assign o[19924] = i[38];
  assign o[19925] = i[38];
  assign o[19926] = i[38];
  assign o[19927] = i[38];
  assign o[19928] = i[38];
  assign o[19929] = i[38];
  assign o[19930] = i[38];
  assign o[19931] = i[38];
  assign o[19932] = i[38];
  assign o[19933] = i[38];
  assign o[19934] = i[38];
  assign o[19935] = i[38];
  assign o[19936] = i[38];
  assign o[19937] = i[38];
  assign o[19938] = i[38];
  assign o[19939] = i[38];
  assign o[19940] = i[38];
  assign o[19941] = i[38];
  assign o[19942] = i[38];
  assign o[19943] = i[38];
  assign o[19944] = i[38];
  assign o[19945] = i[38];
  assign o[19946] = i[38];
  assign o[19947] = i[38];
  assign o[19948] = i[38];
  assign o[19949] = i[38];
  assign o[19950] = i[38];
  assign o[19951] = i[38];
  assign o[19952] = i[38];
  assign o[19953] = i[38];
  assign o[19954] = i[38];
  assign o[19955] = i[38];
  assign o[19956] = i[38];
  assign o[19957] = i[38];
  assign o[19958] = i[38];
  assign o[19959] = i[38];
  assign o[19960] = i[38];
  assign o[19961] = i[38];
  assign o[19962] = i[38];
  assign o[19963] = i[38];
  assign o[19964] = i[38];
  assign o[19965] = i[38];
  assign o[19966] = i[38];
  assign o[19967] = i[38];
  assign o[18944] = i[37];
  assign o[18945] = i[37];
  assign o[18946] = i[37];
  assign o[18947] = i[37];
  assign o[18948] = i[37];
  assign o[18949] = i[37];
  assign o[18950] = i[37];
  assign o[18951] = i[37];
  assign o[18952] = i[37];
  assign o[18953] = i[37];
  assign o[18954] = i[37];
  assign o[18955] = i[37];
  assign o[18956] = i[37];
  assign o[18957] = i[37];
  assign o[18958] = i[37];
  assign o[18959] = i[37];
  assign o[18960] = i[37];
  assign o[18961] = i[37];
  assign o[18962] = i[37];
  assign o[18963] = i[37];
  assign o[18964] = i[37];
  assign o[18965] = i[37];
  assign o[18966] = i[37];
  assign o[18967] = i[37];
  assign o[18968] = i[37];
  assign o[18969] = i[37];
  assign o[18970] = i[37];
  assign o[18971] = i[37];
  assign o[18972] = i[37];
  assign o[18973] = i[37];
  assign o[18974] = i[37];
  assign o[18975] = i[37];
  assign o[18976] = i[37];
  assign o[18977] = i[37];
  assign o[18978] = i[37];
  assign o[18979] = i[37];
  assign o[18980] = i[37];
  assign o[18981] = i[37];
  assign o[18982] = i[37];
  assign o[18983] = i[37];
  assign o[18984] = i[37];
  assign o[18985] = i[37];
  assign o[18986] = i[37];
  assign o[18987] = i[37];
  assign o[18988] = i[37];
  assign o[18989] = i[37];
  assign o[18990] = i[37];
  assign o[18991] = i[37];
  assign o[18992] = i[37];
  assign o[18993] = i[37];
  assign o[18994] = i[37];
  assign o[18995] = i[37];
  assign o[18996] = i[37];
  assign o[18997] = i[37];
  assign o[18998] = i[37];
  assign o[18999] = i[37];
  assign o[19000] = i[37];
  assign o[19001] = i[37];
  assign o[19002] = i[37];
  assign o[19003] = i[37];
  assign o[19004] = i[37];
  assign o[19005] = i[37];
  assign o[19006] = i[37];
  assign o[19007] = i[37];
  assign o[19008] = i[37];
  assign o[19009] = i[37];
  assign o[19010] = i[37];
  assign o[19011] = i[37];
  assign o[19012] = i[37];
  assign o[19013] = i[37];
  assign o[19014] = i[37];
  assign o[19015] = i[37];
  assign o[19016] = i[37];
  assign o[19017] = i[37];
  assign o[19018] = i[37];
  assign o[19019] = i[37];
  assign o[19020] = i[37];
  assign o[19021] = i[37];
  assign o[19022] = i[37];
  assign o[19023] = i[37];
  assign o[19024] = i[37];
  assign o[19025] = i[37];
  assign o[19026] = i[37];
  assign o[19027] = i[37];
  assign o[19028] = i[37];
  assign o[19029] = i[37];
  assign o[19030] = i[37];
  assign o[19031] = i[37];
  assign o[19032] = i[37];
  assign o[19033] = i[37];
  assign o[19034] = i[37];
  assign o[19035] = i[37];
  assign o[19036] = i[37];
  assign o[19037] = i[37];
  assign o[19038] = i[37];
  assign o[19039] = i[37];
  assign o[19040] = i[37];
  assign o[19041] = i[37];
  assign o[19042] = i[37];
  assign o[19043] = i[37];
  assign o[19044] = i[37];
  assign o[19045] = i[37];
  assign o[19046] = i[37];
  assign o[19047] = i[37];
  assign o[19048] = i[37];
  assign o[19049] = i[37];
  assign o[19050] = i[37];
  assign o[19051] = i[37];
  assign o[19052] = i[37];
  assign o[19053] = i[37];
  assign o[19054] = i[37];
  assign o[19055] = i[37];
  assign o[19056] = i[37];
  assign o[19057] = i[37];
  assign o[19058] = i[37];
  assign o[19059] = i[37];
  assign o[19060] = i[37];
  assign o[19061] = i[37];
  assign o[19062] = i[37];
  assign o[19063] = i[37];
  assign o[19064] = i[37];
  assign o[19065] = i[37];
  assign o[19066] = i[37];
  assign o[19067] = i[37];
  assign o[19068] = i[37];
  assign o[19069] = i[37];
  assign o[19070] = i[37];
  assign o[19071] = i[37];
  assign o[19072] = i[37];
  assign o[19073] = i[37];
  assign o[19074] = i[37];
  assign o[19075] = i[37];
  assign o[19076] = i[37];
  assign o[19077] = i[37];
  assign o[19078] = i[37];
  assign o[19079] = i[37];
  assign o[19080] = i[37];
  assign o[19081] = i[37];
  assign o[19082] = i[37];
  assign o[19083] = i[37];
  assign o[19084] = i[37];
  assign o[19085] = i[37];
  assign o[19086] = i[37];
  assign o[19087] = i[37];
  assign o[19088] = i[37];
  assign o[19089] = i[37];
  assign o[19090] = i[37];
  assign o[19091] = i[37];
  assign o[19092] = i[37];
  assign o[19093] = i[37];
  assign o[19094] = i[37];
  assign o[19095] = i[37];
  assign o[19096] = i[37];
  assign o[19097] = i[37];
  assign o[19098] = i[37];
  assign o[19099] = i[37];
  assign o[19100] = i[37];
  assign o[19101] = i[37];
  assign o[19102] = i[37];
  assign o[19103] = i[37];
  assign o[19104] = i[37];
  assign o[19105] = i[37];
  assign o[19106] = i[37];
  assign o[19107] = i[37];
  assign o[19108] = i[37];
  assign o[19109] = i[37];
  assign o[19110] = i[37];
  assign o[19111] = i[37];
  assign o[19112] = i[37];
  assign o[19113] = i[37];
  assign o[19114] = i[37];
  assign o[19115] = i[37];
  assign o[19116] = i[37];
  assign o[19117] = i[37];
  assign o[19118] = i[37];
  assign o[19119] = i[37];
  assign o[19120] = i[37];
  assign o[19121] = i[37];
  assign o[19122] = i[37];
  assign o[19123] = i[37];
  assign o[19124] = i[37];
  assign o[19125] = i[37];
  assign o[19126] = i[37];
  assign o[19127] = i[37];
  assign o[19128] = i[37];
  assign o[19129] = i[37];
  assign o[19130] = i[37];
  assign o[19131] = i[37];
  assign o[19132] = i[37];
  assign o[19133] = i[37];
  assign o[19134] = i[37];
  assign o[19135] = i[37];
  assign o[19136] = i[37];
  assign o[19137] = i[37];
  assign o[19138] = i[37];
  assign o[19139] = i[37];
  assign o[19140] = i[37];
  assign o[19141] = i[37];
  assign o[19142] = i[37];
  assign o[19143] = i[37];
  assign o[19144] = i[37];
  assign o[19145] = i[37];
  assign o[19146] = i[37];
  assign o[19147] = i[37];
  assign o[19148] = i[37];
  assign o[19149] = i[37];
  assign o[19150] = i[37];
  assign o[19151] = i[37];
  assign o[19152] = i[37];
  assign o[19153] = i[37];
  assign o[19154] = i[37];
  assign o[19155] = i[37];
  assign o[19156] = i[37];
  assign o[19157] = i[37];
  assign o[19158] = i[37];
  assign o[19159] = i[37];
  assign o[19160] = i[37];
  assign o[19161] = i[37];
  assign o[19162] = i[37];
  assign o[19163] = i[37];
  assign o[19164] = i[37];
  assign o[19165] = i[37];
  assign o[19166] = i[37];
  assign o[19167] = i[37];
  assign o[19168] = i[37];
  assign o[19169] = i[37];
  assign o[19170] = i[37];
  assign o[19171] = i[37];
  assign o[19172] = i[37];
  assign o[19173] = i[37];
  assign o[19174] = i[37];
  assign o[19175] = i[37];
  assign o[19176] = i[37];
  assign o[19177] = i[37];
  assign o[19178] = i[37];
  assign o[19179] = i[37];
  assign o[19180] = i[37];
  assign o[19181] = i[37];
  assign o[19182] = i[37];
  assign o[19183] = i[37];
  assign o[19184] = i[37];
  assign o[19185] = i[37];
  assign o[19186] = i[37];
  assign o[19187] = i[37];
  assign o[19188] = i[37];
  assign o[19189] = i[37];
  assign o[19190] = i[37];
  assign o[19191] = i[37];
  assign o[19192] = i[37];
  assign o[19193] = i[37];
  assign o[19194] = i[37];
  assign o[19195] = i[37];
  assign o[19196] = i[37];
  assign o[19197] = i[37];
  assign o[19198] = i[37];
  assign o[19199] = i[37];
  assign o[19200] = i[37];
  assign o[19201] = i[37];
  assign o[19202] = i[37];
  assign o[19203] = i[37];
  assign o[19204] = i[37];
  assign o[19205] = i[37];
  assign o[19206] = i[37];
  assign o[19207] = i[37];
  assign o[19208] = i[37];
  assign o[19209] = i[37];
  assign o[19210] = i[37];
  assign o[19211] = i[37];
  assign o[19212] = i[37];
  assign o[19213] = i[37];
  assign o[19214] = i[37];
  assign o[19215] = i[37];
  assign o[19216] = i[37];
  assign o[19217] = i[37];
  assign o[19218] = i[37];
  assign o[19219] = i[37];
  assign o[19220] = i[37];
  assign o[19221] = i[37];
  assign o[19222] = i[37];
  assign o[19223] = i[37];
  assign o[19224] = i[37];
  assign o[19225] = i[37];
  assign o[19226] = i[37];
  assign o[19227] = i[37];
  assign o[19228] = i[37];
  assign o[19229] = i[37];
  assign o[19230] = i[37];
  assign o[19231] = i[37];
  assign o[19232] = i[37];
  assign o[19233] = i[37];
  assign o[19234] = i[37];
  assign o[19235] = i[37];
  assign o[19236] = i[37];
  assign o[19237] = i[37];
  assign o[19238] = i[37];
  assign o[19239] = i[37];
  assign o[19240] = i[37];
  assign o[19241] = i[37];
  assign o[19242] = i[37];
  assign o[19243] = i[37];
  assign o[19244] = i[37];
  assign o[19245] = i[37];
  assign o[19246] = i[37];
  assign o[19247] = i[37];
  assign o[19248] = i[37];
  assign o[19249] = i[37];
  assign o[19250] = i[37];
  assign o[19251] = i[37];
  assign o[19252] = i[37];
  assign o[19253] = i[37];
  assign o[19254] = i[37];
  assign o[19255] = i[37];
  assign o[19256] = i[37];
  assign o[19257] = i[37];
  assign o[19258] = i[37];
  assign o[19259] = i[37];
  assign o[19260] = i[37];
  assign o[19261] = i[37];
  assign o[19262] = i[37];
  assign o[19263] = i[37];
  assign o[19264] = i[37];
  assign o[19265] = i[37];
  assign o[19266] = i[37];
  assign o[19267] = i[37];
  assign o[19268] = i[37];
  assign o[19269] = i[37];
  assign o[19270] = i[37];
  assign o[19271] = i[37];
  assign o[19272] = i[37];
  assign o[19273] = i[37];
  assign o[19274] = i[37];
  assign o[19275] = i[37];
  assign o[19276] = i[37];
  assign o[19277] = i[37];
  assign o[19278] = i[37];
  assign o[19279] = i[37];
  assign o[19280] = i[37];
  assign o[19281] = i[37];
  assign o[19282] = i[37];
  assign o[19283] = i[37];
  assign o[19284] = i[37];
  assign o[19285] = i[37];
  assign o[19286] = i[37];
  assign o[19287] = i[37];
  assign o[19288] = i[37];
  assign o[19289] = i[37];
  assign o[19290] = i[37];
  assign o[19291] = i[37];
  assign o[19292] = i[37];
  assign o[19293] = i[37];
  assign o[19294] = i[37];
  assign o[19295] = i[37];
  assign o[19296] = i[37];
  assign o[19297] = i[37];
  assign o[19298] = i[37];
  assign o[19299] = i[37];
  assign o[19300] = i[37];
  assign o[19301] = i[37];
  assign o[19302] = i[37];
  assign o[19303] = i[37];
  assign o[19304] = i[37];
  assign o[19305] = i[37];
  assign o[19306] = i[37];
  assign o[19307] = i[37];
  assign o[19308] = i[37];
  assign o[19309] = i[37];
  assign o[19310] = i[37];
  assign o[19311] = i[37];
  assign o[19312] = i[37];
  assign o[19313] = i[37];
  assign o[19314] = i[37];
  assign o[19315] = i[37];
  assign o[19316] = i[37];
  assign o[19317] = i[37];
  assign o[19318] = i[37];
  assign o[19319] = i[37];
  assign o[19320] = i[37];
  assign o[19321] = i[37];
  assign o[19322] = i[37];
  assign o[19323] = i[37];
  assign o[19324] = i[37];
  assign o[19325] = i[37];
  assign o[19326] = i[37];
  assign o[19327] = i[37];
  assign o[19328] = i[37];
  assign o[19329] = i[37];
  assign o[19330] = i[37];
  assign o[19331] = i[37];
  assign o[19332] = i[37];
  assign o[19333] = i[37];
  assign o[19334] = i[37];
  assign o[19335] = i[37];
  assign o[19336] = i[37];
  assign o[19337] = i[37];
  assign o[19338] = i[37];
  assign o[19339] = i[37];
  assign o[19340] = i[37];
  assign o[19341] = i[37];
  assign o[19342] = i[37];
  assign o[19343] = i[37];
  assign o[19344] = i[37];
  assign o[19345] = i[37];
  assign o[19346] = i[37];
  assign o[19347] = i[37];
  assign o[19348] = i[37];
  assign o[19349] = i[37];
  assign o[19350] = i[37];
  assign o[19351] = i[37];
  assign o[19352] = i[37];
  assign o[19353] = i[37];
  assign o[19354] = i[37];
  assign o[19355] = i[37];
  assign o[19356] = i[37];
  assign o[19357] = i[37];
  assign o[19358] = i[37];
  assign o[19359] = i[37];
  assign o[19360] = i[37];
  assign o[19361] = i[37];
  assign o[19362] = i[37];
  assign o[19363] = i[37];
  assign o[19364] = i[37];
  assign o[19365] = i[37];
  assign o[19366] = i[37];
  assign o[19367] = i[37];
  assign o[19368] = i[37];
  assign o[19369] = i[37];
  assign o[19370] = i[37];
  assign o[19371] = i[37];
  assign o[19372] = i[37];
  assign o[19373] = i[37];
  assign o[19374] = i[37];
  assign o[19375] = i[37];
  assign o[19376] = i[37];
  assign o[19377] = i[37];
  assign o[19378] = i[37];
  assign o[19379] = i[37];
  assign o[19380] = i[37];
  assign o[19381] = i[37];
  assign o[19382] = i[37];
  assign o[19383] = i[37];
  assign o[19384] = i[37];
  assign o[19385] = i[37];
  assign o[19386] = i[37];
  assign o[19387] = i[37];
  assign o[19388] = i[37];
  assign o[19389] = i[37];
  assign o[19390] = i[37];
  assign o[19391] = i[37];
  assign o[19392] = i[37];
  assign o[19393] = i[37];
  assign o[19394] = i[37];
  assign o[19395] = i[37];
  assign o[19396] = i[37];
  assign o[19397] = i[37];
  assign o[19398] = i[37];
  assign o[19399] = i[37];
  assign o[19400] = i[37];
  assign o[19401] = i[37];
  assign o[19402] = i[37];
  assign o[19403] = i[37];
  assign o[19404] = i[37];
  assign o[19405] = i[37];
  assign o[19406] = i[37];
  assign o[19407] = i[37];
  assign o[19408] = i[37];
  assign o[19409] = i[37];
  assign o[19410] = i[37];
  assign o[19411] = i[37];
  assign o[19412] = i[37];
  assign o[19413] = i[37];
  assign o[19414] = i[37];
  assign o[19415] = i[37];
  assign o[19416] = i[37];
  assign o[19417] = i[37];
  assign o[19418] = i[37];
  assign o[19419] = i[37];
  assign o[19420] = i[37];
  assign o[19421] = i[37];
  assign o[19422] = i[37];
  assign o[19423] = i[37];
  assign o[19424] = i[37];
  assign o[19425] = i[37];
  assign o[19426] = i[37];
  assign o[19427] = i[37];
  assign o[19428] = i[37];
  assign o[19429] = i[37];
  assign o[19430] = i[37];
  assign o[19431] = i[37];
  assign o[19432] = i[37];
  assign o[19433] = i[37];
  assign o[19434] = i[37];
  assign o[19435] = i[37];
  assign o[19436] = i[37];
  assign o[19437] = i[37];
  assign o[19438] = i[37];
  assign o[19439] = i[37];
  assign o[19440] = i[37];
  assign o[19441] = i[37];
  assign o[19442] = i[37];
  assign o[19443] = i[37];
  assign o[19444] = i[37];
  assign o[19445] = i[37];
  assign o[19446] = i[37];
  assign o[19447] = i[37];
  assign o[19448] = i[37];
  assign o[19449] = i[37];
  assign o[19450] = i[37];
  assign o[19451] = i[37];
  assign o[19452] = i[37];
  assign o[19453] = i[37];
  assign o[19454] = i[37];
  assign o[19455] = i[37];
  assign o[18432] = i[36];
  assign o[18433] = i[36];
  assign o[18434] = i[36];
  assign o[18435] = i[36];
  assign o[18436] = i[36];
  assign o[18437] = i[36];
  assign o[18438] = i[36];
  assign o[18439] = i[36];
  assign o[18440] = i[36];
  assign o[18441] = i[36];
  assign o[18442] = i[36];
  assign o[18443] = i[36];
  assign o[18444] = i[36];
  assign o[18445] = i[36];
  assign o[18446] = i[36];
  assign o[18447] = i[36];
  assign o[18448] = i[36];
  assign o[18449] = i[36];
  assign o[18450] = i[36];
  assign o[18451] = i[36];
  assign o[18452] = i[36];
  assign o[18453] = i[36];
  assign o[18454] = i[36];
  assign o[18455] = i[36];
  assign o[18456] = i[36];
  assign o[18457] = i[36];
  assign o[18458] = i[36];
  assign o[18459] = i[36];
  assign o[18460] = i[36];
  assign o[18461] = i[36];
  assign o[18462] = i[36];
  assign o[18463] = i[36];
  assign o[18464] = i[36];
  assign o[18465] = i[36];
  assign o[18466] = i[36];
  assign o[18467] = i[36];
  assign o[18468] = i[36];
  assign o[18469] = i[36];
  assign o[18470] = i[36];
  assign o[18471] = i[36];
  assign o[18472] = i[36];
  assign o[18473] = i[36];
  assign o[18474] = i[36];
  assign o[18475] = i[36];
  assign o[18476] = i[36];
  assign o[18477] = i[36];
  assign o[18478] = i[36];
  assign o[18479] = i[36];
  assign o[18480] = i[36];
  assign o[18481] = i[36];
  assign o[18482] = i[36];
  assign o[18483] = i[36];
  assign o[18484] = i[36];
  assign o[18485] = i[36];
  assign o[18486] = i[36];
  assign o[18487] = i[36];
  assign o[18488] = i[36];
  assign o[18489] = i[36];
  assign o[18490] = i[36];
  assign o[18491] = i[36];
  assign o[18492] = i[36];
  assign o[18493] = i[36];
  assign o[18494] = i[36];
  assign o[18495] = i[36];
  assign o[18496] = i[36];
  assign o[18497] = i[36];
  assign o[18498] = i[36];
  assign o[18499] = i[36];
  assign o[18500] = i[36];
  assign o[18501] = i[36];
  assign o[18502] = i[36];
  assign o[18503] = i[36];
  assign o[18504] = i[36];
  assign o[18505] = i[36];
  assign o[18506] = i[36];
  assign o[18507] = i[36];
  assign o[18508] = i[36];
  assign o[18509] = i[36];
  assign o[18510] = i[36];
  assign o[18511] = i[36];
  assign o[18512] = i[36];
  assign o[18513] = i[36];
  assign o[18514] = i[36];
  assign o[18515] = i[36];
  assign o[18516] = i[36];
  assign o[18517] = i[36];
  assign o[18518] = i[36];
  assign o[18519] = i[36];
  assign o[18520] = i[36];
  assign o[18521] = i[36];
  assign o[18522] = i[36];
  assign o[18523] = i[36];
  assign o[18524] = i[36];
  assign o[18525] = i[36];
  assign o[18526] = i[36];
  assign o[18527] = i[36];
  assign o[18528] = i[36];
  assign o[18529] = i[36];
  assign o[18530] = i[36];
  assign o[18531] = i[36];
  assign o[18532] = i[36];
  assign o[18533] = i[36];
  assign o[18534] = i[36];
  assign o[18535] = i[36];
  assign o[18536] = i[36];
  assign o[18537] = i[36];
  assign o[18538] = i[36];
  assign o[18539] = i[36];
  assign o[18540] = i[36];
  assign o[18541] = i[36];
  assign o[18542] = i[36];
  assign o[18543] = i[36];
  assign o[18544] = i[36];
  assign o[18545] = i[36];
  assign o[18546] = i[36];
  assign o[18547] = i[36];
  assign o[18548] = i[36];
  assign o[18549] = i[36];
  assign o[18550] = i[36];
  assign o[18551] = i[36];
  assign o[18552] = i[36];
  assign o[18553] = i[36];
  assign o[18554] = i[36];
  assign o[18555] = i[36];
  assign o[18556] = i[36];
  assign o[18557] = i[36];
  assign o[18558] = i[36];
  assign o[18559] = i[36];
  assign o[18560] = i[36];
  assign o[18561] = i[36];
  assign o[18562] = i[36];
  assign o[18563] = i[36];
  assign o[18564] = i[36];
  assign o[18565] = i[36];
  assign o[18566] = i[36];
  assign o[18567] = i[36];
  assign o[18568] = i[36];
  assign o[18569] = i[36];
  assign o[18570] = i[36];
  assign o[18571] = i[36];
  assign o[18572] = i[36];
  assign o[18573] = i[36];
  assign o[18574] = i[36];
  assign o[18575] = i[36];
  assign o[18576] = i[36];
  assign o[18577] = i[36];
  assign o[18578] = i[36];
  assign o[18579] = i[36];
  assign o[18580] = i[36];
  assign o[18581] = i[36];
  assign o[18582] = i[36];
  assign o[18583] = i[36];
  assign o[18584] = i[36];
  assign o[18585] = i[36];
  assign o[18586] = i[36];
  assign o[18587] = i[36];
  assign o[18588] = i[36];
  assign o[18589] = i[36];
  assign o[18590] = i[36];
  assign o[18591] = i[36];
  assign o[18592] = i[36];
  assign o[18593] = i[36];
  assign o[18594] = i[36];
  assign o[18595] = i[36];
  assign o[18596] = i[36];
  assign o[18597] = i[36];
  assign o[18598] = i[36];
  assign o[18599] = i[36];
  assign o[18600] = i[36];
  assign o[18601] = i[36];
  assign o[18602] = i[36];
  assign o[18603] = i[36];
  assign o[18604] = i[36];
  assign o[18605] = i[36];
  assign o[18606] = i[36];
  assign o[18607] = i[36];
  assign o[18608] = i[36];
  assign o[18609] = i[36];
  assign o[18610] = i[36];
  assign o[18611] = i[36];
  assign o[18612] = i[36];
  assign o[18613] = i[36];
  assign o[18614] = i[36];
  assign o[18615] = i[36];
  assign o[18616] = i[36];
  assign o[18617] = i[36];
  assign o[18618] = i[36];
  assign o[18619] = i[36];
  assign o[18620] = i[36];
  assign o[18621] = i[36];
  assign o[18622] = i[36];
  assign o[18623] = i[36];
  assign o[18624] = i[36];
  assign o[18625] = i[36];
  assign o[18626] = i[36];
  assign o[18627] = i[36];
  assign o[18628] = i[36];
  assign o[18629] = i[36];
  assign o[18630] = i[36];
  assign o[18631] = i[36];
  assign o[18632] = i[36];
  assign o[18633] = i[36];
  assign o[18634] = i[36];
  assign o[18635] = i[36];
  assign o[18636] = i[36];
  assign o[18637] = i[36];
  assign o[18638] = i[36];
  assign o[18639] = i[36];
  assign o[18640] = i[36];
  assign o[18641] = i[36];
  assign o[18642] = i[36];
  assign o[18643] = i[36];
  assign o[18644] = i[36];
  assign o[18645] = i[36];
  assign o[18646] = i[36];
  assign o[18647] = i[36];
  assign o[18648] = i[36];
  assign o[18649] = i[36];
  assign o[18650] = i[36];
  assign o[18651] = i[36];
  assign o[18652] = i[36];
  assign o[18653] = i[36];
  assign o[18654] = i[36];
  assign o[18655] = i[36];
  assign o[18656] = i[36];
  assign o[18657] = i[36];
  assign o[18658] = i[36];
  assign o[18659] = i[36];
  assign o[18660] = i[36];
  assign o[18661] = i[36];
  assign o[18662] = i[36];
  assign o[18663] = i[36];
  assign o[18664] = i[36];
  assign o[18665] = i[36];
  assign o[18666] = i[36];
  assign o[18667] = i[36];
  assign o[18668] = i[36];
  assign o[18669] = i[36];
  assign o[18670] = i[36];
  assign o[18671] = i[36];
  assign o[18672] = i[36];
  assign o[18673] = i[36];
  assign o[18674] = i[36];
  assign o[18675] = i[36];
  assign o[18676] = i[36];
  assign o[18677] = i[36];
  assign o[18678] = i[36];
  assign o[18679] = i[36];
  assign o[18680] = i[36];
  assign o[18681] = i[36];
  assign o[18682] = i[36];
  assign o[18683] = i[36];
  assign o[18684] = i[36];
  assign o[18685] = i[36];
  assign o[18686] = i[36];
  assign o[18687] = i[36];
  assign o[18688] = i[36];
  assign o[18689] = i[36];
  assign o[18690] = i[36];
  assign o[18691] = i[36];
  assign o[18692] = i[36];
  assign o[18693] = i[36];
  assign o[18694] = i[36];
  assign o[18695] = i[36];
  assign o[18696] = i[36];
  assign o[18697] = i[36];
  assign o[18698] = i[36];
  assign o[18699] = i[36];
  assign o[18700] = i[36];
  assign o[18701] = i[36];
  assign o[18702] = i[36];
  assign o[18703] = i[36];
  assign o[18704] = i[36];
  assign o[18705] = i[36];
  assign o[18706] = i[36];
  assign o[18707] = i[36];
  assign o[18708] = i[36];
  assign o[18709] = i[36];
  assign o[18710] = i[36];
  assign o[18711] = i[36];
  assign o[18712] = i[36];
  assign o[18713] = i[36];
  assign o[18714] = i[36];
  assign o[18715] = i[36];
  assign o[18716] = i[36];
  assign o[18717] = i[36];
  assign o[18718] = i[36];
  assign o[18719] = i[36];
  assign o[18720] = i[36];
  assign o[18721] = i[36];
  assign o[18722] = i[36];
  assign o[18723] = i[36];
  assign o[18724] = i[36];
  assign o[18725] = i[36];
  assign o[18726] = i[36];
  assign o[18727] = i[36];
  assign o[18728] = i[36];
  assign o[18729] = i[36];
  assign o[18730] = i[36];
  assign o[18731] = i[36];
  assign o[18732] = i[36];
  assign o[18733] = i[36];
  assign o[18734] = i[36];
  assign o[18735] = i[36];
  assign o[18736] = i[36];
  assign o[18737] = i[36];
  assign o[18738] = i[36];
  assign o[18739] = i[36];
  assign o[18740] = i[36];
  assign o[18741] = i[36];
  assign o[18742] = i[36];
  assign o[18743] = i[36];
  assign o[18744] = i[36];
  assign o[18745] = i[36];
  assign o[18746] = i[36];
  assign o[18747] = i[36];
  assign o[18748] = i[36];
  assign o[18749] = i[36];
  assign o[18750] = i[36];
  assign o[18751] = i[36];
  assign o[18752] = i[36];
  assign o[18753] = i[36];
  assign o[18754] = i[36];
  assign o[18755] = i[36];
  assign o[18756] = i[36];
  assign o[18757] = i[36];
  assign o[18758] = i[36];
  assign o[18759] = i[36];
  assign o[18760] = i[36];
  assign o[18761] = i[36];
  assign o[18762] = i[36];
  assign o[18763] = i[36];
  assign o[18764] = i[36];
  assign o[18765] = i[36];
  assign o[18766] = i[36];
  assign o[18767] = i[36];
  assign o[18768] = i[36];
  assign o[18769] = i[36];
  assign o[18770] = i[36];
  assign o[18771] = i[36];
  assign o[18772] = i[36];
  assign o[18773] = i[36];
  assign o[18774] = i[36];
  assign o[18775] = i[36];
  assign o[18776] = i[36];
  assign o[18777] = i[36];
  assign o[18778] = i[36];
  assign o[18779] = i[36];
  assign o[18780] = i[36];
  assign o[18781] = i[36];
  assign o[18782] = i[36];
  assign o[18783] = i[36];
  assign o[18784] = i[36];
  assign o[18785] = i[36];
  assign o[18786] = i[36];
  assign o[18787] = i[36];
  assign o[18788] = i[36];
  assign o[18789] = i[36];
  assign o[18790] = i[36];
  assign o[18791] = i[36];
  assign o[18792] = i[36];
  assign o[18793] = i[36];
  assign o[18794] = i[36];
  assign o[18795] = i[36];
  assign o[18796] = i[36];
  assign o[18797] = i[36];
  assign o[18798] = i[36];
  assign o[18799] = i[36];
  assign o[18800] = i[36];
  assign o[18801] = i[36];
  assign o[18802] = i[36];
  assign o[18803] = i[36];
  assign o[18804] = i[36];
  assign o[18805] = i[36];
  assign o[18806] = i[36];
  assign o[18807] = i[36];
  assign o[18808] = i[36];
  assign o[18809] = i[36];
  assign o[18810] = i[36];
  assign o[18811] = i[36];
  assign o[18812] = i[36];
  assign o[18813] = i[36];
  assign o[18814] = i[36];
  assign o[18815] = i[36];
  assign o[18816] = i[36];
  assign o[18817] = i[36];
  assign o[18818] = i[36];
  assign o[18819] = i[36];
  assign o[18820] = i[36];
  assign o[18821] = i[36];
  assign o[18822] = i[36];
  assign o[18823] = i[36];
  assign o[18824] = i[36];
  assign o[18825] = i[36];
  assign o[18826] = i[36];
  assign o[18827] = i[36];
  assign o[18828] = i[36];
  assign o[18829] = i[36];
  assign o[18830] = i[36];
  assign o[18831] = i[36];
  assign o[18832] = i[36];
  assign o[18833] = i[36];
  assign o[18834] = i[36];
  assign o[18835] = i[36];
  assign o[18836] = i[36];
  assign o[18837] = i[36];
  assign o[18838] = i[36];
  assign o[18839] = i[36];
  assign o[18840] = i[36];
  assign o[18841] = i[36];
  assign o[18842] = i[36];
  assign o[18843] = i[36];
  assign o[18844] = i[36];
  assign o[18845] = i[36];
  assign o[18846] = i[36];
  assign o[18847] = i[36];
  assign o[18848] = i[36];
  assign o[18849] = i[36];
  assign o[18850] = i[36];
  assign o[18851] = i[36];
  assign o[18852] = i[36];
  assign o[18853] = i[36];
  assign o[18854] = i[36];
  assign o[18855] = i[36];
  assign o[18856] = i[36];
  assign o[18857] = i[36];
  assign o[18858] = i[36];
  assign o[18859] = i[36];
  assign o[18860] = i[36];
  assign o[18861] = i[36];
  assign o[18862] = i[36];
  assign o[18863] = i[36];
  assign o[18864] = i[36];
  assign o[18865] = i[36];
  assign o[18866] = i[36];
  assign o[18867] = i[36];
  assign o[18868] = i[36];
  assign o[18869] = i[36];
  assign o[18870] = i[36];
  assign o[18871] = i[36];
  assign o[18872] = i[36];
  assign o[18873] = i[36];
  assign o[18874] = i[36];
  assign o[18875] = i[36];
  assign o[18876] = i[36];
  assign o[18877] = i[36];
  assign o[18878] = i[36];
  assign o[18879] = i[36];
  assign o[18880] = i[36];
  assign o[18881] = i[36];
  assign o[18882] = i[36];
  assign o[18883] = i[36];
  assign o[18884] = i[36];
  assign o[18885] = i[36];
  assign o[18886] = i[36];
  assign o[18887] = i[36];
  assign o[18888] = i[36];
  assign o[18889] = i[36];
  assign o[18890] = i[36];
  assign o[18891] = i[36];
  assign o[18892] = i[36];
  assign o[18893] = i[36];
  assign o[18894] = i[36];
  assign o[18895] = i[36];
  assign o[18896] = i[36];
  assign o[18897] = i[36];
  assign o[18898] = i[36];
  assign o[18899] = i[36];
  assign o[18900] = i[36];
  assign o[18901] = i[36];
  assign o[18902] = i[36];
  assign o[18903] = i[36];
  assign o[18904] = i[36];
  assign o[18905] = i[36];
  assign o[18906] = i[36];
  assign o[18907] = i[36];
  assign o[18908] = i[36];
  assign o[18909] = i[36];
  assign o[18910] = i[36];
  assign o[18911] = i[36];
  assign o[18912] = i[36];
  assign o[18913] = i[36];
  assign o[18914] = i[36];
  assign o[18915] = i[36];
  assign o[18916] = i[36];
  assign o[18917] = i[36];
  assign o[18918] = i[36];
  assign o[18919] = i[36];
  assign o[18920] = i[36];
  assign o[18921] = i[36];
  assign o[18922] = i[36];
  assign o[18923] = i[36];
  assign o[18924] = i[36];
  assign o[18925] = i[36];
  assign o[18926] = i[36];
  assign o[18927] = i[36];
  assign o[18928] = i[36];
  assign o[18929] = i[36];
  assign o[18930] = i[36];
  assign o[18931] = i[36];
  assign o[18932] = i[36];
  assign o[18933] = i[36];
  assign o[18934] = i[36];
  assign o[18935] = i[36];
  assign o[18936] = i[36];
  assign o[18937] = i[36];
  assign o[18938] = i[36];
  assign o[18939] = i[36];
  assign o[18940] = i[36];
  assign o[18941] = i[36];
  assign o[18942] = i[36];
  assign o[18943] = i[36];
  assign o[17920] = i[35];
  assign o[17921] = i[35];
  assign o[17922] = i[35];
  assign o[17923] = i[35];
  assign o[17924] = i[35];
  assign o[17925] = i[35];
  assign o[17926] = i[35];
  assign o[17927] = i[35];
  assign o[17928] = i[35];
  assign o[17929] = i[35];
  assign o[17930] = i[35];
  assign o[17931] = i[35];
  assign o[17932] = i[35];
  assign o[17933] = i[35];
  assign o[17934] = i[35];
  assign o[17935] = i[35];
  assign o[17936] = i[35];
  assign o[17937] = i[35];
  assign o[17938] = i[35];
  assign o[17939] = i[35];
  assign o[17940] = i[35];
  assign o[17941] = i[35];
  assign o[17942] = i[35];
  assign o[17943] = i[35];
  assign o[17944] = i[35];
  assign o[17945] = i[35];
  assign o[17946] = i[35];
  assign o[17947] = i[35];
  assign o[17948] = i[35];
  assign o[17949] = i[35];
  assign o[17950] = i[35];
  assign o[17951] = i[35];
  assign o[17952] = i[35];
  assign o[17953] = i[35];
  assign o[17954] = i[35];
  assign o[17955] = i[35];
  assign o[17956] = i[35];
  assign o[17957] = i[35];
  assign o[17958] = i[35];
  assign o[17959] = i[35];
  assign o[17960] = i[35];
  assign o[17961] = i[35];
  assign o[17962] = i[35];
  assign o[17963] = i[35];
  assign o[17964] = i[35];
  assign o[17965] = i[35];
  assign o[17966] = i[35];
  assign o[17967] = i[35];
  assign o[17968] = i[35];
  assign o[17969] = i[35];
  assign o[17970] = i[35];
  assign o[17971] = i[35];
  assign o[17972] = i[35];
  assign o[17973] = i[35];
  assign o[17974] = i[35];
  assign o[17975] = i[35];
  assign o[17976] = i[35];
  assign o[17977] = i[35];
  assign o[17978] = i[35];
  assign o[17979] = i[35];
  assign o[17980] = i[35];
  assign o[17981] = i[35];
  assign o[17982] = i[35];
  assign o[17983] = i[35];
  assign o[17984] = i[35];
  assign o[17985] = i[35];
  assign o[17986] = i[35];
  assign o[17987] = i[35];
  assign o[17988] = i[35];
  assign o[17989] = i[35];
  assign o[17990] = i[35];
  assign o[17991] = i[35];
  assign o[17992] = i[35];
  assign o[17993] = i[35];
  assign o[17994] = i[35];
  assign o[17995] = i[35];
  assign o[17996] = i[35];
  assign o[17997] = i[35];
  assign o[17998] = i[35];
  assign o[17999] = i[35];
  assign o[18000] = i[35];
  assign o[18001] = i[35];
  assign o[18002] = i[35];
  assign o[18003] = i[35];
  assign o[18004] = i[35];
  assign o[18005] = i[35];
  assign o[18006] = i[35];
  assign o[18007] = i[35];
  assign o[18008] = i[35];
  assign o[18009] = i[35];
  assign o[18010] = i[35];
  assign o[18011] = i[35];
  assign o[18012] = i[35];
  assign o[18013] = i[35];
  assign o[18014] = i[35];
  assign o[18015] = i[35];
  assign o[18016] = i[35];
  assign o[18017] = i[35];
  assign o[18018] = i[35];
  assign o[18019] = i[35];
  assign o[18020] = i[35];
  assign o[18021] = i[35];
  assign o[18022] = i[35];
  assign o[18023] = i[35];
  assign o[18024] = i[35];
  assign o[18025] = i[35];
  assign o[18026] = i[35];
  assign o[18027] = i[35];
  assign o[18028] = i[35];
  assign o[18029] = i[35];
  assign o[18030] = i[35];
  assign o[18031] = i[35];
  assign o[18032] = i[35];
  assign o[18033] = i[35];
  assign o[18034] = i[35];
  assign o[18035] = i[35];
  assign o[18036] = i[35];
  assign o[18037] = i[35];
  assign o[18038] = i[35];
  assign o[18039] = i[35];
  assign o[18040] = i[35];
  assign o[18041] = i[35];
  assign o[18042] = i[35];
  assign o[18043] = i[35];
  assign o[18044] = i[35];
  assign o[18045] = i[35];
  assign o[18046] = i[35];
  assign o[18047] = i[35];
  assign o[18048] = i[35];
  assign o[18049] = i[35];
  assign o[18050] = i[35];
  assign o[18051] = i[35];
  assign o[18052] = i[35];
  assign o[18053] = i[35];
  assign o[18054] = i[35];
  assign o[18055] = i[35];
  assign o[18056] = i[35];
  assign o[18057] = i[35];
  assign o[18058] = i[35];
  assign o[18059] = i[35];
  assign o[18060] = i[35];
  assign o[18061] = i[35];
  assign o[18062] = i[35];
  assign o[18063] = i[35];
  assign o[18064] = i[35];
  assign o[18065] = i[35];
  assign o[18066] = i[35];
  assign o[18067] = i[35];
  assign o[18068] = i[35];
  assign o[18069] = i[35];
  assign o[18070] = i[35];
  assign o[18071] = i[35];
  assign o[18072] = i[35];
  assign o[18073] = i[35];
  assign o[18074] = i[35];
  assign o[18075] = i[35];
  assign o[18076] = i[35];
  assign o[18077] = i[35];
  assign o[18078] = i[35];
  assign o[18079] = i[35];
  assign o[18080] = i[35];
  assign o[18081] = i[35];
  assign o[18082] = i[35];
  assign o[18083] = i[35];
  assign o[18084] = i[35];
  assign o[18085] = i[35];
  assign o[18086] = i[35];
  assign o[18087] = i[35];
  assign o[18088] = i[35];
  assign o[18089] = i[35];
  assign o[18090] = i[35];
  assign o[18091] = i[35];
  assign o[18092] = i[35];
  assign o[18093] = i[35];
  assign o[18094] = i[35];
  assign o[18095] = i[35];
  assign o[18096] = i[35];
  assign o[18097] = i[35];
  assign o[18098] = i[35];
  assign o[18099] = i[35];
  assign o[18100] = i[35];
  assign o[18101] = i[35];
  assign o[18102] = i[35];
  assign o[18103] = i[35];
  assign o[18104] = i[35];
  assign o[18105] = i[35];
  assign o[18106] = i[35];
  assign o[18107] = i[35];
  assign o[18108] = i[35];
  assign o[18109] = i[35];
  assign o[18110] = i[35];
  assign o[18111] = i[35];
  assign o[18112] = i[35];
  assign o[18113] = i[35];
  assign o[18114] = i[35];
  assign o[18115] = i[35];
  assign o[18116] = i[35];
  assign o[18117] = i[35];
  assign o[18118] = i[35];
  assign o[18119] = i[35];
  assign o[18120] = i[35];
  assign o[18121] = i[35];
  assign o[18122] = i[35];
  assign o[18123] = i[35];
  assign o[18124] = i[35];
  assign o[18125] = i[35];
  assign o[18126] = i[35];
  assign o[18127] = i[35];
  assign o[18128] = i[35];
  assign o[18129] = i[35];
  assign o[18130] = i[35];
  assign o[18131] = i[35];
  assign o[18132] = i[35];
  assign o[18133] = i[35];
  assign o[18134] = i[35];
  assign o[18135] = i[35];
  assign o[18136] = i[35];
  assign o[18137] = i[35];
  assign o[18138] = i[35];
  assign o[18139] = i[35];
  assign o[18140] = i[35];
  assign o[18141] = i[35];
  assign o[18142] = i[35];
  assign o[18143] = i[35];
  assign o[18144] = i[35];
  assign o[18145] = i[35];
  assign o[18146] = i[35];
  assign o[18147] = i[35];
  assign o[18148] = i[35];
  assign o[18149] = i[35];
  assign o[18150] = i[35];
  assign o[18151] = i[35];
  assign o[18152] = i[35];
  assign o[18153] = i[35];
  assign o[18154] = i[35];
  assign o[18155] = i[35];
  assign o[18156] = i[35];
  assign o[18157] = i[35];
  assign o[18158] = i[35];
  assign o[18159] = i[35];
  assign o[18160] = i[35];
  assign o[18161] = i[35];
  assign o[18162] = i[35];
  assign o[18163] = i[35];
  assign o[18164] = i[35];
  assign o[18165] = i[35];
  assign o[18166] = i[35];
  assign o[18167] = i[35];
  assign o[18168] = i[35];
  assign o[18169] = i[35];
  assign o[18170] = i[35];
  assign o[18171] = i[35];
  assign o[18172] = i[35];
  assign o[18173] = i[35];
  assign o[18174] = i[35];
  assign o[18175] = i[35];
  assign o[18176] = i[35];
  assign o[18177] = i[35];
  assign o[18178] = i[35];
  assign o[18179] = i[35];
  assign o[18180] = i[35];
  assign o[18181] = i[35];
  assign o[18182] = i[35];
  assign o[18183] = i[35];
  assign o[18184] = i[35];
  assign o[18185] = i[35];
  assign o[18186] = i[35];
  assign o[18187] = i[35];
  assign o[18188] = i[35];
  assign o[18189] = i[35];
  assign o[18190] = i[35];
  assign o[18191] = i[35];
  assign o[18192] = i[35];
  assign o[18193] = i[35];
  assign o[18194] = i[35];
  assign o[18195] = i[35];
  assign o[18196] = i[35];
  assign o[18197] = i[35];
  assign o[18198] = i[35];
  assign o[18199] = i[35];
  assign o[18200] = i[35];
  assign o[18201] = i[35];
  assign o[18202] = i[35];
  assign o[18203] = i[35];
  assign o[18204] = i[35];
  assign o[18205] = i[35];
  assign o[18206] = i[35];
  assign o[18207] = i[35];
  assign o[18208] = i[35];
  assign o[18209] = i[35];
  assign o[18210] = i[35];
  assign o[18211] = i[35];
  assign o[18212] = i[35];
  assign o[18213] = i[35];
  assign o[18214] = i[35];
  assign o[18215] = i[35];
  assign o[18216] = i[35];
  assign o[18217] = i[35];
  assign o[18218] = i[35];
  assign o[18219] = i[35];
  assign o[18220] = i[35];
  assign o[18221] = i[35];
  assign o[18222] = i[35];
  assign o[18223] = i[35];
  assign o[18224] = i[35];
  assign o[18225] = i[35];
  assign o[18226] = i[35];
  assign o[18227] = i[35];
  assign o[18228] = i[35];
  assign o[18229] = i[35];
  assign o[18230] = i[35];
  assign o[18231] = i[35];
  assign o[18232] = i[35];
  assign o[18233] = i[35];
  assign o[18234] = i[35];
  assign o[18235] = i[35];
  assign o[18236] = i[35];
  assign o[18237] = i[35];
  assign o[18238] = i[35];
  assign o[18239] = i[35];
  assign o[18240] = i[35];
  assign o[18241] = i[35];
  assign o[18242] = i[35];
  assign o[18243] = i[35];
  assign o[18244] = i[35];
  assign o[18245] = i[35];
  assign o[18246] = i[35];
  assign o[18247] = i[35];
  assign o[18248] = i[35];
  assign o[18249] = i[35];
  assign o[18250] = i[35];
  assign o[18251] = i[35];
  assign o[18252] = i[35];
  assign o[18253] = i[35];
  assign o[18254] = i[35];
  assign o[18255] = i[35];
  assign o[18256] = i[35];
  assign o[18257] = i[35];
  assign o[18258] = i[35];
  assign o[18259] = i[35];
  assign o[18260] = i[35];
  assign o[18261] = i[35];
  assign o[18262] = i[35];
  assign o[18263] = i[35];
  assign o[18264] = i[35];
  assign o[18265] = i[35];
  assign o[18266] = i[35];
  assign o[18267] = i[35];
  assign o[18268] = i[35];
  assign o[18269] = i[35];
  assign o[18270] = i[35];
  assign o[18271] = i[35];
  assign o[18272] = i[35];
  assign o[18273] = i[35];
  assign o[18274] = i[35];
  assign o[18275] = i[35];
  assign o[18276] = i[35];
  assign o[18277] = i[35];
  assign o[18278] = i[35];
  assign o[18279] = i[35];
  assign o[18280] = i[35];
  assign o[18281] = i[35];
  assign o[18282] = i[35];
  assign o[18283] = i[35];
  assign o[18284] = i[35];
  assign o[18285] = i[35];
  assign o[18286] = i[35];
  assign o[18287] = i[35];
  assign o[18288] = i[35];
  assign o[18289] = i[35];
  assign o[18290] = i[35];
  assign o[18291] = i[35];
  assign o[18292] = i[35];
  assign o[18293] = i[35];
  assign o[18294] = i[35];
  assign o[18295] = i[35];
  assign o[18296] = i[35];
  assign o[18297] = i[35];
  assign o[18298] = i[35];
  assign o[18299] = i[35];
  assign o[18300] = i[35];
  assign o[18301] = i[35];
  assign o[18302] = i[35];
  assign o[18303] = i[35];
  assign o[18304] = i[35];
  assign o[18305] = i[35];
  assign o[18306] = i[35];
  assign o[18307] = i[35];
  assign o[18308] = i[35];
  assign o[18309] = i[35];
  assign o[18310] = i[35];
  assign o[18311] = i[35];
  assign o[18312] = i[35];
  assign o[18313] = i[35];
  assign o[18314] = i[35];
  assign o[18315] = i[35];
  assign o[18316] = i[35];
  assign o[18317] = i[35];
  assign o[18318] = i[35];
  assign o[18319] = i[35];
  assign o[18320] = i[35];
  assign o[18321] = i[35];
  assign o[18322] = i[35];
  assign o[18323] = i[35];
  assign o[18324] = i[35];
  assign o[18325] = i[35];
  assign o[18326] = i[35];
  assign o[18327] = i[35];
  assign o[18328] = i[35];
  assign o[18329] = i[35];
  assign o[18330] = i[35];
  assign o[18331] = i[35];
  assign o[18332] = i[35];
  assign o[18333] = i[35];
  assign o[18334] = i[35];
  assign o[18335] = i[35];
  assign o[18336] = i[35];
  assign o[18337] = i[35];
  assign o[18338] = i[35];
  assign o[18339] = i[35];
  assign o[18340] = i[35];
  assign o[18341] = i[35];
  assign o[18342] = i[35];
  assign o[18343] = i[35];
  assign o[18344] = i[35];
  assign o[18345] = i[35];
  assign o[18346] = i[35];
  assign o[18347] = i[35];
  assign o[18348] = i[35];
  assign o[18349] = i[35];
  assign o[18350] = i[35];
  assign o[18351] = i[35];
  assign o[18352] = i[35];
  assign o[18353] = i[35];
  assign o[18354] = i[35];
  assign o[18355] = i[35];
  assign o[18356] = i[35];
  assign o[18357] = i[35];
  assign o[18358] = i[35];
  assign o[18359] = i[35];
  assign o[18360] = i[35];
  assign o[18361] = i[35];
  assign o[18362] = i[35];
  assign o[18363] = i[35];
  assign o[18364] = i[35];
  assign o[18365] = i[35];
  assign o[18366] = i[35];
  assign o[18367] = i[35];
  assign o[18368] = i[35];
  assign o[18369] = i[35];
  assign o[18370] = i[35];
  assign o[18371] = i[35];
  assign o[18372] = i[35];
  assign o[18373] = i[35];
  assign o[18374] = i[35];
  assign o[18375] = i[35];
  assign o[18376] = i[35];
  assign o[18377] = i[35];
  assign o[18378] = i[35];
  assign o[18379] = i[35];
  assign o[18380] = i[35];
  assign o[18381] = i[35];
  assign o[18382] = i[35];
  assign o[18383] = i[35];
  assign o[18384] = i[35];
  assign o[18385] = i[35];
  assign o[18386] = i[35];
  assign o[18387] = i[35];
  assign o[18388] = i[35];
  assign o[18389] = i[35];
  assign o[18390] = i[35];
  assign o[18391] = i[35];
  assign o[18392] = i[35];
  assign o[18393] = i[35];
  assign o[18394] = i[35];
  assign o[18395] = i[35];
  assign o[18396] = i[35];
  assign o[18397] = i[35];
  assign o[18398] = i[35];
  assign o[18399] = i[35];
  assign o[18400] = i[35];
  assign o[18401] = i[35];
  assign o[18402] = i[35];
  assign o[18403] = i[35];
  assign o[18404] = i[35];
  assign o[18405] = i[35];
  assign o[18406] = i[35];
  assign o[18407] = i[35];
  assign o[18408] = i[35];
  assign o[18409] = i[35];
  assign o[18410] = i[35];
  assign o[18411] = i[35];
  assign o[18412] = i[35];
  assign o[18413] = i[35];
  assign o[18414] = i[35];
  assign o[18415] = i[35];
  assign o[18416] = i[35];
  assign o[18417] = i[35];
  assign o[18418] = i[35];
  assign o[18419] = i[35];
  assign o[18420] = i[35];
  assign o[18421] = i[35];
  assign o[18422] = i[35];
  assign o[18423] = i[35];
  assign o[18424] = i[35];
  assign o[18425] = i[35];
  assign o[18426] = i[35];
  assign o[18427] = i[35];
  assign o[18428] = i[35];
  assign o[18429] = i[35];
  assign o[18430] = i[35];
  assign o[18431] = i[35];
  assign o[17408] = i[34];
  assign o[17409] = i[34];
  assign o[17410] = i[34];
  assign o[17411] = i[34];
  assign o[17412] = i[34];
  assign o[17413] = i[34];
  assign o[17414] = i[34];
  assign o[17415] = i[34];
  assign o[17416] = i[34];
  assign o[17417] = i[34];
  assign o[17418] = i[34];
  assign o[17419] = i[34];
  assign o[17420] = i[34];
  assign o[17421] = i[34];
  assign o[17422] = i[34];
  assign o[17423] = i[34];
  assign o[17424] = i[34];
  assign o[17425] = i[34];
  assign o[17426] = i[34];
  assign o[17427] = i[34];
  assign o[17428] = i[34];
  assign o[17429] = i[34];
  assign o[17430] = i[34];
  assign o[17431] = i[34];
  assign o[17432] = i[34];
  assign o[17433] = i[34];
  assign o[17434] = i[34];
  assign o[17435] = i[34];
  assign o[17436] = i[34];
  assign o[17437] = i[34];
  assign o[17438] = i[34];
  assign o[17439] = i[34];
  assign o[17440] = i[34];
  assign o[17441] = i[34];
  assign o[17442] = i[34];
  assign o[17443] = i[34];
  assign o[17444] = i[34];
  assign o[17445] = i[34];
  assign o[17446] = i[34];
  assign o[17447] = i[34];
  assign o[17448] = i[34];
  assign o[17449] = i[34];
  assign o[17450] = i[34];
  assign o[17451] = i[34];
  assign o[17452] = i[34];
  assign o[17453] = i[34];
  assign o[17454] = i[34];
  assign o[17455] = i[34];
  assign o[17456] = i[34];
  assign o[17457] = i[34];
  assign o[17458] = i[34];
  assign o[17459] = i[34];
  assign o[17460] = i[34];
  assign o[17461] = i[34];
  assign o[17462] = i[34];
  assign o[17463] = i[34];
  assign o[17464] = i[34];
  assign o[17465] = i[34];
  assign o[17466] = i[34];
  assign o[17467] = i[34];
  assign o[17468] = i[34];
  assign o[17469] = i[34];
  assign o[17470] = i[34];
  assign o[17471] = i[34];
  assign o[17472] = i[34];
  assign o[17473] = i[34];
  assign o[17474] = i[34];
  assign o[17475] = i[34];
  assign o[17476] = i[34];
  assign o[17477] = i[34];
  assign o[17478] = i[34];
  assign o[17479] = i[34];
  assign o[17480] = i[34];
  assign o[17481] = i[34];
  assign o[17482] = i[34];
  assign o[17483] = i[34];
  assign o[17484] = i[34];
  assign o[17485] = i[34];
  assign o[17486] = i[34];
  assign o[17487] = i[34];
  assign o[17488] = i[34];
  assign o[17489] = i[34];
  assign o[17490] = i[34];
  assign o[17491] = i[34];
  assign o[17492] = i[34];
  assign o[17493] = i[34];
  assign o[17494] = i[34];
  assign o[17495] = i[34];
  assign o[17496] = i[34];
  assign o[17497] = i[34];
  assign o[17498] = i[34];
  assign o[17499] = i[34];
  assign o[17500] = i[34];
  assign o[17501] = i[34];
  assign o[17502] = i[34];
  assign o[17503] = i[34];
  assign o[17504] = i[34];
  assign o[17505] = i[34];
  assign o[17506] = i[34];
  assign o[17507] = i[34];
  assign o[17508] = i[34];
  assign o[17509] = i[34];
  assign o[17510] = i[34];
  assign o[17511] = i[34];
  assign o[17512] = i[34];
  assign o[17513] = i[34];
  assign o[17514] = i[34];
  assign o[17515] = i[34];
  assign o[17516] = i[34];
  assign o[17517] = i[34];
  assign o[17518] = i[34];
  assign o[17519] = i[34];
  assign o[17520] = i[34];
  assign o[17521] = i[34];
  assign o[17522] = i[34];
  assign o[17523] = i[34];
  assign o[17524] = i[34];
  assign o[17525] = i[34];
  assign o[17526] = i[34];
  assign o[17527] = i[34];
  assign o[17528] = i[34];
  assign o[17529] = i[34];
  assign o[17530] = i[34];
  assign o[17531] = i[34];
  assign o[17532] = i[34];
  assign o[17533] = i[34];
  assign o[17534] = i[34];
  assign o[17535] = i[34];
  assign o[17536] = i[34];
  assign o[17537] = i[34];
  assign o[17538] = i[34];
  assign o[17539] = i[34];
  assign o[17540] = i[34];
  assign o[17541] = i[34];
  assign o[17542] = i[34];
  assign o[17543] = i[34];
  assign o[17544] = i[34];
  assign o[17545] = i[34];
  assign o[17546] = i[34];
  assign o[17547] = i[34];
  assign o[17548] = i[34];
  assign o[17549] = i[34];
  assign o[17550] = i[34];
  assign o[17551] = i[34];
  assign o[17552] = i[34];
  assign o[17553] = i[34];
  assign o[17554] = i[34];
  assign o[17555] = i[34];
  assign o[17556] = i[34];
  assign o[17557] = i[34];
  assign o[17558] = i[34];
  assign o[17559] = i[34];
  assign o[17560] = i[34];
  assign o[17561] = i[34];
  assign o[17562] = i[34];
  assign o[17563] = i[34];
  assign o[17564] = i[34];
  assign o[17565] = i[34];
  assign o[17566] = i[34];
  assign o[17567] = i[34];
  assign o[17568] = i[34];
  assign o[17569] = i[34];
  assign o[17570] = i[34];
  assign o[17571] = i[34];
  assign o[17572] = i[34];
  assign o[17573] = i[34];
  assign o[17574] = i[34];
  assign o[17575] = i[34];
  assign o[17576] = i[34];
  assign o[17577] = i[34];
  assign o[17578] = i[34];
  assign o[17579] = i[34];
  assign o[17580] = i[34];
  assign o[17581] = i[34];
  assign o[17582] = i[34];
  assign o[17583] = i[34];
  assign o[17584] = i[34];
  assign o[17585] = i[34];
  assign o[17586] = i[34];
  assign o[17587] = i[34];
  assign o[17588] = i[34];
  assign o[17589] = i[34];
  assign o[17590] = i[34];
  assign o[17591] = i[34];
  assign o[17592] = i[34];
  assign o[17593] = i[34];
  assign o[17594] = i[34];
  assign o[17595] = i[34];
  assign o[17596] = i[34];
  assign o[17597] = i[34];
  assign o[17598] = i[34];
  assign o[17599] = i[34];
  assign o[17600] = i[34];
  assign o[17601] = i[34];
  assign o[17602] = i[34];
  assign o[17603] = i[34];
  assign o[17604] = i[34];
  assign o[17605] = i[34];
  assign o[17606] = i[34];
  assign o[17607] = i[34];
  assign o[17608] = i[34];
  assign o[17609] = i[34];
  assign o[17610] = i[34];
  assign o[17611] = i[34];
  assign o[17612] = i[34];
  assign o[17613] = i[34];
  assign o[17614] = i[34];
  assign o[17615] = i[34];
  assign o[17616] = i[34];
  assign o[17617] = i[34];
  assign o[17618] = i[34];
  assign o[17619] = i[34];
  assign o[17620] = i[34];
  assign o[17621] = i[34];
  assign o[17622] = i[34];
  assign o[17623] = i[34];
  assign o[17624] = i[34];
  assign o[17625] = i[34];
  assign o[17626] = i[34];
  assign o[17627] = i[34];
  assign o[17628] = i[34];
  assign o[17629] = i[34];
  assign o[17630] = i[34];
  assign o[17631] = i[34];
  assign o[17632] = i[34];
  assign o[17633] = i[34];
  assign o[17634] = i[34];
  assign o[17635] = i[34];
  assign o[17636] = i[34];
  assign o[17637] = i[34];
  assign o[17638] = i[34];
  assign o[17639] = i[34];
  assign o[17640] = i[34];
  assign o[17641] = i[34];
  assign o[17642] = i[34];
  assign o[17643] = i[34];
  assign o[17644] = i[34];
  assign o[17645] = i[34];
  assign o[17646] = i[34];
  assign o[17647] = i[34];
  assign o[17648] = i[34];
  assign o[17649] = i[34];
  assign o[17650] = i[34];
  assign o[17651] = i[34];
  assign o[17652] = i[34];
  assign o[17653] = i[34];
  assign o[17654] = i[34];
  assign o[17655] = i[34];
  assign o[17656] = i[34];
  assign o[17657] = i[34];
  assign o[17658] = i[34];
  assign o[17659] = i[34];
  assign o[17660] = i[34];
  assign o[17661] = i[34];
  assign o[17662] = i[34];
  assign o[17663] = i[34];
  assign o[17664] = i[34];
  assign o[17665] = i[34];
  assign o[17666] = i[34];
  assign o[17667] = i[34];
  assign o[17668] = i[34];
  assign o[17669] = i[34];
  assign o[17670] = i[34];
  assign o[17671] = i[34];
  assign o[17672] = i[34];
  assign o[17673] = i[34];
  assign o[17674] = i[34];
  assign o[17675] = i[34];
  assign o[17676] = i[34];
  assign o[17677] = i[34];
  assign o[17678] = i[34];
  assign o[17679] = i[34];
  assign o[17680] = i[34];
  assign o[17681] = i[34];
  assign o[17682] = i[34];
  assign o[17683] = i[34];
  assign o[17684] = i[34];
  assign o[17685] = i[34];
  assign o[17686] = i[34];
  assign o[17687] = i[34];
  assign o[17688] = i[34];
  assign o[17689] = i[34];
  assign o[17690] = i[34];
  assign o[17691] = i[34];
  assign o[17692] = i[34];
  assign o[17693] = i[34];
  assign o[17694] = i[34];
  assign o[17695] = i[34];
  assign o[17696] = i[34];
  assign o[17697] = i[34];
  assign o[17698] = i[34];
  assign o[17699] = i[34];
  assign o[17700] = i[34];
  assign o[17701] = i[34];
  assign o[17702] = i[34];
  assign o[17703] = i[34];
  assign o[17704] = i[34];
  assign o[17705] = i[34];
  assign o[17706] = i[34];
  assign o[17707] = i[34];
  assign o[17708] = i[34];
  assign o[17709] = i[34];
  assign o[17710] = i[34];
  assign o[17711] = i[34];
  assign o[17712] = i[34];
  assign o[17713] = i[34];
  assign o[17714] = i[34];
  assign o[17715] = i[34];
  assign o[17716] = i[34];
  assign o[17717] = i[34];
  assign o[17718] = i[34];
  assign o[17719] = i[34];
  assign o[17720] = i[34];
  assign o[17721] = i[34];
  assign o[17722] = i[34];
  assign o[17723] = i[34];
  assign o[17724] = i[34];
  assign o[17725] = i[34];
  assign o[17726] = i[34];
  assign o[17727] = i[34];
  assign o[17728] = i[34];
  assign o[17729] = i[34];
  assign o[17730] = i[34];
  assign o[17731] = i[34];
  assign o[17732] = i[34];
  assign o[17733] = i[34];
  assign o[17734] = i[34];
  assign o[17735] = i[34];
  assign o[17736] = i[34];
  assign o[17737] = i[34];
  assign o[17738] = i[34];
  assign o[17739] = i[34];
  assign o[17740] = i[34];
  assign o[17741] = i[34];
  assign o[17742] = i[34];
  assign o[17743] = i[34];
  assign o[17744] = i[34];
  assign o[17745] = i[34];
  assign o[17746] = i[34];
  assign o[17747] = i[34];
  assign o[17748] = i[34];
  assign o[17749] = i[34];
  assign o[17750] = i[34];
  assign o[17751] = i[34];
  assign o[17752] = i[34];
  assign o[17753] = i[34];
  assign o[17754] = i[34];
  assign o[17755] = i[34];
  assign o[17756] = i[34];
  assign o[17757] = i[34];
  assign o[17758] = i[34];
  assign o[17759] = i[34];
  assign o[17760] = i[34];
  assign o[17761] = i[34];
  assign o[17762] = i[34];
  assign o[17763] = i[34];
  assign o[17764] = i[34];
  assign o[17765] = i[34];
  assign o[17766] = i[34];
  assign o[17767] = i[34];
  assign o[17768] = i[34];
  assign o[17769] = i[34];
  assign o[17770] = i[34];
  assign o[17771] = i[34];
  assign o[17772] = i[34];
  assign o[17773] = i[34];
  assign o[17774] = i[34];
  assign o[17775] = i[34];
  assign o[17776] = i[34];
  assign o[17777] = i[34];
  assign o[17778] = i[34];
  assign o[17779] = i[34];
  assign o[17780] = i[34];
  assign o[17781] = i[34];
  assign o[17782] = i[34];
  assign o[17783] = i[34];
  assign o[17784] = i[34];
  assign o[17785] = i[34];
  assign o[17786] = i[34];
  assign o[17787] = i[34];
  assign o[17788] = i[34];
  assign o[17789] = i[34];
  assign o[17790] = i[34];
  assign o[17791] = i[34];
  assign o[17792] = i[34];
  assign o[17793] = i[34];
  assign o[17794] = i[34];
  assign o[17795] = i[34];
  assign o[17796] = i[34];
  assign o[17797] = i[34];
  assign o[17798] = i[34];
  assign o[17799] = i[34];
  assign o[17800] = i[34];
  assign o[17801] = i[34];
  assign o[17802] = i[34];
  assign o[17803] = i[34];
  assign o[17804] = i[34];
  assign o[17805] = i[34];
  assign o[17806] = i[34];
  assign o[17807] = i[34];
  assign o[17808] = i[34];
  assign o[17809] = i[34];
  assign o[17810] = i[34];
  assign o[17811] = i[34];
  assign o[17812] = i[34];
  assign o[17813] = i[34];
  assign o[17814] = i[34];
  assign o[17815] = i[34];
  assign o[17816] = i[34];
  assign o[17817] = i[34];
  assign o[17818] = i[34];
  assign o[17819] = i[34];
  assign o[17820] = i[34];
  assign o[17821] = i[34];
  assign o[17822] = i[34];
  assign o[17823] = i[34];
  assign o[17824] = i[34];
  assign o[17825] = i[34];
  assign o[17826] = i[34];
  assign o[17827] = i[34];
  assign o[17828] = i[34];
  assign o[17829] = i[34];
  assign o[17830] = i[34];
  assign o[17831] = i[34];
  assign o[17832] = i[34];
  assign o[17833] = i[34];
  assign o[17834] = i[34];
  assign o[17835] = i[34];
  assign o[17836] = i[34];
  assign o[17837] = i[34];
  assign o[17838] = i[34];
  assign o[17839] = i[34];
  assign o[17840] = i[34];
  assign o[17841] = i[34];
  assign o[17842] = i[34];
  assign o[17843] = i[34];
  assign o[17844] = i[34];
  assign o[17845] = i[34];
  assign o[17846] = i[34];
  assign o[17847] = i[34];
  assign o[17848] = i[34];
  assign o[17849] = i[34];
  assign o[17850] = i[34];
  assign o[17851] = i[34];
  assign o[17852] = i[34];
  assign o[17853] = i[34];
  assign o[17854] = i[34];
  assign o[17855] = i[34];
  assign o[17856] = i[34];
  assign o[17857] = i[34];
  assign o[17858] = i[34];
  assign o[17859] = i[34];
  assign o[17860] = i[34];
  assign o[17861] = i[34];
  assign o[17862] = i[34];
  assign o[17863] = i[34];
  assign o[17864] = i[34];
  assign o[17865] = i[34];
  assign o[17866] = i[34];
  assign o[17867] = i[34];
  assign o[17868] = i[34];
  assign o[17869] = i[34];
  assign o[17870] = i[34];
  assign o[17871] = i[34];
  assign o[17872] = i[34];
  assign o[17873] = i[34];
  assign o[17874] = i[34];
  assign o[17875] = i[34];
  assign o[17876] = i[34];
  assign o[17877] = i[34];
  assign o[17878] = i[34];
  assign o[17879] = i[34];
  assign o[17880] = i[34];
  assign o[17881] = i[34];
  assign o[17882] = i[34];
  assign o[17883] = i[34];
  assign o[17884] = i[34];
  assign o[17885] = i[34];
  assign o[17886] = i[34];
  assign o[17887] = i[34];
  assign o[17888] = i[34];
  assign o[17889] = i[34];
  assign o[17890] = i[34];
  assign o[17891] = i[34];
  assign o[17892] = i[34];
  assign o[17893] = i[34];
  assign o[17894] = i[34];
  assign o[17895] = i[34];
  assign o[17896] = i[34];
  assign o[17897] = i[34];
  assign o[17898] = i[34];
  assign o[17899] = i[34];
  assign o[17900] = i[34];
  assign o[17901] = i[34];
  assign o[17902] = i[34];
  assign o[17903] = i[34];
  assign o[17904] = i[34];
  assign o[17905] = i[34];
  assign o[17906] = i[34];
  assign o[17907] = i[34];
  assign o[17908] = i[34];
  assign o[17909] = i[34];
  assign o[17910] = i[34];
  assign o[17911] = i[34];
  assign o[17912] = i[34];
  assign o[17913] = i[34];
  assign o[17914] = i[34];
  assign o[17915] = i[34];
  assign o[17916] = i[34];
  assign o[17917] = i[34];
  assign o[17918] = i[34];
  assign o[17919] = i[34];
  assign o[16896] = i[33];
  assign o[16897] = i[33];
  assign o[16898] = i[33];
  assign o[16899] = i[33];
  assign o[16900] = i[33];
  assign o[16901] = i[33];
  assign o[16902] = i[33];
  assign o[16903] = i[33];
  assign o[16904] = i[33];
  assign o[16905] = i[33];
  assign o[16906] = i[33];
  assign o[16907] = i[33];
  assign o[16908] = i[33];
  assign o[16909] = i[33];
  assign o[16910] = i[33];
  assign o[16911] = i[33];
  assign o[16912] = i[33];
  assign o[16913] = i[33];
  assign o[16914] = i[33];
  assign o[16915] = i[33];
  assign o[16916] = i[33];
  assign o[16917] = i[33];
  assign o[16918] = i[33];
  assign o[16919] = i[33];
  assign o[16920] = i[33];
  assign o[16921] = i[33];
  assign o[16922] = i[33];
  assign o[16923] = i[33];
  assign o[16924] = i[33];
  assign o[16925] = i[33];
  assign o[16926] = i[33];
  assign o[16927] = i[33];
  assign o[16928] = i[33];
  assign o[16929] = i[33];
  assign o[16930] = i[33];
  assign o[16931] = i[33];
  assign o[16932] = i[33];
  assign o[16933] = i[33];
  assign o[16934] = i[33];
  assign o[16935] = i[33];
  assign o[16936] = i[33];
  assign o[16937] = i[33];
  assign o[16938] = i[33];
  assign o[16939] = i[33];
  assign o[16940] = i[33];
  assign o[16941] = i[33];
  assign o[16942] = i[33];
  assign o[16943] = i[33];
  assign o[16944] = i[33];
  assign o[16945] = i[33];
  assign o[16946] = i[33];
  assign o[16947] = i[33];
  assign o[16948] = i[33];
  assign o[16949] = i[33];
  assign o[16950] = i[33];
  assign o[16951] = i[33];
  assign o[16952] = i[33];
  assign o[16953] = i[33];
  assign o[16954] = i[33];
  assign o[16955] = i[33];
  assign o[16956] = i[33];
  assign o[16957] = i[33];
  assign o[16958] = i[33];
  assign o[16959] = i[33];
  assign o[16960] = i[33];
  assign o[16961] = i[33];
  assign o[16962] = i[33];
  assign o[16963] = i[33];
  assign o[16964] = i[33];
  assign o[16965] = i[33];
  assign o[16966] = i[33];
  assign o[16967] = i[33];
  assign o[16968] = i[33];
  assign o[16969] = i[33];
  assign o[16970] = i[33];
  assign o[16971] = i[33];
  assign o[16972] = i[33];
  assign o[16973] = i[33];
  assign o[16974] = i[33];
  assign o[16975] = i[33];
  assign o[16976] = i[33];
  assign o[16977] = i[33];
  assign o[16978] = i[33];
  assign o[16979] = i[33];
  assign o[16980] = i[33];
  assign o[16981] = i[33];
  assign o[16982] = i[33];
  assign o[16983] = i[33];
  assign o[16984] = i[33];
  assign o[16985] = i[33];
  assign o[16986] = i[33];
  assign o[16987] = i[33];
  assign o[16988] = i[33];
  assign o[16989] = i[33];
  assign o[16990] = i[33];
  assign o[16991] = i[33];
  assign o[16992] = i[33];
  assign o[16993] = i[33];
  assign o[16994] = i[33];
  assign o[16995] = i[33];
  assign o[16996] = i[33];
  assign o[16997] = i[33];
  assign o[16998] = i[33];
  assign o[16999] = i[33];
  assign o[17000] = i[33];
  assign o[17001] = i[33];
  assign o[17002] = i[33];
  assign o[17003] = i[33];
  assign o[17004] = i[33];
  assign o[17005] = i[33];
  assign o[17006] = i[33];
  assign o[17007] = i[33];
  assign o[17008] = i[33];
  assign o[17009] = i[33];
  assign o[17010] = i[33];
  assign o[17011] = i[33];
  assign o[17012] = i[33];
  assign o[17013] = i[33];
  assign o[17014] = i[33];
  assign o[17015] = i[33];
  assign o[17016] = i[33];
  assign o[17017] = i[33];
  assign o[17018] = i[33];
  assign o[17019] = i[33];
  assign o[17020] = i[33];
  assign o[17021] = i[33];
  assign o[17022] = i[33];
  assign o[17023] = i[33];
  assign o[17024] = i[33];
  assign o[17025] = i[33];
  assign o[17026] = i[33];
  assign o[17027] = i[33];
  assign o[17028] = i[33];
  assign o[17029] = i[33];
  assign o[17030] = i[33];
  assign o[17031] = i[33];
  assign o[17032] = i[33];
  assign o[17033] = i[33];
  assign o[17034] = i[33];
  assign o[17035] = i[33];
  assign o[17036] = i[33];
  assign o[17037] = i[33];
  assign o[17038] = i[33];
  assign o[17039] = i[33];
  assign o[17040] = i[33];
  assign o[17041] = i[33];
  assign o[17042] = i[33];
  assign o[17043] = i[33];
  assign o[17044] = i[33];
  assign o[17045] = i[33];
  assign o[17046] = i[33];
  assign o[17047] = i[33];
  assign o[17048] = i[33];
  assign o[17049] = i[33];
  assign o[17050] = i[33];
  assign o[17051] = i[33];
  assign o[17052] = i[33];
  assign o[17053] = i[33];
  assign o[17054] = i[33];
  assign o[17055] = i[33];
  assign o[17056] = i[33];
  assign o[17057] = i[33];
  assign o[17058] = i[33];
  assign o[17059] = i[33];
  assign o[17060] = i[33];
  assign o[17061] = i[33];
  assign o[17062] = i[33];
  assign o[17063] = i[33];
  assign o[17064] = i[33];
  assign o[17065] = i[33];
  assign o[17066] = i[33];
  assign o[17067] = i[33];
  assign o[17068] = i[33];
  assign o[17069] = i[33];
  assign o[17070] = i[33];
  assign o[17071] = i[33];
  assign o[17072] = i[33];
  assign o[17073] = i[33];
  assign o[17074] = i[33];
  assign o[17075] = i[33];
  assign o[17076] = i[33];
  assign o[17077] = i[33];
  assign o[17078] = i[33];
  assign o[17079] = i[33];
  assign o[17080] = i[33];
  assign o[17081] = i[33];
  assign o[17082] = i[33];
  assign o[17083] = i[33];
  assign o[17084] = i[33];
  assign o[17085] = i[33];
  assign o[17086] = i[33];
  assign o[17087] = i[33];
  assign o[17088] = i[33];
  assign o[17089] = i[33];
  assign o[17090] = i[33];
  assign o[17091] = i[33];
  assign o[17092] = i[33];
  assign o[17093] = i[33];
  assign o[17094] = i[33];
  assign o[17095] = i[33];
  assign o[17096] = i[33];
  assign o[17097] = i[33];
  assign o[17098] = i[33];
  assign o[17099] = i[33];
  assign o[17100] = i[33];
  assign o[17101] = i[33];
  assign o[17102] = i[33];
  assign o[17103] = i[33];
  assign o[17104] = i[33];
  assign o[17105] = i[33];
  assign o[17106] = i[33];
  assign o[17107] = i[33];
  assign o[17108] = i[33];
  assign o[17109] = i[33];
  assign o[17110] = i[33];
  assign o[17111] = i[33];
  assign o[17112] = i[33];
  assign o[17113] = i[33];
  assign o[17114] = i[33];
  assign o[17115] = i[33];
  assign o[17116] = i[33];
  assign o[17117] = i[33];
  assign o[17118] = i[33];
  assign o[17119] = i[33];
  assign o[17120] = i[33];
  assign o[17121] = i[33];
  assign o[17122] = i[33];
  assign o[17123] = i[33];
  assign o[17124] = i[33];
  assign o[17125] = i[33];
  assign o[17126] = i[33];
  assign o[17127] = i[33];
  assign o[17128] = i[33];
  assign o[17129] = i[33];
  assign o[17130] = i[33];
  assign o[17131] = i[33];
  assign o[17132] = i[33];
  assign o[17133] = i[33];
  assign o[17134] = i[33];
  assign o[17135] = i[33];
  assign o[17136] = i[33];
  assign o[17137] = i[33];
  assign o[17138] = i[33];
  assign o[17139] = i[33];
  assign o[17140] = i[33];
  assign o[17141] = i[33];
  assign o[17142] = i[33];
  assign o[17143] = i[33];
  assign o[17144] = i[33];
  assign o[17145] = i[33];
  assign o[17146] = i[33];
  assign o[17147] = i[33];
  assign o[17148] = i[33];
  assign o[17149] = i[33];
  assign o[17150] = i[33];
  assign o[17151] = i[33];
  assign o[17152] = i[33];
  assign o[17153] = i[33];
  assign o[17154] = i[33];
  assign o[17155] = i[33];
  assign o[17156] = i[33];
  assign o[17157] = i[33];
  assign o[17158] = i[33];
  assign o[17159] = i[33];
  assign o[17160] = i[33];
  assign o[17161] = i[33];
  assign o[17162] = i[33];
  assign o[17163] = i[33];
  assign o[17164] = i[33];
  assign o[17165] = i[33];
  assign o[17166] = i[33];
  assign o[17167] = i[33];
  assign o[17168] = i[33];
  assign o[17169] = i[33];
  assign o[17170] = i[33];
  assign o[17171] = i[33];
  assign o[17172] = i[33];
  assign o[17173] = i[33];
  assign o[17174] = i[33];
  assign o[17175] = i[33];
  assign o[17176] = i[33];
  assign o[17177] = i[33];
  assign o[17178] = i[33];
  assign o[17179] = i[33];
  assign o[17180] = i[33];
  assign o[17181] = i[33];
  assign o[17182] = i[33];
  assign o[17183] = i[33];
  assign o[17184] = i[33];
  assign o[17185] = i[33];
  assign o[17186] = i[33];
  assign o[17187] = i[33];
  assign o[17188] = i[33];
  assign o[17189] = i[33];
  assign o[17190] = i[33];
  assign o[17191] = i[33];
  assign o[17192] = i[33];
  assign o[17193] = i[33];
  assign o[17194] = i[33];
  assign o[17195] = i[33];
  assign o[17196] = i[33];
  assign o[17197] = i[33];
  assign o[17198] = i[33];
  assign o[17199] = i[33];
  assign o[17200] = i[33];
  assign o[17201] = i[33];
  assign o[17202] = i[33];
  assign o[17203] = i[33];
  assign o[17204] = i[33];
  assign o[17205] = i[33];
  assign o[17206] = i[33];
  assign o[17207] = i[33];
  assign o[17208] = i[33];
  assign o[17209] = i[33];
  assign o[17210] = i[33];
  assign o[17211] = i[33];
  assign o[17212] = i[33];
  assign o[17213] = i[33];
  assign o[17214] = i[33];
  assign o[17215] = i[33];
  assign o[17216] = i[33];
  assign o[17217] = i[33];
  assign o[17218] = i[33];
  assign o[17219] = i[33];
  assign o[17220] = i[33];
  assign o[17221] = i[33];
  assign o[17222] = i[33];
  assign o[17223] = i[33];
  assign o[17224] = i[33];
  assign o[17225] = i[33];
  assign o[17226] = i[33];
  assign o[17227] = i[33];
  assign o[17228] = i[33];
  assign o[17229] = i[33];
  assign o[17230] = i[33];
  assign o[17231] = i[33];
  assign o[17232] = i[33];
  assign o[17233] = i[33];
  assign o[17234] = i[33];
  assign o[17235] = i[33];
  assign o[17236] = i[33];
  assign o[17237] = i[33];
  assign o[17238] = i[33];
  assign o[17239] = i[33];
  assign o[17240] = i[33];
  assign o[17241] = i[33];
  assign o[17242] = i[33];
  assign o[17243] = i[33];
  assign o[17244] = i[33];
  assign o[17245] = i[33];
  assign o[17246] = i[33];
  assign o[17247] = i[33];
  assign o[17248] = i[33];
  assign o[17249] = i[33];
  assign o[17250] = i[33];
  assign o[17251] = i[33];
  assign o[17252] = i[33];
  assign o[17253] = i[33];
  assign o[17254] = i[33];
  assign o[17255] = i[33];
  assign o[17256] = i[33];
  assign o[17257] = i[33];
  assign o[17258] = i[33];
  assign o[17259] = i[33];
  assign o[17260] = i[33];
  assign o[17261] = i[33];
  assign o[17262] = i[33];
  assign o[17263] = i[33];
  assign o[17264] = i[33];
  assign o[17265] = i[33];
  assign o[17266] = i[33];
  assign o[17267] = i[33];
  assign o[17268] = i[33];
  assign o[17269] = i[33];
  assign o[17270] = i[33];
  assign o[17271] = i[33];
  assign o[17272] = i[33];
  assign o[17273] = i[33];
  assign o[17274] = i[33];
  assign o[17275] = i[33];
  assign o[17276] = i[33];
  assign o[17277] = i[33];
  assign o[17278] = i[33];
  assign o[17279] = i[33];
  assign o[17280] = i[33];
  assign o[17281] = i[33];
  assign o[17282] = i[33];
  assign o[17283] = i[33];
  assign o[17284] = i[33];
  assign o[17285] = i[33];
  assign o[17286] = i[33];
  assign o[17287] = i[33];
  assign o[17288] = i[33];
  assign o[17289] = i[33];
  assign o[17290] = i[33];
  assign o[17291] = i[33];
  assign o[17292] = i[33];
  assign o[17293] = i[33];
  assign o[17294] = i[33];
  assign o[17295] = i[33];
  assign o[17296] = i[33];
  assign o[17297] = i[33];
  assign o[17298] = i[33];
  assign o[17299] = i[33];
  assign o[17300] = i[33];
  assign o[17301] = i[33];
  assign o[17302] = i[33];
  assign o[17303] = i[33];
  assign o[17304] = i[33];
  assign o[17305] = i[33];
  assign o[17306] = i[33];
  assign o[17307] = i[33];
  assign o[17308] = i[33];
  assign o[17309] = i[33];
  assign o[17310] = i[33];
  assign o[17311] = i[33];
  assign o[17312] = i[33];
  assign o[17313] = i[33];
  assign o[17314] = i[33];
  assign o[17315] = i[33];
  assign o[17316] = i[33];
  assign o[17317] = i[33];
  assign o[17318] = i[33];
  assign o[17319] = i[33];
  assign o[17320] = i[33];
  assign o[17321] = i[33];
  assign o[17322] = i[33];
  assign o[17323] = i[33];
  assign o[17324] = i[33];
  assign o[17325] = i[33];
  assign o[17326] = i[33];
  assign o[17327] = i[33];
  assign o[17328] = i[33];
  assign o[17329] = i[33];
  assign o[17330] = i[33];
  assign o[17331] = i[33];
  assign o[17332] = i[33];
  assign o[17333] = i[33];
  assign o[17334] = i[33];
  assign o[17335] = i[33];
  assign o[17336] = i[33];
  assign o[17337] = i[33];
  assign o[17338] = i[33];
  assign o[17339] = i[33];
  assign o[17340] = i[33];
  assign o[17341] = i[33];
  assign o[17342] = i[33];
  assign o[17343] = i[33];
  assign o[17344] = i[33];
  assign o[17345] = i[33];
  assign o[17346] = i[33];
  assign o[17347] = i[33];
  assign o[17348] = i[33];
  assign o[17349] = i[33];
  assign o[17350] = i[33];
  assign o[17351] = i[33];
  assign o[17352] = i[33];
  assign o[17353] = i[33];
  assign o[17354] = i[33];
  assign o[17355] = i[33];
  assign o[17356] = i[33];
  assign o[17357] = i[33];
  assign o[17358] = i[33];
  assign o[17359] = i[33];
  assign o[17360] = i[33];
  assign o[17361] = i[33];
  assign o[17362] = i[33];
  assign o[17363] = i[33];
  assign o[17364] = i[33];
  assign o[17365] = i[33];
  assign o[17366] = i[33];
  assign o[17367] = i[33];
  assign o[17368] = i[33];
  assign o[17369] = i[33];
  assign o[17370] = i[33];
  assign o[17371] = i[33];
  assign o[17372] = i[33];
  assign o[17373] = i[33];
  assign o[17374] = i[33];
  assign o[17375] = i[33];
  assign o[17376] = i[33];
  assign o[17377] = i[33];
  assign o[17378] = i[33];
  assign o[17379] = i[33];
  assign o[17380] = i[33];
  assign o[17381] = i[33];
  assign o[17382] = i[33];
  assign o[17383] = i[33];
  assign o[17384] = i[33];
  assign o[17385] = i[33];
  assign o[17386] = i[33];
  assign o[17387] = i[33];
  assign o[17388] = i[33];
  assign o[17389] = i[33];
  assign o[17390] = i[33];
  assign o[17391] = i[33];
  assign o[17392] = i[33];
  assign o[17393] = i[33];
  assign o[17394] = i[33];
  assign o[17395] = i[33];
  assign o[17396] = i[33];
  assign o[17397] = i[33];
  assign o[17398] = i[33];
  assign o[17399] = i[33];
  assign o[17400] = i[33];
  assign o[17401] = i[33];
  assign o[17402] = i[33];
  assign o[17403] = i[33];
  assign o[17404] = i[33];
  assign o[17405] = i[33];
  assign o[17406] = i[33];
  assign o[17407] = i[33];
  assign o[16384] = i[32];
  assign o[16385] = i[32];
  assign o[16386] = i[32];
  assign o[16387] = i[32];
  assign o[16388] = i[32];
  assign o[16389] = i[32];
  assign o[16390] = i[32];
  assign o[16391] = i[32];
  assign o[16392] = i[32];
  assign o[16393] = i[32];
  assign o[16394] = i[32];
  assign o[16395] = i[32];
  assign o[16396] = i[32];
  assign o[16397] = i[32];
  assign o[16398] = i[32];
  assign o[16399] = i[32];
  assign o[16400] = i[32];
  assign o[16401] = i[32];
  assign o[16402] = i[32];
  assign o[16403] = i[32];
  assign o[16404] = i[32];
  assign o[16405] = i[32];
  assign o[16406] = i[32];
  assign o[16407] = i[32];
  assign o[16408] = i[32];
  assign o[16409] = i[32];
  assign o[16410] = i[32];
  assign o[16411] = i[32];
  assign o[16412] = i[32];
  assign o[16413] = i[32];
  assign o[16414] = i[32];
  assign o[16415] = i[32];
  assign o[16416] = i[32];
  assign o[16417] = i[32];
  assign o[16418] = i[32];
  assign o[16419] = i[32];
  assign o[16420] = i[32];
  assign o[16421] = i[32];
  assign o[16422] = i[32];
  assign o[16423] = i[32];
  assign o[16424] = i[32];
  assign o[16425] = i[32];
  assign o[16426] = i[32];
  assign o[16427] = i[32];
  assign o[16428] = i[32];
  assign o[16429] = i[32];
  assign o[16430] = i[32];
  assign o[16431] = i[32];
  assign o[16432] = i[32];
  assign o[16433] = i[32];
  assign o[16434] = i[32];
  assign o[16435] = i[32];
  assign o[16436] = i[32];
  assign o[16437] = i[32];
  assign o[16438] = i[32];
  assign o[16439] = i[32];
  assign o[16440] = i[32];
  assign o[16441] = i[32];
  assign o[16442] = i[32];
  assign o[16443] = i[32];
  assign o[16444] = i[32];
  assign o[16445] = i[32];
  assign o[16446] = i[32];
  assign o[16447] = i[32];
  assign o[16448] = i[32];
  assign o[16449] = i[32];
  assign o[16450] = i[32];
  assign o[16451] = i[32];
  assign o[16452] = i[32];
  assign o[16453] = i[32];
  assign o[16454] = i[32];
  assign o[16455] = i[32];
  assign o[16456] = i[32];
  assign o[16457] = i[32];
  assign o[16458] = i[32];
  assign o[16459] = i[32];
  assign o[16460] = i[32];
  assign o[16461] = i[32];
  assign o[16462] = i[32];
  assign o[16463] = i[32];
  assign o[16464] = i[32];
  assign o[16465] = i[32];
  assign o[16466] = i[32];
  assign o[16467] = i[32];
  assign o[16468] = i[32];
  assign o[16469] = i[32];
  assign o[16470] = i[32];
  assign o[16471] = i[32];
  assign o[16472] = i[32];
  assign o[16473] = i[32];
  assign o[16474] = i[32];
  assign o[16475] = i[32];
  assign o[16476] = i[32];
  assign o[16477] = i[32];
  assign o[16478] = i[32];
  assign o[16479] = i[32];
  assign o[16480] = i[32];
  assign o[16481] = i[32];
  assign o[16482] = i[32];
  assign o[16483] = i[32];
  assign o[16484] = i[32];
  assign o[16485] = i[32];
  assign o[16486] = i[32];
  assign o[16487] = i[32];
  assign o[16488] = i[32];
  assign o[16489] = i[32];
  assign o[16490] = i[32];
  assign o[16491] = i[32];
  assign o[16492] = i[32];
  assign o[16493] = i[32];
  assign o[16494] = i[32];
  assign o[16495] = i[32];
  assign o[16496] = i[32];
  assign o[16497] = i[32];
  assign o[16498] = i[32];
  assign o[16499] = i[32];
  assign o[16500] = i[32];
  assign o[16501] = i[32];
  assign o[16502] = i[32];
  assign o[16503] = i[32];
  assign o[16504] = i[32];
  assign o[16505] = i[32];
  assign o[16506] = i[32];
  assign o[16507] = i[32];
  assign o[16508] = i[32];
  assign o[16509] = i[32];
  assign o[16510] = i[32];
  assign o[16511] = i[32];
  assign o[16512] = i[32];
  assign o[16513] = i[32];
  assign o[16514] = i[32];
  assign o[16515] = i[32];
  assign o[16516] = i[32];
  assign o[16517] = i[32];
  assign o[16518] = i[32];
  assign o[16519] = i[32];
  assign o[16520] = i[32];
  assign o[16521] = i[32];
  assign o[16522] = i[32];
  assign o[16523] = i[32];
  assign o[16524] = i[32];
  assign o[16525] = i[32];
  assign o[16526] = i[32];
  assign o[16527] = i[32];
  assign o[16528] = i[32];
  assign o[16529] = i[32];
  assign o[16530] = i[32];
  assign o[16531] = i[32];
  assign o[16532] = i[32];
  assign o[16533] = i[32];
  assign o[16534] = i[32];
  assign o[16535] = i[32];
  assign o[16536] = i[32];
  assign o[16537] = i[32];
  assign o[16538] = i[32];
  assign o[16539] = i[32];
  assign o[16540] = i[32];
  assign o[16541] = i[32];
  assign o[16542] = i[32];
  assign o[16543] = i[32];
  assign o[16544] = i[32];
  assign o[16545] = i[32];
  assign o[16546] = i[32];
  assign o[16547] = i[32];
  assign o[16548] = i[32];
  assign o[16549] = i[32];
  assign o[16550] = i[32];
  assign o[16551] = i[32];
  assign o[16552] = i[32];
  assign o[16553] = i[32];
  assign o[16554] = i[32];
  assign o[16555] = i[32];
  assign o[16556] = i[32];
  assign o[16557] = i[32];
  assign o[16558] = i[32];
  assign o[16559] = i[32];
  assign o[16560] = i[32];
  assign o[16561] = i[32];
  assign o[16562] = i[32];
  assign o[16563] = i[32];
  assign o[16564] = i[32];
  assign o[16565] = i[32];
  assign o[16566] = i[32];
  assign o[16567] = i[32];
  assign o[16568] = i[32];
  assign o[16569] = i[32];
  assign o[16570] = i[32];
  assign o[16571] = i[32];
  assign o[16572] = i[32];
  assign o[16573] = i[32];
  assign o[16574] = i[32];
  assign o[16575] = i[32];
  assign o[16576] = i[32];
  assign o[16577] = i[32];
  assign o[16578] = i[32];
  assign o[16579] = i[32];
  assign o[16580] = i[32];
  assign o[16581] = i[32];
  assign o[16582] = i[32];
  assign o[16583] = i[32];
  assign o[16584] = i[32];
  assign o[16585] = i[32];
  assign o[16586] = i[32];
  assign o[16587] = i[32];
  assign o[16588] = i[32];
  assign o[16589] = i[32];
  assign o[16590] = i[32];
  assign o[16591] = i[32];
  assign o[16592] = i[32];
  assign o[16593] = i[32];
  assign o[16594] = i[32];
  assign o[16595] = i[32];
  assign o[16596] = i[32];
  assign o[16597] = i[32];
  assign o[16598] = i[32];
  assign o[16599] = i[32];
  assign o[16600] = i[32];
  assign o[16601] = i[32];
  assign o[16602] = i[32];
  assign o[16603] = i[32];
  assign o[16604] = i[32];
  assign o[16605] = i[32];
  assign o[16606] = i[32];
  assign o[16607] = i[32];
  assign o[16608] = i[32];
  assign o[16609] = i[32];
  assign o[16610] = i[32];
  assign o[16611] = i[32];
  assign o[16612] = i[32];
  assign o[16613] = i[32];
  assign o[16614] = i[32];
  assign o[16615] = i[32];
  assign o[16616] = i[32];
  assign o[16617] = i[32];
  assign o[16618] = i[32];
  assign o[16619] = i[32];
  assign o[16620] = i[32];
  assign o[16621] = i[32];
  assign o[16622] = i[32];
  assign o[16623] = i[32];
  assign o[16624] = i[32];
  assign o[16625] = i[32];
  assign o[16626] = i[32];
  assign o[16627] = i[32];
  assign o[16628] = i[32];
  assign o[16629] = i[32];
  assign o[16630] = i[32];
  assign o[16631] = i[32];
  assign o[16632] = i[32];
  assign o[16633] = i[32];
  assign o[16634] = i[32];
  assign o[16635] = i[32];
  assign o[16636] = i[32];
  assign o[16637] = i[32];
  assign o[16638] = i[32];
  assign o[16639] = i[32];
  assign o[16640] = i[32];
  assign o[16641] = i[32];
  assign o[16642] = i[32];
  assign o[16643] = i[32];
  assign o[16644] = i[32];
  assign o[16645] = i[32];
  assign o[16646] = i[32];
  assign o[16647] = i[32];
  assign o[16648] = i[32];
  assign o[16649] = i[32];
  assign o[16650] = i[32];
  assign o[16651] = i[32];
  assign o[16652] = i[32];
  assign o[16653] = i[32];
  assign o[16654] = i[32];
  assign o[16655] = i[32];
  assign o[16656] = i[32];
  assign o[16657] = i[32];
  assign o[16658] = i[32];
  assign o[16659] = i[32];
  assign o[16660] = i[32];
  assign o[16661] = i[32];
  assign o[16662] = i[32];
  assign o[16663] = i[32];
  assign o[16664] = i[32];
  assign o[16665] = i[32];
  assign o[16666] = i[32];
  assign o[16667] = i[32];
  assign o[16668] = i[32];
  assign o[16669] = i[32];
  assign o[16670] = i[32];
  assign o[16671] = i[32];
  assign o[16672] = i[32];
  assign o[16673] = i[32];
  assign o[16674] = i[32];
  assign o[16675] = i[32];
  assign o[16676] = i[32];
  assign o[16677] = i[32];
  assign o[16678] = i[32];
  assign o[16679] = i[32];
  assign o[16680] = i[32];
  assign o[16681] = i[32];
  assign o[16682] = i[32];
  assign o[16683] = i[32];
  assign o[16684] = i[32];
  assign o[16685] = i[32];
  assign o[16686] = i[32];
  assign o[16687] = i[32];
  assign o[16688] = i[32];
  assign o[16689] = i[32];
  assign o[16690] = i[32];
  assign o[16691] = i[32];
  assign o[16692] = i[32];
  assign o[16693] = i[32];
  assign o[16694] = i[32];
  assign o[16695] = i[32];
  assign o[16696] = i[32];
  assign o[16697] = i[32];
  assign o[16698] = i[32];
  assign o[16699] = i[32];
  assign o[16700] = i[32];
  assign o[16701] = i[32];
  assign o[16702] = i[32];
  assign o[16703] = i[32];
  assign o[16704] = i[32];
  assign o[16705] = i[32];
  assign o[16706] = i[32];
  assign o[16707] = i[32];
  assign o[16708] = i[32];
  assign o[16709] = i[32];
  assign o[16710] = i[32];
  assign o[16711] = i[32];
  assign o[16712] = i[32];
  assign o[16713] = i[32];
  assign o[16714] = i[32];
  assign o[16715] = i[32];
  assign o[16716] = i[32];
  assign o[16717] = i[32];
  assign o[16718] = i[32];
  assign o[16719] = i[32];
  assign o[16720] = i[32];
  assign o[16721] = i[32];
  assign o[16722] = i[32];
  assign o[16723] = i[32];
  assign o[16724] = i[32];
  assign o[16725] = i[32];
  assign o[16726] = i[32];
  assign o[16727] = i[32];
  assign o[16728] = i[32];
  assign o[16729] = i[32];
  assign o[16730] = i[32];
  assign o[16731] = i[32];
  assign o[16732] = i[32];
  assign o[16733] = i[32];
  assign o[16734] = i[32];
  assign o[16735] = i[32];
  assign o[16736] = i[32];
  assign o[16737] = i[32];
  assign o[16738] = i[32];
  assign o[16739] = i[32];
  assign o[16740] = i[32];
  assign o[16741] = i[32];
  assign o[16742] = i[32];
  assign o[16743] = i[32];
  assign o[16744] = i[32];
  assign o[16745] = i[32];
  assign o[16746] = i[32];
  assign o[16747] = i[32];
  assign o[16748] = i[32];
  assign o[16749] = i[32];
  assign o[16750] = i[32];
  assign o[16751] = i[32];
  assign o[16752] = i[32];
  assign o[16753] = i[32];
  assign o[16754] = i[32];
  assign o[16755] = i[32];
  assign o[16756] = i[32];
  assign o[16757] = i[32];
  assign o[16758] = i[32];
  assign o[16759] = i[32];
  assign o[16760] = i[32];
  assign o[16761] = i[32];
  assign o[16762] = i[32];
  assign o[16763] = i[32];
  assign o[16764] = i[32];
  assign o[16765] = i[32];
  assign o[16766] = i[32];
  assign o[16767] = i[32];
  assign o[16768] = i[32];
  assign o[16769] = i[32];
  assign o[16770] = i[32];
  assign o[16771] = i[32];
  assign o[16772] = i[32];
  assign o[16773] = i[32];
  assign o[16774] = i[32];
  assign o[16775] = i[32];
  assign o[16776] = i[32];
  assign o[16777] = i[32];
  assign o[16778] = i[32];
  assign o[16779] = i[32];
  assign o[16780] = i[32];
  assign o[16781] = i[32];
  assign o[16782] = i[32];
  assign o[16783] = i[32];
  assign o[16784] = i[32];
  assign o[16785] = i[32];
  assign o[16786] = i[32];
  assign o[16787] = i[32];
  assign o[16788] = i[32];
  assign o[16789] = i[32];
  assign o[16790] = i[32];
  assign o[16791] = i[32];
  assign o[16792] = i[32];
  assign o[16793] = i[32];
  assign o[16794] = i[32];
  assign o[16795] = i[32];
  assign o[16796] = i[32];
  assign o[16797] = i[32];
  assign o[16798] = i[32];
  assign o[16799] = i[32];
  assign o[16800] = i[32];
  assign o[16801] = i[32];
  assign o[16802] = i[32];
  assign o[16803] = i[32];
  assign o[16804] = i[32];
  assign o[16805] = i[32];
  assign o[16806] = i[32];
  assign o[16807] = i[32];
  assign o[16808] = i[32];
  assign o[16809] = i[32];
  assign o[16810] = i[32];
  assign o[16811] = i[32];
  assign o[16812] = i[32];
  assign o[16813] = i[32];
  assign o[16814] = i[32];
  assign o[16815] = i[32];
  assign o[16816] = i[32];
  assign o[16817] = i[32];
  assign o[16818] = i[32];
  assign o[16819] = i[32];
  assign o[16820] = i[32];
  assign o[16821] = i[32];
  assign o[16822] = i[32];
  assign o[16823] = i[32];
  assign o[16824] = i[32];
  assign o[16825] = i[32];
  assign o[16826] = i[32];
  assign o[16827] = i[32];
  assign o[16828] = i[32];
  assign o[16829] = i[32];
  assign o[16830] = i[32];
  assign o[16831] = i[32];
  assign o[16832] = i[32];
  assign o[16833] = i[32];
  assign o[16834] = i[32];
  assign o[16835] = i[32];
  assign o[16836] = i[32];
  assign o[16837] = i[32];
  assign o[16838] = i[32];
  assign o[16839] = i[32];
  assign o[16840] = i[32];
  assign o[16841] = i[32];
  assign o[16842] = i[32];
  assign o[16843] = i[32];
  assign o[16844] = i[32];
  assign o[16845] = i[32];
  assign o[16846] = i[32];
  assign o[16847] = i[32];
  assign o[16848] = i[32];
  assign o[16849] = i[32];
  assign o[16850] = i[32];
  assign o[16851] = i[32];
  assign o[16852] = i[32];
  assign o[16853] = i[32];
  assign o[16854] = i[32];
  assign o[16855] = i[32];
  assign o[16856] = i[32];
  assign o[16857] = i[32];
  assign o[16858] = i[32];
  assign o[16859] = i[32];
  assign o[16860] = i[32];
  assign o[16861] = i[32];
  assign o[16862] = i[32];
  assign o[16863] = i[32];
  assign o[16864] = i[32];
  assign o[16865] = i[32];
  assign o[16866] = i[32];
  assign o[16867] = i[32];
  assign o[16868] = i[32];
  assign o[16869] = i[32];
  assign o[16870] = i[32];
  assign o[16871] = i[32];
  assign o[16872] = i[32];
  assign o[16873] = i[32];
  assign o[16874] = i[32];
  assign o[16875] = i[32];
  assign o[16876] = i[32];
  assign o[16877] = i[32];
  assign o[16878] = i[32];
  assign o[16879] = i[32];
  assign o[16880] = i[32];
  assign o[16881] = i[32];
  assign o[16882] = i[32];
  assign o[16883] = i[32];
  assign o[16884] = i[32];
  assign o[16885] = i[32];
  assign o[16886] = i[32];
  assign o[16887] = i[32];
  assign o[16888] = i[32];
  assign o[16889] = i[32];
  assign o[16890] = i[32];
  assign o[16891] = i[32];
  assign o[16892] = i[32];
  assign o[16893] = i[32];
  assign o[16894] = i[32];
  assign o[16895] = i[32];
  assign o[15872] = i[31];
  assign o[15873] = i[31];
  assign o[15874] = i[31];
  assign o[15875] = i[31];
  assign o[15876] = i[31];
  assign o[15877] = i[31];
  assign o[15878] = i[31];
  assign o[15879] = i[31];
  assign o[15880] = i[31];
  assign o[15881] = i[31];
  assign o[15882] = i[31];
  assign o[15883] = i[31];
  assign o[15884] = i[31];
  assign o[15885] = i[31];
  assign o[15886] = i[31];
  assign o[15887] = i[31];
  assign o[15888] = i[31];
  assign o[15889] = i[31];
  assign o[15890] = i[31];
  assign o[15891] = i[31];
  assign o[15892] = i[31];
  assign o[15893] = i[31];
  assign o[15894] = i[31];
  assign o[15895] = i[31];
  assign o[15896] = i[31];
  assign o[15897] = i[31];
  assign o[15898] = i[31];
  assign o[15899] = i[31];
  assign o[15900] = i[31];
  assign o[15901] = i[31];
  assign o[15902] = i[31];
  assign o[15903] = i[31];
  assign o[15904] = i[31];
  assign o[15905] = i[31];
  assign o[15906] = i[31];
  assign o[15907] = i[31];
  assign o[15908] = i[31];
  assign o[15909] = i[31];
  assign o[15910] = i[31];
  assign o[15911] = i[31];
  assign o[15912] = i[31];
  assign o[15913] = i[31];
  assign o[15914] = i[31];
  assign o[15915] = i[31];
  assign o[15916] = i[31];
  assign o[15917] = i[31];
  assign o[15918] = i[31];
  assign o[15919] = i[31];
  assign o[15920] = i[31];
  assign o[15921] = i[31];
  assign o[15922] = i[31];
  assign o[15923] = i[31];
  assign o[15924] = i[31];
  assign o[15925] = i[31];
  assign o[15926] = i[31];
  assign o[15927] = i[31];
  assign o[15928] = i[31];
  assign o[15929] = i[31];
  assign o[15930] = i[31];
  assign o[15931] = i[31];
  assign o[15932] = i[31];
  assign o[15933] = i[31];
  assign o[15934] = i[31];
  assign o[15935] = i[31];
  assign o[15936] = i[31];
  assign o[15937] = i[31];
  assign o[15938] = i[31];
  assign o[15939] = i[31];
  assign o[15940] = i[31];
  assign o[15941] = i[31];
  assign o[15942] = i[31];
  assign o[15943] = i[31];
  assign o[15944] = i[31];
  assign o[15945] = i[31];
  assign o[15946] = i[31];
  assign o[15947] = i[31];
  assign o[15948] = i[31];
  assign o[15949] = i[31];
  assign o[15950] = i[31];
  assign o[15951] = i[31];
  assign o[15952] = i[31];
  assign o[15953] = i[31];
  assign o[15954] = i[31];
  assign o[15955] = i[31];
  assign o[15956] = i[31];
  assign o[15957] = i[31];
  assign o[15958] = i[31];
  assign o[15959] = i[31];
  assign o[15960] = i[31];
  assign o[15961] = i[31];
  assign o[15962] = i[31];
  assign o[15963] = i[31];
  assign o[15964] = i[31];
  assign o[15965] = i[31];
  assign o[15966] = i[31];
  assign o[15967] = i[31];
  assign o[15968] = i[31];
  assign o[15969] = i[31];
  assign o[15970] = i[31];
  assign o[15971] = i[31];
  assign o[15972] = i[31];
  assign o[15973] = i[31];
  assign o[15974] = i[31];
  assign o[15975] = i[31];
  assign o[15976] = i[31];
  assign o[15977] = i[31];
  assign o[15978] = i[31];
  assign o[15979] = i[31];
  assign o[15980] = i[31];
  assign o[15981] = i[31];
  assign o[15982] = i[31];
  assign o[15983] = i[31];
  assign o[15984] = i[31];
  assign o[15985] = i[31];
  assign o[15986] = i[31];
  assign o[15987] = i[31];
  assign o[15988] = i[31];
  assign o[15989] = i[31];
  assign o[15990] = i[31];
  assign o[15991] = i[31];
  assign o[15992] = i[31];
  assign o[15993] = i[31];
  assign o[15994] = i[31];
  assign o[15995] = i[31];
  assign o[15996] = i[31];
  assign o[15997] = i[31];
  assign o[15998] = i[31];
  assign o[15999] = i[31];
  assign o[16000] = i[31];
  assign o[16001] = i[31];
  assign o[16002] = i[31];
  assign o[16003] = i[31];
  assign o[16004] = i[31];
  assign o[16005] = i[31];
  assign o[16006] = i[31];
  assign o[16007] = i[31];
  assign o[16008] = i[31];
  assign o[16009] = i[31];
  assign o[16010] = i[31];
  assign o[16011] = i[31];
  assign o[16012] = i[31];
  assign o[16013] = i[31];
  assign o[16014] = i[31];
  assign o[16015] = i[31];
  assign o[16016] = i[31];
  assign o[16017] = i[31];
  assign o[16018] = i[31];
  assign o[16019] = i[31];
  assign o[16020] = i[31];
  assign o[16021] = i[31];
  assign o[16022] = i[31];
  assign o[16023] = i[31];
  assign o[16024] = i[31];
  assign o[16025] = i[31];
  assign o[16026] = i[31];
  assign o[16027] = i[31];
  assign o[16028] = i[31];
  assign o[16029] = i[31];
  assign o[16030] = i[31];
  assign o[16031] = i[31];
  assign o[16032] = i[31];
  assign o[16033] = i[31];
  assign o[16034] = i[31];
  assign o[16035] = i[31];
  assign o[16036] = i[31];
  assign o[16037] = i[31];
  assign o[16038] = i[31];
  assign o[16039] = i[31];
  assign o[16040] = i[31];
  assign o[16041] = i[31];
  assign o[16042] = i[31];
  assign o[16043] = i[31];
  assign o[16044] = i[31];
  assign o[16045] = i[31];
  assign o[16046] = i[31];
  assign o[16047] = i[31];
  assign o[16048] = i[31];
  assign o[16049] = i[31];
  assign o[16050] = i[31];
  assign o[16051] = i[31];
  assign o[16052] = i[31];
  assign o[16053] = i[31];
  assign o[16054] = i[31];
  assign o[16055] = i[31];
  assign o[16056] = i[31];
  assign o[16057] = i[31];
  assign o[16058] = i[31];
  assign o[16059] = i[31];
  assign o[16060] = i[31];
  assign o[16061] = i[31];
  assign o[16062] = i[31];
  assign o[16063] = i[31];
  assign o[16064] = i[31];
  assign o[16065] = i[31];
  assign o[16066] = i[31];
  assign o[16067] = i[31];
  assign o[16068] = i[31];
  assign o[16069] = i[31];
  assign o[16070] = i[31];
  assign o[16071] = i[31];
  assign o[16072] = i[31];
  assign o[16073] = i[31];
  assign o[16074] = i[31];
  assign o[16075] = i[31];
  assign o[16076] = i[31];
  assign o[16077] = i[31];
  assign o[16078] = i[31];
  assign o[16079] = i[31];
  assign o[16080] = i[31];
  assign o[16081] = i[31];
  assign o[16082] = i[31];
  assign o[16083] = i[31];
  assign o[16084] = i[31];
  assign o[16085] = i[31];
  assign o[16086] = i[31];
  assign o[16087] = i[31];
  assign o[16088] = i[31];
  assign o[16089] = i[31];
  assign o[16090] = i[31];
  assign o[16091] = i[31];
  assign o[16092] = i[31];
  assign o[16093] = i[31];
  assign o[16094] = i[31];
  assign o[16095] = i[31];
  assign o[16096] = i[31];
  assign o[16097] = i[31];
  assign o[16098] = i[31];
  assign o[16099] = i[31];
  assign o[16100] = i[31];
  assign o[16101] = i[31];
  assign o[16102] = i[31];
  assign o[16103] = i[31];
  assign o[16104] = i[31];
  assign o[16105] = i[31];
  assign o[16106] = i[31];
  assign o[16107] = i[31];
  assign o[16108] = i[31];
  assign o[16109] = i[31];
  assign o[16110] = i[31];
  assign o[16111] = i[31];
  assign o[16112] = i[31];
  assign o[16113] = i[31];
  assign o[16114] = i[31];
  assign o[16115] = i[31];
  assign o[16116] = i[31];
  assign o[16117] = i[31];
  assign o[16118] = i[31];
  assign o[16119] = i[31];
  assign o[16120] = i[31];
  assign o[16121] = i[31];
  assign o[16122] = i[31];
  assign o[16123] = i[31];
  assign o[16124] = i[31];
  assign o[16125] = i[31];
  assign o[16126] = i[31];
  assign o[16127] = i[31];
  assign o[16128] = i[31];
  assign o[16129] = i[31];
  assign o[16130] = i[31];
  assign o[16131] = i[31];
  assign o[16132] = i[31];
  assign o[16133] = i[31];
  assign o[16134] = i[31];
  assign o[16135] = i[31];
  assign o[16136] = i[31];
  assign o[16137] = i[31];
  assign o[16138] = i[31];
  assign o[16139] = i[31];
  assign o[16140] = i[31];
  assign o[16141] = i[31];
  assign o[16142] = i[31];
  assign o[16143] = i[31];
  assign o[16144] = i[31];
  assign o[16145] = i[31];
  assign o[16146] = i[31];
  assign o[16147] = i[31];
  assign o[16148] = i[31];
  assign o[16149] = i[31];
  assign o[16150] = i[31];
  assign o[16151] = i[31];
  assign o[16152] = i[31];
  assign o[16153] = i[31];
  assign o[16154] = i[31];
  assign o[16155] = i[31];
  assign o[16156] = i[31];
  assign o[16157] = i[31];
  assign o[16158] = i[31];
  assign o[16159] = i[31];
  assign o[16160] = i[31];
  assign o[16161] = i[31];
  assign o[16162] = i[31];
  assign o[16163] = i[31];
  assign o[16164] = i[31];
  assign o[16165] = i[31];
  assign o[16166] = i[31];
  assign o[16167] = i[31];
  assign o[16168] = i[31];
  assign o[16169] = i[31];
  assign o[16170] = i[31];
  assign o[16171] = i[31];
  assign o[16172] = i[31];
  assign o[16173] = i[31];
  assign o[16174] = i[31];
  assign o[16175] = i[31];
  assign o[16176] = i[31];
  assign o[16177] = i[31];
  assign o[16178] = i[31];
  assign o[16179] = i[31];
  assign o[16180] = i[31];
  assign o[16181] = i[31];
  assign o[16182] = i[31];
  assign o[16183] = i[31];
  assign o[16184] = i[31];
  assign o[16185] = i[31];
  assign o[16186] = i[31];
  assign o[16187] = i[31];
  assign o[16188] = i[31];
  assign o[16189] = i[31];
  assign o[16190] = i[31];
  assign o[16191] = i[31];
  assign o[16192] = i[31];
  assign o[16193] = i[31];
  assign o[16194] = i[31];
  assign o[16195] = i[31];
  assign o[16196] = i[31];
  assign o[16197] = i[31];
  assign o[16198] = i[31];
  assign o[16199] = i[31];
  assign o[16200] = i[31];
  assign o[16201] = i[31];
  assign o[16202] = i[31];
  assign o[16203] = i[31];
  assign o[16204] = i[31];
  assign o[16205] = i[31];
  assign o[16206] = i[31];
  assign o[16207] = i[31];
  assign o[16208] = i[31];
  assign o[16209] = i[31];
  assign o[16210] = i[31];
  assign o[16211] = i[31];
  assign o[16212] = i[31];
  assign o[16213] = i[31];
  assign o[16214] = i[31];
  assign o[16215] = i[31];
  assign o[16216] = i[31];
  assign o[16217] = i[31];
  assign o[16218] = i[31];
  assign o[16219] = i[31];
  assign o[16220] = i[31];
  assign o[16221] = i[31];
  assign o[16222] = i[31];
  assign o[16223] = i[31];
  assign o[16224] = i[31];
  assign o[16225] = i[31];
  assign o[16226] = i[31];
  assign o[16227] = i[31];
  assign o[16228] = i[31];
  assign o[16229] = i[31];
  assign o[16230] = i[31];
  assign o[16231] = i[31];
  assign o[16232] = i[31];
  assign o[16233] = i[31];
  assign o[16234] = i[31];
  assign o[16235] = i[31];
  assign o[16236] = i[31];
  assign o[16237] = i[31];
  assign o[16238] = i[31];
  assign o[16239] = i[31];
  assign o[16240] = i[31];
  assign o[16241] = i[31];
  assign o[16242] = i[31];
  assign o[16243] = i[31];
  assign o[16244] = i[31];
  assign o[16245] = i[31];
  assign o[16246] = i[31];
  assign o[16247] = i[31];
  assign o[16248] = i[31];
  assign o[16249] = i[31];
  assign o[16250] = i[31];
  assign o[16251] = i[31];
  assign o[16252] = i[31];
  assign o[16253] = i[31];
  assign o[16254] = i[31];
  assign o[16255] = i[31];
  assign o[16256] = i[31];
  assign o[16257] = i[31];
  assign o[16258] = i[31];
  assign o[16259] = i[31];
  assign o[16260] = i[31];
  assign o[16261] = i[31];
  assign o[16262] = i[31];
  assign o[16263] = i[31];
  assign o[16264] = i[31];
  assign o[16265] = i[31];
  assign o[16266] = i[31];
  assign o[16267] = i[31];
  assign o[16268] = i[31];
  assign o[16269] = i[31];
  assign o[16270] = i[31];
  assign o[16271] = i[31];
  assign o[16272] = i[31];
  assign o[16273] = i[31];
  assign o[16274] = i[31];
  assign o[16275] = i[31];
  assign o[16276] = i[31];
  assign o[16277] = i[31];
  assign o[16278] = i[31];
  assign o[16279] = i[31];
  assign o[16280] = i[31];
  assign o[16281] = i[31];
  assign o[16282] = i[31];
  assign o[16283] = i[31];
  assign o[16284] = i[31];
  assign o[16285] = i[31];
  assign o[16286] = i[31];
  assign o[16287] = i[31];
  assign o[16288] = i[31];
  assign o[16289] = i[31];
  assign o[16290] = i[31];
  assign o[16291] = i[31];
  assign o[16292] = i[31];
  assign o[16293] = i[31];
  assign o[16294] = i[31];
  assign o[16295] = i[31];
  assign o[16296] = i[31];
  assign o[16297] = i[31];
  assign o[16298] = i[31];
  assign o[16299] = i[31];
  assign o[16300] = i[31];
  assign o[16301] = i[31];
  assign o[16302] = i[31];
  assign o[16303] = i[31];
  assign o[16304] = i[31];
  assign o[16305] = i[31];
  assign o[16306] = i[31];
  assign o[16307] = i[31];
  assign o[16308] = i[31];
  assign o[16309] = i[31];
  assign o[16310] = i[31];
  assign o[16311] = i[31];
  assign o[16312] = i[31];
  assign o[16313] = i[31];
  assign o[16314] = i[31];
  assign o[16315] = i[31];
  assign o[16316] = i[31];
  assign o[16317] = i[31];
  assign o[16318] = i[31];
  assign o[16319] = i[31];
  assign o[16320] = i[31];
  assign o[16321] = i[31];
  assign o[16322] = i[31];
  assign o[16323] = i[31];
  assign o[16324] = i[31];
  assign o[16325] = i[31];
  assign o[16326] = i[31];
  assign o[16327] = i[31];
  assign o[16328] = i[31];
  assign o[16329] = i[31];
  assign o[16330] = i[31];
  assign o[16331] = i[31];
  assign o[16332] = i[31];
  assign o[16333] = i[31];
  assign o[16334] = i[31];
  assign o[16335] = i[31];
  assign o[16336] = i[31];
  assign o[16337] = i[31];
  assign o[16338] = i[31];
  assign o[16339] = i[31];
  assign o[16340] = i[31];
  assign o[16341] = i[31];
  assign o[16342] = i[31];
  assign o[16343] = i[31];
  assign o[16344] = i[31];
  assign o[16345] = i[31];
  assign o[16346] = i[31];
  assign o[16347] = i[31];
  assign o[16348] = i[31];
  assign o[16349] = i[31];
  assign o[16350] = i[31];
  assign o[16351] = i[31];
  assign o[16352] = i[31];
  assign o[16353] = i[31];
  assign o[16354] = i[31];
  assign o[16355] = i[31];
  assign o[16356] = i[31];
  assign o[16357] = i[31];
  assign o[16358] = i[31];
  assign o[16359] = i[31];
  assign o[16360] = i[31];
  assign o[16361] = i[31];
  assign o[16362] = i[31];
  assign o[16363] = i[31];
  assign o[16364] = i[31];
  assign o[16365] = i[31];
  assign o[16366] = i[31];
  assign o[16367] = i[31];
  assign o[16368] = i[31];
  assign o[16369] = i[31];
  assign o[16370] = i[31];
  assign o[16371] = i[31];
  assign o[16372] = i[31];
  assign o[16373] = i[31];
  assign o[16374] = i[31];
  assign o[16375] = i[31];
  assign o[16376] = i[31];
  assign o[16377] = i[31];
  assign o[16378] = i[31];
  assign o[16379] = i[31];
  assign o[16380] = i[31];
  assign o[16381] = i[31];
  assign o[16382] = i[31];
  assign o[16383] = i[31];
  assign o[15360] = i[30];
  assign o[15361] = i[30];
  assign o[15362] = i[30];
  assign o[15363] = i[30];
  assign o[15364] = i[30];
  assign o[15365] = i[30];
  assign o[15366] = i[30];
  assign o[15367] = i[30];
  assign o[15368] = i[30];
  assign o[15369] = i[30];
  assign o[15370] = i[30];
  assign o[15371] = i[30];
  assign o[15372] = i[30];
  assign o[15373] = i[30];
  assign o[15374] = i[30];
  assign o[15375] = i[30];
  assign o[15376] = i[30];
  assign o[15377] = i[30];
  assign o[15378] = i[30];
  assign o[15379] = i[30];
  assign o[15380] = i[30];
  assign o[15381] = i[30];
  assign o[15382] = i[30];
  assign o[15383] = i[30];
  assign o[15384] = i[30];
  assign o[15385] = i[30];
  assign o[15386] = i[30];
  assign o[15387] = i[30];
  assign o[15388] = i[30];
  assign o[15389] = i[30];
  assign o[15390] = i[30];
  assign o[15391] = i[30];
  assign o[15392] = i[30];
  assign o[15393] = i[30];
  assign o[15394] = i[30];
  assign o[15395] = i[30];
  assign o[15396] = i[30];
  assign o[15397] = i[30];
  assign o[15398] = i[30];
  assign o[15399] = i[30];
  assign o[15400] = i[30];
  assign o[15401] = i[30];
  assign o[15402] = i[30];
  assign o[15403] = i[30];
  assign o[15404] = i[30];
  assign o[15405] = i[30];
  assign o[15406] = i[30];
  assign o[15407] = i[30];
  assign o[15408] = i[30];
  assign o[15409] = i[30];
  assign o[15410] = i[30];
  assign o[15411] = i[30];
  assign o[15412] = i[30];
  assign o[15413] = i[30];
  assign o[15414] = i[30];
  assign o[15415] = i[30];
  assign o[15416] = i[30];
  assign o[15417] = i[30];
  assign o[15418] = i[30];
  assign o[15419] = i[30];
  assign o[15420] = i[30];
  assign o[15421] = i[30];
  assign o[15422] = i[30];
  assign o[15423] = i[30];
  assign o[15424] = i[30];
  assign o[15425] = i[30];
  assign o[15426] = i[30];
  assign o[15427] = i[30];
  assign o[15428] = i[30];
  assign o[15429] = i[30];
  assign o[15430] = i[30];
  assign o[15431] = i[30];
  assign o[15432] = i[30];
  assign o[15433] = i[30];
  assign o[15434] = i[30];
  assign o[15435] = i[30];
  assign o[15436] = i[30];
  assign o[15437] = i[30];
  assign o[15438] = i[30];
  assign o[15439] = i[30];
  assign o[15440] = i[30];
  assign o[15441] = i[30];
  assign o[15442] = i[30];
  assign o[15443] = i[30];
  assign o[15444] = i[30];
  assign o[15445] = i[30];
  assign o[15446] = i[30];
  assign o[15447] = i[30];
  assign o[15448] = i[30];
  assign o[15449] = i[30];
  assign o[15450] = i[30];
  assign o[15451] = i[30];
  assign o[15452] = i[30];
  assign o[15453] = i[30];
  assign o[15454] = i[30];
  assign o[15455] = i[30];
  assign o[15456] = i[30];
  assign o[15457] = i[30];
  assign o[15458] = i[30];
  assign o[15459] = i[30];
  assign o[15460] = i[30];
  assign o[15461] = i[30];
  assign o[15462] = i[30];
  assign o[15463] = i[30];
  assign o[15464] = i[30];
  assign o[15465] = i[30];
  assign o[15466] = i[30];
  assign o[15467] = i[30];
  assign o[15468] = i[30];
  assign o[15469] = i[30];
  assign o[15470] = i[30];
  assign o[15471] = i[30];
  assign o[15472] = i[30];
  assign o[15473] = i[30];
  assign o[15474] = i[30];
  assign o[15475] = i[30];
  assign o[15476] = i[30];
  assign o[15477] = i[30];
  assign o[15478] = i[30];
  assign o[15479] = i[30];
  assign o[15480] = i[30];
  assign o[15481] = i[30];
  assign o[15482] = i[30];
  assign o[15483] = i[30];
  assign o[15484] = i[30];
  assign o[15485] = i[30];
  assign o[15486] = i[30];
  assign o[15487] = i[30];
  assign o[15488] = i[30];
  assign o[15489] = i[30];
  assign o[15490] = i[30];
  assign o[15491] = i[30];
  assign o[15492] = i[30];
  assign o[15493] = i[30];
  assign o[15494] = i[30];
  assign o[15495] = i[30];
  assign o[15496] = i[30];
  assign o[15497] = i[30];
  assign o[15498] = i[30];
  assign o[15499] = i[30];
  assign o[15500] = i[30];
  assign o[15501] = i[30];
  assign o[15502] = i[30];
  assign o[15503] = i[30];
  assign o[15504] = i[30];
  assign o[15505] = i[30];
  assign o[15506] = i[30];
  assign o[15507] = i[30];
  assign o[15508] = i[30];
  assign o[15509] = i[30];
  assign o[15510] = i[30];
  assign o[15511] = i[30];
  assign o[15512] = i[30];
  assign o[15513] = i[30];
  assign o[15514] = i[30];
  assign o[15515] = i[30];
  assign o[15516] = i[30];
  assign o[15517] = i[30];
  assign o[15518] = i[30];
  assign o[15519] = i[30];
  assign o[15520] = i[30];
  assign o[15521] = i[30];
  assign o[15522] = i[30];
  assign o[15523] = i[30];
  assign o[15524] = i[30];
  assign o[15525] = i[30];
  assign o[15526] = i[30];
  assign o[15527] = i[30];
  assign o[15528] = i[30];
  assign o[15529] = i[30];
  assign o[15530] = i[30];
  assign o[15531] = i[30];
  assign o[15532] = i[30];
  assign o[15533] = i[30];
  assign o[15534] = i[30];
  assign o[15535] = i[30];
  assign o[15536] = i[30];
  assign o[15537] = i[30];
  assign o[15538] = i[30];
  assign o[15539] = i[30];
  assign o[15540] = i[30];
  assign o[15541] = i[30];
  assign o[15542] = i[30];
  assign o[15543] = i[30];
  assign o[15544] = i[30];
  assign o[15545] = i[30];
  assign o[15546] = i[30];
  assign o[15547] = i[30];
  assign o[15548] = i[30];
  assign o[15549] = i[30];
  assign o[15550] = i[30];
  assign o[15551] = i[30];
  assign o[15552] = i[30];
  assign o[15553] = i[30];
  assign o[15554] = i[30];
  assign o[15555] = i[30];
  assign o[15556] = i[30];
  assign o[15557] = i[30];
  assign o[15558] = i[30];
  assign o[15559] = i[30];
  assign o[15560] = i[30];
  assign o[15561] = i[30];
  assign o[15562] = i[30];
  assign o[15563] = i[30];
  assign o[15564] = i[30];
  assign o[15565] = i[30];
  assign o[15566] = i[30];
  assign o[15567] = i[30];
  assign o[15568] = i[30];
  assign o[15569] = i[30];
  assign o[15570] = i[30];
  assign o[15571] = i[30];
  assign o[15572] = i[30];
  assign o[15573] = i[30];
  assign o[15574] = i[30];
  assign o[15575] = i[30];
  assign o[15576] = i[30];
  assign o[15577] = i[30];
  assign o[15578] = i[30];
  assign o[15579] = i[30];
  assign o[15580] = i[30];
  assign o[15581] = i[30];
  assign o[15582] = i[30];
  assign o[15583] = i[30];
  assign o[15584] = i[30];
  assign o[15585] = i[30];
  assign o[15586] = i[30];
  assign o[15587] = i[30];
  assign o[15588] = i[30];
  assign o[15589] = i[30];
  assign o[15590] = i[30];
  assign o[15591] = i[30];
  assign o[15592] = i[30];
  assign o[15593] = i[30];
  assign o[15594] = i[30];
  assign o[15595] = i[30];
  assign o[15596] = i[30];
  assign o[15597] = i[30];
  assign o[15598] = i[30];
  assign o[15599] = i[30];
  assign o[15600] = i[30];
  assign o[15601] = i[30];
  assign o[15602] = i[30];
  assign o[15603] = i[30];
  assign o[15604] = i[30];
  assign o[15605] = i[30];
  assign o[15606] = i[30];
  assign o[15607] = i[30];
  assign o[15608] = i[30];
  assign o[15609] = i[30];
  assign o[15610] = i[30];
  assign o[15611] = i[30];
  assign o[15612] = i[30];
  assign o[15613] = i[30];
  assign o[15614] = i[30];
  assign o[15615] = i[30];
  assign o[15616] = i[30];
  assign o[15617] = i[30];
  assign o[15618] = i[30];
  assign o[15619] = i[30];
  assign o[15620] = i[30];
  assign o[15621] = i[30];
  assign o[15622] = i[30];
  assign o[15623] = i[30];
  assign o[15624] = i[30];
  assign o[15625] = i[30];
  assign o[15626] = i[30];
  assign o[15627] = i[30];
  assign o[15628] = i[30];
  assign o[15629] = i[30];
  assign o[15630] = i[30];
  assign o[15631] = i[30];
  assign o[15632] = i[30];
  assign o[15633] = i[30];
  assign o[15634] = i[30];
  assign o[15635] = i[30];
  assign o[15636] = i[30];
  assign o[15637] = i[30];
  assign o[15638] = i[30];
  assign o[15639] = i[30];
  assign o[15640] = i[30];
  assign o[15641] = i[30];
  assign o[15642] = i[30];
  assign o[15643] = i[30];
  assign o[15644] = i[30];
  assign o[15645] = i[30];
  assign o[15646] = i[30];
  assign o[15647] = i[30];
  assign o[15648] = i[30];
  assign o[15649] = i[30];
  assign o[15650] = i[30];
  assign o[15651] = i[30];
  assign o[15652] = i[30];
  assign o[15653] = i[30];
  assign o[15654] = i[30];
  assign o[15655] = i[30];
  assign o[15656] = i[30];
  assign o[15657] = i[30];
  assign o[15658] = i[30];
  assign o[15659] = i[30];
  assign o[15660] = i[30];
  assign o[15661] = i[30];
  assign o[15662] = i[30];
  assign o[15663] = i[30];
  assign o[15664] = i[30];
  assign o[15665] = i[30];
  assign o[15666] = i[30];
  assign o[15667] = i[30];
  assign o[15668] = i[30];
  assign o[15669] = i[30];
  assign o[15670] = i[30];
  assign o[15671] = i[30];
  assign o[15672] = i[30];
  assign o[15673] = i[30];
  assign o[15674] = i[30];
  assign o[15675] = i[30];
  assign o[15676] = i[30];
  assign o[15677] = i[30];
  assign o[15678] = i[30];
  assign o[15679] = i[30];
  assign o[15680] = i[30];
  assign o[15681] = i[30];
  assign o[15682] = i[30];
  assign o[15683] = i[30];
  assign o[15684] = i[30];
  assign o[15685] = i[30];
  assign o[15686] = i[30];
  assign o[15687] = i[30];
  assign o[15688] = i[30];
  assign o[15689] = i[30];
  assign o[15690] = i[30];
  assign o[15691] = i[30];
  assign o[15692] = i[30];
  assign o[15693] = i[30];
  assign o[15694] = i[30];
  assign o[15695] = i[30];
  assign o[15696] = i[30];
  assign o[15697] = i[30];
  assign o[15698] = i[30];
  assign o[15699] = i[30];
  assign o[15700] = i[30];
  assign o[15701] = i[30];
  assign o[15702] = i[30];
  assign o[15703] = i[30];
  assign o[15704] = i[30];
  assign o[15705] = i[30];
  assign o[15706] = i[30];
  assign o[15707] = i[30];
  assign o[15708] = i[30];
  assign o[15709] = i[30];
  assign o[15710] = i[30];
  assign o[15711] = i[30];
  assign o[15712] = i[30];
  assign o[15713] = i[30];
  assign o[15714] = i[30];
  assign o[15715] = i[30];
  assign o[15716] = i[30];
  assign o[15717] = i[30];
  assign o[15718] = i[30];
  assign o[15719] = i[30];
  assign o[15720] = i[30];
  assign o[15721] = i[30];
  assign o[15722] = i[30];
  assign o[15723] = i[30];
  assign o[15724] = i[30];
  assign o[15725] = i[30];
  assign o[15726] = i[30];
  assign o[15727] = i[30];
  assign o[15728] = i[30];
  assign o[15729] = i[30];
  assign o[15730] = i[30];
  assign o[15731] = i[30];
  assign o[15732] = i[30];
  assign o[15733] = i[30];
  assign o[15734] = i[30];
  assign o[15735] = i[30];
  assign o[15736] = i[30];
  assign o[15737] = i[30];
  assign o[15738] = i[30];
  assign o[15739] = i[30];
  assign o[15740] = i[30];
  assign o[15741] = i[30];
  assign o[15742] = i[30];
  assign o[15743] = i[30];
  assign o[15744] = i[30];
  assign o[15745] = i[30];
  assign o[15746] = i[30];
  assign o[15747] = i[30];
  assign o[15748] = i[30];
  assign o[15749] = i[30];
  assign o[15750] = i[30];
  assign o[15751] = i[30];
  assign o[15752] = i[30];
  assign o[15753] = i[30];
  assign o[15754] = i[30];
  assign o[15755] = i[30];
  assign o[15756] = i[30];
  assign o[15757] = i[30];
  assign o[15758] = i[30];
  assign o[15759] = i[30];
  assign o[15760] = i[30];
  assign o[15761] = i[30];
  assign o[15762] = i[30];
  assign o[15763] = i[30];
  assign o[15764] = i[30];
  assign o[15765] = i[30];
  assign o[15766] = i[30];
  assign o[15767] = i[30];
  assign o[15768] = i[30];
  assign o[15769] = i[30];
  assign o[15770] = i[30];
  assign o[15771] = i[30];
  assign o[15772] = i[30];
  assign o[15773] = i[30];
  assign o[15774] = i[30];
  assign o[15775] = i[30];
  assign o[15776] = i[30];
  assign o[15777] = i[30];
  assign o[15778] = i[30];
  assign o[15779] = i[30];
  assign o[15780] = i[30];
  assign o[15781] = i[30];
  assign o[15782] = i[30];
  assign o[15783] = i[30];
  assign o[15784] = i[30];
  assign o[15785] = i[30];
  assign o[15786] = i[30];
  assign o[15787] = i[30];
  assign o[15788] = i[30];
  assign o[15789] = i[30];
  assign o[15790] = i[30];
  assign o[15791] = i[30];
  assign o[15792] = i[30];
  assign o[15793] = i[30];
  assign o[15794] = i[30];
  assign o[15795] = i[30];
  assign o[15796] = i[30];
  assign o[15797] = i[30];
  assign o[15798] = i[30];
  assign o[15799] = i[30];
  assign o[15800] = i[30];
  assign o[15801] = i[30];
  assign o[15802] = i[30];
  assign o[15803] = i[30];
  assign o[15804] = i[30];
  assign o[15805] = i[30];
  assign o[15806] = i[30];
  assign o[15807] = i[30];
  assign o[15808] = i[30];
  assign o[15809] = i[30];
  assign o[15810] = i[30];
  assign o[15811] = i[30];
  assign o[15812] = i[30];
  assign o[15813] = i[30];
  assign o[15814] = i[30];
  assign o[15815] = i[30];
  assign o[15816] = i[30];
  assign o[15817] = i[30];
  assign o[15818] = i[30];
  assign o[15819] = i[30];
  assign o[15820] = i[30];
  assign o[15821] = i[30];
  assign o[15822] = i[30];
  assign o[15823] = i[30];
  assign o[15824] = i[30];
  assign o[15825] = i[30];
  assign o[15826] = i[30];
  assign o[15827] = i[30];
  assign o[15828] = i[30];
  assign o[15829] = i[30];
  assign o[15830] = i[30];
  assign o[15831] = i[30];
  assign o[15832] = i[30];
  assign o[15833] = i[30];
  assign o[15834] = i[30];
  assign o[15835] = i[30];
  assign o[15836] = i[30];
  assign o[15837] = i[30];
  assign o[15838] = i[30];
  assign o[15839] = i[30];
  assign o[15840] = i[30];
  assign o[15841] = i[30];
  assign o[15842] = i[30];
  assign o[15843] = i[30];
  assign o[15844] = i[30];
  assign o[15845] = i[30];
  assign o[15846] = i[30];
  assign o[15847] = i[30];
  assign o[15848] = i[30];
  assign o[15849] = i[30];
  assign o[15850] = i[30];
  assign o[15851] = i[30];
  assign o[15852] = i[30];
  assign o[15853] = i[30];
  assign o[15854] = i[30];
  assign o[15855] = i[30];
  assign o[15856] = i[30];
  assign o[15857] = i[30];
  assign o[15858] = i[30];
  assign o[15859] = i[30];
  assign o[15860] = i[30];
  assign o[15861] = i[30];
  assign o[15862] = i[30];
  assign o[15863] = i[30];
  assign o[15864] = i[30];
  assign o[15865] = i[30];
  assign o[15866] = i[30];
  assign o[15867] = i[30];
  assign o[15868] = i[30];
  assign o[15869] = i[30];
  assign o[15870] = i[30];
  assign o[15871] = i[30];
  assign o[14848] = i[29];
  assign o[14849] = i[29];
  assign o[14850] = i[29];
  assign o[14851] = i[29];
  assign o[14852] = i[29];
  assign o[14853] = i[29];
  assign o[14854] = i[29];
  assign o[14855] = i[29];
  assign o[14856] = i[29];
  assign o[14857] = i[29];
  assign o[14858] = i[29];
  assign o[14859] = i[29];
  assign o[14860] = i[29];
  assign o[14861] = i[29];
  assign o[14862] = i[29];
  assign o[14863] = i[29];
  assign o[14864] = i[29];
  assign o[14865] = i[29];
  assign o[14866] = i[29];
  assign o[14867] = i[29];
  assign o[14868] = i[29];
  assign o[14869] = i[29];
  assign o[14870] = i[29];
  assign o[14871] = i[29];
  assign o[14872] = i[29];
  assign o[14873] = i[29];
  assign o[14874] = i[29];
  assign o[14875] = i[29];
  assign o[14876] = i[29];
  assign o[14877] = i[29];
  assign o[14878] = i[29];
  assign o[14879] = i[29];
  assign o[14880] = i[29];
  assign o[14881] = i[29];
  assign o[14882] = i[29];
  assign o[14883] = i[29];
  assign o[14884] = i[29];
  assign o[14885] = i[29];
  assign o[14886] = i[29];
  assign o[14887] = i[29];
  assign o[14888] = i[29];
  assign o[14889] = i[29];
  assign o[14890] = i[29];
  assign o[14891] = i[29];
  assign o[14892] = i[29];
  assign o[14893] = i[29];
  assign o[14894] = i[29];
  assign o[14895] = i[29];
  assign o[14896] = i[29];
  assign o[14897] = i[29];
  assign o[14898] = i[29];
  assign o[14899] = i[29];
  assign o[14900] = i[29];
  assign o[14901] = i[29];
  assign o[14902] = i[29];
  assign o[14903] = i[29];
  assign o[14904] = i[29];
  assign o[14905] = i[29];
  assign o[14906] = i[29];
  assign o[14907] = i[29];
  assign o[14908] = i[29];
  assign o[14909] = i[29];
  assign o[14910] = i[29];
  assign o[14911] = i[29];
  assign o[14912] = i[29];
  assign o[14913] = i[29];
  assign o[14914] = i[29];
  assign o[14915] = i[29];
  assign o[14916] = i[29];
  assign o[14917] = i[29];
  assign o[14918] = i[29];
  assign o[14919] = i[29];
  assign o[14920] = i[29];
  assign o[14921] = i[29];
  assign o[14922] = i[29];
  assign o[14923] = i[29];
  assign o[14924] = i[29];
  assign o[14925] = i[29];
  assign o[14926] = i[29];
  assign o[14927] = i[29];
  assign o[14928] = i[29];
  assign o[14929] = i[29];
  assign o[14930] = i[29];
  assign o[14931] = i[29];
  assign o[14932] = i[29];
  assign o[14933] = i[29];
  assign o[14934] = i[29];
  assign o[14935] = i[29];
  assign o[14936] = i[29];
  assign o[14937] = i[29];
  assign o[14938] = i[29];
  assign o[14939] = i[29];
  assign o[14940] = i[29];
  assign o[14941] = i[29];
  assign o[14942] = i[29];
  assign o[14943] = i[29];
  assign o[14944] = i[29];
  assign o[14945] = i[29];
  assign o[14946] = i[29];
  assign o[14947] = i[29];
  assign o[14948] = i[29];
  assign o[14949] = i[29];
  assign o[14950] = i[29];
  assign o[14951] = i[29];
  assign o[14952] = i[29];
  assign o[14953] = i[29];
  assign o[14954] = i[29];
  assign o[14955] = i[29];
  assign o[14956] = i[29];
  assign o[14957] = i[29];
  assign o[14958] = i[29];
  assign o[14959] = i[29];
  assign o[14960] = i[29];
  assign o[14961] = i[29];
  assign o[14962] = i[29];
  assign o[14963] = i[29];
  assign o[14964] = i[29];
  assign o[14965] = i[29];
  assign o[14966] = i[29];
  assign o[14967] = i[29];
  assign o[14968] = i[29];
  assign o[14969] = i[29];
  assign o[14970] = i[29];
  assign o[14971] = i[29];
  assign o[14972] = i[29];
  assign o[14973] = i[29];
  assign o[14974] = i[29];
  assign o[14975] = i[29];
  assign o[14976] = i[29];
  assign o[14977] = i[29];
  assign o[14978] = i[29];
  assign o[14979] = i[29];
  assign o[14980] = i[29];
  assign o[14981] = i[29];
  assign o[14982] = i[29];
  assign o[14983] = i[29];
  assign o[14984] = i[29];
  assign o[14985] = i[29];
  assign o[14986] = i[29];
  assign o[14987] = i[29];
  assign o[14988] = i[29];
  assign o[14989] = i[29];
  assign o[14990] = i[29];
  assign o[14991] = i[29];
  assign o[14992] = i[29];
  assign o[14993] = i[29];
  assign o[14994] = i[29];
  assign o[14995] = i[29];
  assign o[14996] = i[29];
  assign o[14997] = i[29];
  assign o[14998] = i[29];
  assign o[14999] = i[29];
  assign o[15000] = i[29];
  assign o[15001] = i[29];
  assign o[15002] = i[29];
  assign o[15003] = i[29];
  assign o[15004] = i[29];
  assign o[15005] = i[29];
  assign o[15006] = i[29];
  assign o[15007] = i[29];
  assign o[15008] = i[29];
  assign o[15009] = i[29];
  assign o[15010] = i[29];
  assign o[15011] = i[29];
  assign o[15012] = i[29];
  assign o[15013] = i[29];
  assign o[15014] = i[29];
  assign o[15015] = i[29];
  assign o[15016] = i[29];
  assign o[15017] = i[29];
  assign o[15018] = i[29];
  assign o[15019] = i[29];
  assign o[15020] = i[29];
  assign o[15021] = i[29];
  assign o[15022] = i[29];
  assign o[15023] = i[29];
  assign o[15024] = i[29];
  assign o[15025] = i[29];
  assign o[15026] = i[29];
  assign o[15027] = i[29];
  assign o[15028] = i[29];
  assign o[15029] = i[29];
  assign o[15030] = i[29];
  assign o[15031] = i[29];
  assign o[15032] = i[29];
  assign o[15033] = i[29];
  assign o[15034] = i[29];
  assign o[15035] = i[29];
  assign o[15036] = i[29];
  assign o[15037] = i[29];
  assign o[15038] = i[29];
  assign o[15039] = i[29];
  assign o[15040] = i[29];
  assign o[15041] = i[29];
  assign o[15042] = i[29];
  assign o[15043] = i[29];
  assign o[15044] = i[29];
  assign o[15045] = i[29];
  assign o[15046] = i[29];
  assign o[15047] = i[29];
  assign o[15048] = i[29];
  assign o[15049] = i[29];
  assign o[15050] = i[29];
  assign o[15051] = i[29];
  assign o[15052] = i[29];
  assign o[15053] = i[29];
  assign o[15054] = i[29];
  assign o[15055] = i[29];
  assign o[15056] = i[29];
  assign o[15057] = i[29];
  assign o[15058] = i[29];
  assign o[15059] = i[29];
  assign o[15060] = i[29];
  assign o[15061] = i[29];
  assign o[15062] = i[29];
  assign o[15063] = i[29];
  assign o[15064] = i[29];
  assign o[15065] = i[29];
  assign o[15066] = i[29];
  assign o[15067] = i[29];
  assign o[15068] = i[29];
  assign o[15069] = i[29];
  assign o[15070] = i[29];
  assign o[15071] = i[29];
  assign o[15072] = i[29];
  assign o[15073] = i[29];
  assign o[15074] = i[29];
  assign o[15075] = i[29];
  assign o[15076] = i[29];
  assign o[15077] = i[29];
  assign o[15078] = i[29];
  assign o[15079] = i[29];
  assign o[15080] = i[29];
  assign o[15081] = i[29];
  assign o[15082] = i[29];
  assign o[15083] = i[29];
  assign o[15084] = i[29];
  assign o[15085] = i[29];
  assign o[15086] = i[29];
  assign o[15087] = i[29];
  assign o[15088] = i[29];
  assign o[15089] = i[29];
  assign o[15090] = i[29];
  assign o[15091] = i[29];
  assign o[15092] = i[29];
  assign o[15093] = i[29];
  assign o[15094] = i[29];
  assign o[15095] = i[29];
  assign o[15096] = i[29];
  assign o[15097] = i[29];
  assign o[15098] = i[29];
  assign o[15099] = i[29];
  assign o[15100] = i[29];
  assign o[15101] = i[29];
  assign o[15102] = i[29];
  assign o[15103] = i[29];
  assign o[15104] = i[29];
  assign o[15105] = i[29];
  assign o[15106] = i[29];
  assign o[15107] = i[29];
  assign o[15108] = i[29];
  assign o[15109] = i[29];
  assign o[15110] = i[29];
  assign o[15111] = i[29];
  assign o[15112] = i[29];
  assign o[15113] = i[29];
  assign o[15114] = i[29];
  assign o[15115] = i[29];
  assign o[15116] = i[29];
  assign o[15117] = i[29];
  assign o[15118] = i[29];
  assign o[15119] = i[29];
  assign o[15120] = i[29];
  assign o[15121] = i[29];
  assign o[15122] = i[29];
  assign o[15123] = i[29];
  assign o[15124] = i[29];
  assign o[15125] = i[29];
  assign o[15126] = i[29];
  assign o[15127] = i[29];
  assign o[15128] = i[29];
  assign o[15129] = i[29];
  assign o[15130] = i[29];
  assign o[15131] = i[29];
  assign o[15132] = i[29];
  assign o[15133] = i[29];
  assign o[15134] = i[29];
  assign o[15135] = i[29];
  assign o[15136] = i[29];
  assign o[15137] = i[29];
  assign o[15138] = i[29];
  assign o[15139] = i[29];
  assign o[15140] = i[29];
  assign o[15141] = i[29];
  assign o[15142] = i[29];
  assign o[15143] = i[29];
  assign o[15144] = i[29];
  assign o[15145] = i[29];
  assign o[15146] = i[29];
  assign o[15147] = i[29];
  assign o[15148] = i[29];
  assign o[15149] = i[29];
  assign o[15150] = i[29];
  assign o[15151] = i[29];
  assign o[15152] = i[29];
  assign o[15153] = i[29];
  assign o[15154] = i[29];
  assign o[15155] = i[29];
  assign o[15156] = i[29];
  assign o[15157] = i[29];
  assign o[15158] = i[29];
  assign o[15159] = i[29];
  assign o[15160] = i[29];
  assign o[15161] = i[29];
  assign o[15162] = i[29];
  assign o[15163] = i[29];
  assign o[15164] = i[29];
  assign o[15165] = i[29];
  assign o[15166] = i[29];
  assign o[15167] = i[29];
  assign o[15168] = i[29];
  assign o[15169] = i[29];
  assign o[15170] = i[29];
  assign o[15171] = i[29];
  assign o[15172] = i[29];
  assign o[15173] = i[29];
  assign o[15174] = i[29];
  assign o[15175] = i[29];
  assign o[15176] = i[29];
  assign o[15177] = i[29];
  assign o[15178] = i[29];
  assign o[15179] = i[29];
  assign o[15180] = i[29];
  assign o[15181] = i[29];
  assign o[15182] = i[29];
  assign o[15183] = i[29];
  assign o[15184] = i[29];
  assign o[15185] = i[29];
  assign o[15186] = i[29];
  assign o[15187] = i[29];
  assign o[15188] = i[29];
  assign o[15189] = i[29];
  assign o[15190] = i[29];
  assign o[15191] = i[29];
  assign o[15192] = i[29];
  assign o[15193] = i[29];
  assign o[15194] = i[29];
  assign o[15195] = i[29];
  assign o[15196] = i[29];
  assign o[15197] = i[29];
  assign o[15198] = i[29];
  assign o[15199] = i[29];
  assign o[15200] = i[29];
  assign o[15201] = i[29];
  assign o[15202] = i[29];
  assign o[15203] = i[29];
  assign o[15204] = i[29];
  assign o[15205] = i[29];
  assign o[15206] = i[29];
  assign o[15207] = i[29];
  assign o[15208] = i[29];
  assign o[15209] = i[29];
  assign o[15210] = i[29];
  assign o[15211] = i[29];
  assign o[15212] = i[29];
  assign o[15213] = i[29];
  assign o[15214] = i[29];
  assign o[15215] = i[29];
  assign o[15216] = i[29];
  assign o[15217] = i[29];
  assign o[15218] = i[29];
  assign o[15219] = i[29];
  assign o[15220] = i[29];
  assign o[15221] = i[29];
  assign o[15222] = i[29];
  assign o[15223] = i[29];
  assign o[15224] = i[29];
  assign o[15225] = i[29];
  assign o[15226] = i[29];
  assign o[15227] = i[29];
  assign o[15228] = i[29];
  assign o[15229] = i[29];
  assign o[15230] = i[29];
  assign o[15231] = i[29];
  assign o[15232] = i[29];
  assign o[15233] = i[29];
  assign o[15234] = i[29];
  assign o[15235] = i[29];
  assign o[15236] = i[29];
  assign o[15237] = i[29];
  assign o[15238] = i[29];
  assign o[15239] = i[29];
  assign o[15240] = i[29];
  assign o[15241] = i[29];
  assign o[15242] = i[29];
  assign o[15243] = i[29];
  assign o[15244] = i[29];
  assign o[15245] = i[29];
  assign o[15246] = i[29];
  assign o[15247] = i[29];
  assign o[15248] = i[29];
  assign o[15249] = i[29];
  assign o[15250] = i[29];
  assign o[15251] = i[29];
  assign o[15252] = i[29];
  assign o[15253] = i[29];
  assign o[15254] = i[29];
  assign o[15255] = i[29];
  assign o[15256] = i[29];
  assign o[15257] = i[29];
  assign o[15258] = i[29];
  assign o[15259] = i[29];
  assign o[15260] = i[29];
  assign o[15261] = i[29];
  assign o[15262] = i[29];
  assign o[15263] = i[29];
  assign o[15264] = i[29];
  assign o[15265] = i[29];
  assign o[15266] = i[29];
  assign o[15267] = i[29];
  assign o[15268] = i[29];
  assign o[15269] = i[29];
  assign o[15270] = i[29];
  assign o[15271] = i[29];
  assign o[15272] = i[29];
  assign o[15273] = i[29];
  assign o[15274] = i[29];
  assign o[15275] = i[29];
  assign o[15276] = i[29];
  assign o[15277] = i[29];
  assign o[15278] = i[29];
  assign o[15279] = i[29];
  assign o[15280] = i[29];
  assign o[15281] = i[29];
  assign o[15282] = i[29];
  assign o[15283] = i[29];
  assign o[15284] = i[29];
  assign o[15285] = i[29];
  assign o[15286] = i[29];
  assign o[15287] = i[29];
  assign o[15288] = i[29];
  assign o[15289] = i[29];
  assign o[15290] = i[29];
  assign o[15291] = i[29];
  assign o[15292] = i[29];
  assign o[15293] = i[29];
  assign o[15294] = i[29];
  assign o[15295] = i[29];
  assign o[15296] = i[29];
  assign o[15297] = i[29];
  assign o[15298] = i[29];
  assign o[15299] = i[29];
  assign o[15300] = i[29];
  assign o[15301] = i[29];
  assign o[15302] = i[29];
  assign o[15303] = i[29];
  assign o[15304] = i[29];
  assign o[15305] = i[29];
  assign o[15306] = i[29];
  assign o[15307] = i[29];
  assign o[15308] = i[29];
  assign o[15309] = i[29];
  assign o[15310] = i[29];
  assign o[15311] = i[29];
  assign o[15312] = i[29];
  assign o[15313] = i[29];
  assign o[15314] = i[29];
  assign o[15315] = i[29];
  assign o[15316] = i[29];
  assign o[15317] = i[29];
  assign o[15318] = i[29];
  assign o[15319] = i[29];
  assign o[15320] = i[29];
  assign o[15321] = i[29];
  assign o[15322] = i[29];
  assign o[15323] = i[29];
  assign o[15324] = i[29];
  assign o[15325] = i[29];
  assign o[15326] = i[29];
  assign o[15327] = i[29];
  assign o[15328] = i[29];
  assign o[15329] = i[29];
  assign o[15330] = i[29];
  assign o[15331] = i[29];
  assign o[15332] = i[29];
  assign o[15333] = i[29];
  assign o[15334] = i[29];
  assign o[15335] = i[29];
  assign o[15336] = i[29];
  assign o[15337] = i[29];
  assign o[15338] = i[29];
  assign o[15339] = i[29];
  assign o[15340] = i[29];
  assign o[15341] = i[29];
  assign o[15342] = i[29];
  assign o[15343] = i[29];
  assign o[15344] = i[29];
  assign o[15345] = i[29];
  assign o[15346] = i[29];
  assign o[15347] = i[29];
  assign o[15348] = i[29];
  assign o[15349] = i[29];
  assign o[15350] = i[29];
  assign o[15351] = i[29];
  assign o[15352] = i[29];
  assign o[15353] = i[29];
  assign o[15354] = i[29];
  assign o[15355] = i[29];
  assign o[15356] = i[29];
  assign o[15357] = i[29];
  assign o[15358] = i[29];
  assign o[15359] = i[29];
  assign o[14336] = i[28];
  assign o[14337] = i[28];
  assign o[14338] = i[28];
  assign o[14339] = i[28];
  assign o[14340] = i[28];
  assign o[14341] = i[28];
  assign o[14342] = i[28];
  assign o[14343] = i[28];
  assign o[14344] = i[28];
  assign o[14345] = i[28];
  assign o[14346] = i[28];
  assign o[14347] = i[28];
  assign o[14348] = i[28];
  assign o[14349] = i[28];
  assign o[14350] = i[28];
  assign o[14351] = i[28];
  assign o[14352] = i[28];
  assign o[14353] = i[28];
  assign o[14354] = i[28];
  assign o[14355] = i[28];
  assign o[14356] = i[28];
  assign o[14357] = i[28];
  assign o[14358] = i[28];
  assign o[14359] = i[28];
  assign o[14360] = i[28];
  assign o[14361] = i[28];
  assign o[14362] = i[28];
  assign o[14363] = i[28];
  assign o[14364] = i[28];
  assign o[14365] = i[28];
  assign o[14366] = i[28];
  assign o[14367] = i[28];
  assign o[14368] = i[28];
  assign o[14369] = i[28];
  assign o[14370] = i[28];
  assign o[14371] = i[28];
  assign o[14372] = i[28];
  assign o[14373] = i[28];
  assign o[14374] = i[28];
  assign o[14375] = i[28];
  assign o[14376] = i[28];
  assign o[14377] = i[28];
  assign o[14378] = i[28];
  assign o[14379] = i[28];
  assign o[14380] = i[28];
  assign o[14381] = i[28];
  assign o[14382] = i[28];
  assign o[14383] = i[28];
  assign o[14384] = i[28];
  assign o[14385] = i[28];
  assign o[14386] = i[28];
  assign o[14387] = i[28];
  assign o[14388] = i[28];
  assign o[14389] = i[28];
  assign o[14390] = i[28];
  assign o[14391] = i[28];
  assign o[14392] = i[28];
  assign o[14393] = i[28];
  assign o[14394] = i[28];
  assign o[14395] = i[28];
  assign o[14396] = i[28];
  assign o[14397] = i[28];
  assign o[14398] = i[28];
  assign o[14399] = i[28];
  assign o[14400] = i[28];
  assign o[14401] = i[28];
  assign o[14402] = i[28];
  assign o[14403] = i[28];
  assign o[14404] = i[28];
  assign o[14405] = i[28];
  assign o[14406] = i[28];
  assign o[14407] = i[28];
  assign o[14408] = i[28];
  assign o[14409] = i[28];
  assign o[14410] = i[28];
  assign o[14411] = i[28];
  assign o[14412] = i[28];
  assign o[14413] = i[28];
  assign o[14414] = i[28];
  assign o[14415] = i[28];
  assign o[14416] = i[28];
  assign o[14417] = i[28];
  assign o[14418] = i[28];
  assign o[14419] = i[28];
  assign o[14420] = i[28];
  assign o[14421] = i[28];
  assign o[14422] = i[28];
  assign o[14423] = i[28];
  assign o[14424] = i[28];
  assign o[14425] = i[28];
  assign o[14426] = i[28];
  assign o[14427] = i[28];
  assign o[14428] = i[28];
  assign o[14429] = i[28];
  assign o[14430] = i[28];
  assign o[14431] = i[28];
  assign o[14432] = i[28];
  assign o[14433] = i[28];
  assign o[14434] = i[28];
  assign o[14435] = i[28];
  assign o[14436] = i[28];
  assign o[14437] = i[28];
  assign o[14438] = i[28];
  assign o[14439] = i[28];
  assign o[14440] = i[28];
  assign o[14441] = i[28];
  assign o[14442] = i[28];
  assign o[14443] = i[28];
  assign o[14444] = i[28];
  assign o[14445] = i[28];
  assign o[14446] = i[28];
  assign o[14447] = i[28];
  assign o[14448] = i[28];
  assign o[14449] = i[28];
  assign o[14450] = i[28];
  assign o[14451] = i[28];
  assign o[14452] = i[28];
  assign o[14453] = i[28];
  assign o[14454] = i[28];
  assign o[14455] = i[28];
  assign o[14456] = i[28];
  assign o[14457] = i[28];
  assign o[14458] = i[28];
  assign o[14459] = i[28];
  assign o[14460] = i[28];
  assign o[14461] = i[28];
  assign o[14462] = i[28];
  assign o[14463] = i[28];
  assign o[14464] = i[28];
  assign o[14465] = i[28];
  assign o[14466] = i[28];
  assign o[14467] = i[28];
  assign o[14468] = i[28];
  assign o[14469] = i[28];
  assign o[14470] = i[28];
  assign o[14471] = i[28];
  assign o[14472] = i[28];
  assign o[14473] = i[28];
  assign o[14474] = i[28];
  assign o[14475] = i[28];
  assign o[14476] = i[28];
  assign o[14477] = i[28];
  assign o[14478] = i[28];
  assign o[14479] = i[28];
  assign o[14480] = i[28];
  assign o[14481] = i[28];
  assign o[14482] = i[28];
  assign o[14483] = i[28];
  assign o[14484] = i[28];
  assign o[14485] = i[28];
  assign o[14486] = i[28];
  assign o[14487] = i[28];
  assign o[14488] = i[28];
  assign o[14489] = i[28];
  assign o[14490] = i[28];
  assign o[14491] = i[28];
  assign o[14492] = i[28];
  assign o[14493] = i[28];
  assign o[14494] = i[28];
  assign o[14495] = i[28];
  assign o[14496] = i[28];
  assign o[14497] = i[28];
  assign o[14498] = i[28];
  assign o[14499] = i[28];
  assign o[14500] = i[28];
  assign o[14501] = i[28];
  assign o[14502] = i[28];
  assign o[14503] = i[28];
  assign o[14504] = i[28];
  assign o[14505] = i[28];
  assign o[14506] = i[28];
  assign o[14507] = i[28];
  assign o[14508] = i[28];
  assign o[14509] = i[28];
  assign o[14510] = i[28];
  assign o[14511] = i[28];
  assign o[14512] = i[28];
  assign o[14513] = i[28];
  assign o[14514] = i[28];
  assign o[14515] = i[28];
  assign o[14516] = i[28];
  assign o[14517] = i[28];
  assign o[14518] = i[28];
  assign o[14519] = i[28];
  assign o[14520] = i[28];
  assign o[14521] = i[28];
  assign o[14522] = i[28];
  assign o[14523] = i[28];
  assign o[14524] = i[28];
  assign o[14525] = i[28];
  assign o[14526] = i[28];
  assign o[14527] = i[28];
  assign o[14528] = i[28];
  assign o[14529] = i[28];
  assign o[14530] = i[28];
  assign o[14531] = i[28];
  assign o[14532] = i[28];
  assign o[14533] = i[28];
  assign o[14534] = i[28];
  assign o[14535] = i[28];
  assign o[14536] = i[28];
  assign o[14537] = i[28];
  assign o[14538] = i[28];
  assign o[14539] = i[28];
  assign o[14540] = i[28];
  assign o[14541] = i[28];
  assign o[14542] = i[28];
  assign o[14543] = i[28];
  assign o[14544] = i[28];
  assign o[14545] = i[28];
  assign o[14546] = i[28];
  assign o[14547] = i[28];
  assign o[14548] = i[28];
  assign o[14549] = i[28];
  assign o[14550] = i[28];
  assign o[14551] = i[28];
  assign o[14552] = i[28];
  assign o[14553] = i[28];
  assign o[14554] = i[28];
  assign o[14555] = i[28];
  assign o[14556] = i[28];
  assign o[14557] = i[28];
  assign o[14558] = i[28];
  assign o[14559] = i[28];
  assign o[14560] = i[28];
  assign o[14561] = i[28];
  assign o[14562] = i[28];
  assign o[14563] = i[28];
  assign o[14564] = i[28];
  assign o[14565] = i[28];
  assign o[14566] = i[28];
  assign o[14567] = i[28];
  assign o[14568] = i[28];
  assign o[14569] = i[28];
  assign o[14570] = i[28];
  assign o[14571] = i[28];
  assign o[14572] = i[28];
  assign o[14573] = i[28];
  assign o[14574] = i[28];
  assign o[14575] = i[28];
  assign o[14576] = i[28];
  assign o[14577] = i[28];
  assign o[14578] = i[28];
  assign o[14579] = i[28];
  assign o[14580] = i[28];
  assign o[14581] = i[28];
  assign o[14582] = i[28];
  assign o[14583] = i[28];
  assign o[14584] = i[28];
  assign o[14585] = i[28];
  assign o[14586] = i[28];
  assign o[14587] = i[28];
  assign o[14588] = i[28];
  assign o[14589] = i[28];
  assign o[14590] = i[28];
  assign o[14591] = i[28];
  assign o[14592] = i[28];
  assign o[14593] = i[28];
  assign o[14594] = i[28];
  assign o[14595] = i[28];
  assign o[14596] = i[28];
  assign o[14597] = i[28];
  assign o[14598] = i[28];
  assign o[14599] = i[28];
  assign o[14600] = i[28];
  assign o[14601] = i[28];
  assign o[14602] = i[28];
  assign o[14603] = i[28];
  assign o[14604] = i[28];
  assign o[14605] = i[28];
  assign o[14606] = i[28];
  assign o[14607] = i[28];
  assign o[14608] = i[28];
  assign o[14609] = i[28];
  assign o[14610] = i[28];
  assign o[14611] = i[28];
  assign o[14612] = i[28];
  assign o[14613] = i[28];
  assign o[14614] = i[28];
  assign o[14615] = i[28];
  assign o[14616] = i[28];
  assign o[14617] = i[28];
  assign o[14618] = i[28];
  assign o[14619] = i[28];
  assign o[14620] = i[28];
  assign o[14621] = i[28];
  assign o[14622] = i[28];
  assign o[14623] = i[28];
  assign o[14624] = i[28];
  assign o[14625] = i[28];
  assign o[14626] = i[28];
  assign o[14627] = i[28];
  assign o[14628] = i[28];
  assign o[14629] = i[28];
  assign o[14630] = i[28];
  assign o[14631] = i[28];
  assign o[14632] = i[28];
  assign o[14633] = i[28];
  assign o[14634] = i[28];
  assign o[14635] = i[28];
  assign o[14636] = i[28];
  assign o[14637] = i[28];
  assign o[14638] = i[28];
  assign o[14639] = i[28];
  assign o[14640] = i[28];
  assign o[14641] = i[28];
  assign o[14642] = i[28];
  assign o[14643] = i[28];
  assign o[14644] = i[28];
  assign o[14645] = i[28];
  assign o[14646] = i[28];
  assign o[14647] = i[28];
  assign o[14648] = i[28];
  assign o[14649] = i[28];
  assign o[14650] = i[28];
  assign o[14651] = i[28];
  assign o[14652] = i[28];
  assign o[14653] = i[28];
  assign o[14654] = i[28];
  assign o[14655] = i[28];
  assign o[14656] = i[28];
  assign o[14657] = i[28];
  assign o[14658] = i[28];
  assign o[14659] = i[28];
  assign o[14660] = i[28];
  assign o[14661] = i[28];
  assign o[14662] = i[28];
  assign o[14663] = i[28];
  assign o[14664] = i[28];
  assign o[14665] = i[28];
  assign o[14666] = i[28];
  assign o[14667] = i[28];
  assign o[14668] = i[28];
  assign o[14669] = i[28];
  assign o[14670] = i[28];
  assign o[14671] = i[28];
  assign o[14672] = i[28];
  assign o[14673] = i[28];
  assign o[14674] = i[28];
  assign o[14675] = i[28];
  assign o[14676] = i[28];
  assign o[14677] = i[28];
  assign o[14678] = i[28];
  assign o[14679] = i[28];
  assign o[14680] = i[28];
  assign o[14681] = i[28];
  assign o[14682] = i[28];
  assign o[14683] = i[28];
  assign o[14684] = i[28];
  assign o[14685] = i[28];
  assign o[14686] = i[28];
  assign o[14687] = i[28];
  assign o[14688] = i[28];
  assign o[14689] = i[28];
  assign o[14690] = i[28];
  assign o[14691] = i[28];
  assign o[14692] = i[28];
  assign o[14693] = i[28];
  assign o[14694] = i[28];
  assign o[14695] = i[28];
  assign o[14696] = i[28];
  assign o[14697] = i[28];
  assign o[14698] = i[28];
  assign o[14699] = i[28];
  assign o[14700] = i[28];
  assign o[14701] = i[28];
  assign o[14702] = i[28];
  assign o[14703] = i[28];
  assign o[14704] = i[28];
  assign o[14705] = i[28];
  assign o[14706] = i[28];
  assign o[14707] = i[28];
  assign o[14708] = i[28];
  assign o[14709] = i[28];
  assign o[14710] = i[28];
  assign o[14711] = i[28];
  assign o[14712] = i[28];
  assign o[14713] = i[28];
  assign o[14714] = i[28];
  assign o[14715] = i[28];
  assign o[14716] = i[28];
  assign o[14717] = i[28];
  assign o[14718] = i[28];
  assign o[14719] = i[28];
  assign o[14720] = i[28];
  assign o[14721] = i[28];
  assign o[14722] = i[28];
  assign o[14723] = i[28];
  assign o[14724] = i[28];
  assign o[14725] = i[28];
  assign o[14726] = i[28];
  assign o[14727] = i[28];
  assign o[14728] = i[28];
  assign o[14729] = i[28];
  assign o[14730] = i[28];
  assign o[14731] = i[28];
  assign o[14732] = i[28];
  assign o[14733] = i[28];
  assign o[14734] = i[28];
  assign o[14735] = i[28];
  assign o[14736] = i[28];
  assign o[14737] = i[28];
  assign o[14738] = i[28];
  assign o[14739] = i[28];
  assign o[14740] = i[28];
  assign o[14741] = i[28];
  assign o[14742] = i[28];
  assign o[14743] = i[28];
  assign o[14744] = i[28];
  assign o[14745] = i[28];
  assign o[14746] = i[28];
  assign o[14747] = i[28];
  assign o[14748] = i[28];
  assign o[14749] = i[28];
  assign o[14750] = i[28];
  assign o[14751] = i[28];
  assign o[14752] = i[28];
  assign o[14753] = i[28];
  assign o[14754] = i[28];
  assign o[14755] = i[28];
  assign o[14756] = i[28];
  assign o[14757] = i[28];
  assign o[14758] = i[28];
  assign o[14759] = i[28];
  assign o[14760] = i[28];
  assign o[14761] = i[28];
  assign o[14762] = i[28];
  assign o[14763] = i[28];
  assign o[14764] = i[28];
  assign o[14765] = i[28];
  assign o[14766] = i[28];
  assign o[14767] = i[28];
  assign o[14768] = i[28];
  assign o[14769] = i[28];
  assign o[14770] = i[28];
  assign o[14771] = i[28];
  assign o[14772] = i[28];
  assign o[14773] = i[28];
  assign o[14774] = i[28];
  assign o[14775] = i[28];
  assign o[14776] = i[28];
  assign o[14777] = i[28];
  assign o[14778] = i[28];
  assign o[14779] = i[28];
  assign o[14780] = i[28];
  assign o[14781] = i[28];
  assign o[14782] = i[28];
  assign o[14783] = i[28];
  assign o[14784] = i[28];
  assign o[14785] = i[28];
  assign o[14786] = i[28];
  assign o[14787] = i[28];
  assign o[14788] = i[28];
  assign o[14789] = i[28];
  assign o[14790] = i[28];
  assign o[14791] = i[28];
  assign o[14792] = i[28];
  assign o[14793] = i[28];
  assign o[14794] = i[28];
  assign o[14795] = i[28];
  assign o[14796] = i[28];
  assign o[14797] = i[28];
  assign o[14798] = i[28];
  assign o[14799] = i[28];
  assign o[14800] = i[28];
  assign o[14801] = i[28];
  assign o[14802] = i[28];
  assign o[14803] = i[28];
  assign o[14804] = i[28];
  assign o[14805] = i[28];
  assign o[14806] = i[28];
  assign o[14807] = i[28];
  assign o[14808] = i[28];
  assign o[14809] = i[28];
  assign o[14810] = i[28];
  assign o[14811] = i[28];
  assign o[14812] = i[28];
  assign o[14813] = i[28];
  assign o[14814] = i[28];
  assign o[14815] = i[28];
  assign o[14816] = i[28];
  assign o[14817] = i[28];
  assign o[14818] = i[28];
  assign o[14819] = i[28];
  assign o[14820] = i[28];
  assign o[14821] = i[28];
  assign o[14822] = i[28];
  assign o[14823] = i[28];
  assign o[14824] = i[28];
  assign o[14825] = i[28];
  assign o[14826] = i[28];
  assign o[14827] = i[28];
  assign o[14828] = i[28];
  assign o[14829] = i[28];
  assign o[14830] = i[28];
  assign o[14831] = i[28];
  assign o[14832] = i[28];
  assign o[14833] = i[28];
  assign o[14834] = i[28];
  assign o[14835] = i[28];
  assign o[14836] = i[28];
  assign o[14837] = i[28];
  assign o[14838] = i[28];
  assign o[14839] = i[28];
  assign o[14840] = i[28];
  assign o[14841] = i[28];
  assign o[14842] = i[28];
  assign o[14843] = i[28];
  assign o[14844] = i[28];
  assign o[14845] = i[28];
  assign o[14846] = i[28];
  assign o[14847] = i[28];
  assign o[13824] = i[27];
  assign o[13825] = i[27];
  assign o[13826] = i[27];
  assign o[13827] = i[27];
  assign o[13828] = i[27];
  assign o[13829] = i[27];
  assign o[13830] = i[27];
  assign o[13831] = i[27];
  assign o[13832] = i[27];
  assign o[13833] = i[27];
  assign o[13834] = i[27];
  assign o[13835] = i[27];
  assign o[13836] = i[27];
  assign o[13837] = i[27];
  assign o[13838] = i[27];
  assign o[13839] = i[27];
  assign o[13840] = i[27];
  assign o[13841] = i[27];
  assign o[13842] = i[27];
  assign o[13843] = i[27];
  assign o[13844] = i[27];
  assign o[13845] = i[27];
  assign o[13846] = i[27];
  assign o[13847] = i[27];
  assign o[13848] = i[27];
  assign o[13849] = i[27];
  assign o[13850] = i[27];
  assign o[13851] = i[27];
  assign o[13852] = i[27];
  assign o[13853] = i[27];
  assign o[13854] = i[27];
  assign o[13855] = i[27];
  assign o[13856] = i[27];
  assign o[13857] = i[27];
  assign o[13858] = i[27];
  assign o[13859] = i[27];
  assign o[13860] = i[27];
  assign o[13861] = i[27];
  assign o[13862] = i[27];
  assign o[13863] = i[27];
  assign o[13864] = i[27];
  assign o[13865] = i[27];
  assign o[13866] = i[27];
  assign o[13867] = i[27];
  assign o[13868] = i[27];
  assign o[13869] = i[27];
  assign o[13870] = i[27];
  assign o[13871] = i[27];
  assign o[13872] = i[27];
  assign o[13873] = i[27];
  assign o[13874] = i[27];
  assign o[13875] = i[27];
  assign o[13876] = i[27];
  assign o[13877] = i[27];
  assign o[13878] = i[27];
  assign o[13879] = i[27];
  assign o[13880] = i[27];
  assign o[13881] = i[27];
  assign o[13882] = i[27];
  assign o[13883] = i[27];
  assign o[13884] = i[27];
  assign o[13885] = i[27];
  assign o[13886] = i[27];
  assign o[13887] = i[27];
  assign o[13888] = i[27];
  assign o[13889] = i[27];
  assign o[13890] = i[27];
  assign o[13891] = i[27];
  assign o[13892] = i[27];
  assign o[13893] = i[27];
  assign o[13894] = i[27];
  assign o[13895] = i[27];
  assign o[13896] = i[27];
  assign o[13897] = i[27];
  assign o[13898] = i[27];
  assign o[13899] = i[27];
  assign o[13900] = i[27];
  assign o[13901] = i[27];
  assign o[13902] = i[27];
  assign o[13903] = i[27];
  assign o[13904] = i[27];
  assign o[13905] = i[27];
  assign o[13906] = i[27];
  assign o[13907] = i[27];
  assign o[13908] = i[27];
  assign o[13909] = i[27];
  assign o[13910] = i[27];
  assign o[13911] = i[27];
  assign o[13912] = i[27];
  assign o[13913] = i[27];
  assign o[13914] = i[27];
  assign o[13915] = i[27];
  assign o[13916] = i[27];
  assign o[13917] = i[27];
  assign o[13918] = i[27];
  assign o[13919] = i[27];
  assign o[13920] = i[27];
  assign o[13921] = i[27];
  assign o[13922] = i[27];
  assign o[13923] = i[27];
  assign o[13924] = i[27];
  assign o[13925] = i[27];
  assign o[13926] = i[27];
  assign o[13927] = i[27];
  assign o[13928] = i[27];
  assign o[13929] = i[27];
  assign o[13930] = i[27];
  assign o[13931] = i[27];
  assign o[13932] = i[27];
  assign o[13933] = i[27];
  assign o[13934] = i[27];
  assign o[13935] = i[27];
  assign o[13936] = i[27];
  assign o[13937] = i[27];
  assign o[13938] = i[27];
  assign o[13939] = i[27];
  assign o[13940] = i[27];
  assign o[13941] = i[27];
  assign o[13942] = i[27];
  assign o[13943] = i[27];
  assign o[13944] = i[27];
  assign o[13945] = i[27];
  assign o[13946] = i[27];
  assign o[13947] = i[27];
  assign o[13948] = i[27];
  assign o[13949] = i[27];
  assign o[13950] = i[27];
  assign o[13951] = i[27];
  assign o[13952] = i[27];
  assign o[13953] = i[27];
  assign o[13954] = i[27];
  assign o[13955] = i[27];
  assign o[13956] = i[27];
  assign o[13957] = i[27];
  assign o[13958] = i[27];
  assign o[13959] = i[27];
  assign o[13960] = i[27];
  assign o[13961] = i[27];
  assign o[13962] = i[27];
  assign o[13963] = i[27];
  assign o[13964] = i[27];
  assign o[13965] = i[27];
  assign o[13966] = i[27];
  assign o[13967] = i[27];
  assign o[13968] = i[27];
  assign o[13969] = i[27];
  assign o[13970] = i[27];
  assign o[13971] = i[27];
  assign o[13972] = i[27];
  assign o[13973] = i[27];
  assign o[13974] = i[27];
  assign o[13975] = i[27];
  assign o[13976] = i[27];
  assign o[13977] = i[27];
  assign o[13978] = i[27];
  assign o[13979] = i[27];
  assign o[13980] = i[27];
  assign o[13981] = i[27];
  assign o[13982] = i[27];
  assign o[13983] = i[27];
  assign o[13984] = i[27];
  assign o[13985] = i[27];
  assign o[13986] = i[27];
  assign o[13987] = i[27];
  assign o[13988] = i[27];
  assign o[13989] = i[27];
  assign o[13990] = i[27];
  assign o[13991] = i[27];
  assign o[13992] = i[27];
  assign o[13993] = i[27];
  assign o[13994] = i[27];
  assign o[13995] = i[27];
  assign o[13996] = i[27];
  assign o[13997] = i[27];
  assign o[13998] = i[27];
  assign o[13999] = i[27];
  assign o[14000] = i[27];
  assign o[14001] = i[27];
  assign o[14002] = i[27];
  assign o[14003] = i[27];
  assign o[14004] = i[27];
  assign o[14005] = i[27];
  assign o[14006] = i[27];
  assign o[14007] = i[27];
  assign o[14008] = i[27];
  assign o[14009] = i[27];
  assign o[14010] = i[27];
  assign o[14011] = i[27];
  assign o[14012] = i[27];
  assign o[14013] = i[27];
  assign o[14014] = i[27];
  assign o[14015] = i[27];
  assign o[14016] = i[27];
  assign o[14017] = i[27];
  assign o[14018] = i[27];
  assign o[14019] = i[27];
  assign o[14020] = i[27];
  assign o[14021] = i[27];
  assign o[14022] = i[27];
  assign o[14023] = i[27];
  assign o[14024] = i[27];
  assign o[14025] = i[27];
  assign o[14026] = i[27];
  assign o[14027] = i[27];
  assign o[14028] = i[27];
  assign o[14029] = i[27];
  assign o[14030] = i[27];
  assign o[14031] = i[27];
  assign o[14032] = i[27];
  assign o[14033] = i[27];
  assign o[14034] = i[27];
  assign o[14035] = i[27];
  assign o[14036] = i[27];
  assign o[14037] = i[27];
  assign o[14038] = i[27];
  assign o[14039] = i[27];
  assign o[14040] = i[27];
  assign o[14041] = i[27];
  assign o[14042] = i[27];
  assign o[14043] = i[27];
  assign o[14044] = i[27];
  assign o[14045] = i[27];
  assign o[14046] = i[27];
  assign o[14047] = i[27];
  assign o[14048] = i[27];
  assign o[14049] = i[27];
  assign o[14050] = i[27];
  assign o[14051] = i[27];
  assign o[14052] = i[27];
  assign o[14053] = i[27];
  assign o[14054] = i[27];
  assign o[14055] = i[27];
  assign o[14056] = i[27];
  assign o[14057] = i[27];
  assign o[14058] = i[27];
  assign o[14059] = i[27];
  assign o[14060] = i[27];
  assign o[14061] = i[27];
  assign o[14062] = i[27];
  assign o[14063] = i[27];
  assign o[14064] = i[27];
  assign o[14065] = i[27];
  assign o[14066] = i[27];
  assign o[14067] = i[27];
  assign o[14068] = i[27];
  assign o[14069] = i[27];
  assign o[14070] = i[27];
  assign o[14071] = i[27];
  assign o[14072] = i[27];
  assign o[14073] = i[27];
  assign o[14074] = i[27];
  assign o[14075] = i[27];
  assign o[14076] = i[27];
  assign o[14077] = i[27];
  assign o[14078] = i[27];
  assign o[14079] = i[27];
  assign o[14080] = i[27];
  assign o[14081] = i[27];
  assign o[14082] = i[27];
  assign o[14083] = i[27];
  assign o[14084] = i[27];
  assign o[14085] = i[27];
  assign o[14086] = i[27];
  assign o[14087] = i[27];
  assign o[14088] = i[27];
  assign o[14089] = i[27];
  assign o[14090] = i[27];
  assign o[14091] = i[27];
  assign o[14092] = i[27];
  assign o[14093] = i[27];
  assign o[14094] = i[27];
  assign o[14095] = i[27];
  assign o[14096] = i[27];
  assign o[14097] = i[27];
  assign o[14098] = i[27];
  assign o[14099] = i[27];
  assign o[14100] = i[27];
  assign o[14101] = i[27];
  assign o[14102] = i[27];
  assign o[14103] = i[27];
  assign o[14104] = i[27];
  assign o[14105] = i[27];
  assign o[14106] = i[27];
  assign o[14107] = i[27];
  assign o[14108] = i[27];
  assign o[14109] = i[27];
  assign o[14110] = i[27];
  assign o[14111] = i[27];
  assign o[14112] = i[27];
  assign o[14113] = i[27];
  assign o[14114] = i[27];
  assign o[14115] = i[27];
  assign o[14116] = i[27];
  assign o[14117] = i[27];
  assign o[14118] = i[27];
  assign o[14119] = i[27];
  assign o[14120] = i[27];
  assign o[14121] = i[27];
  assign o[14122] = i[27];
  assign o[14123] = i[27];
  assign o[14124] = i[27];
  assign o[14125] = i[27];
  assign o[14126] = i[27];
  assign o[14127] = i[27];
  assign o[14128] = i[27];
  assign o[14129] = i[27];
  assign o[14130] = i[27];
  assign o[14131] = i[27];
  assign o[14132] = i[27];
  assign o[14133] = i[27];
  assign o[14134] = i[27];
  assign o[14135] = i[27];
  assign o[14136] = i[27];
  assign o[14137] = i[27];
  assign o[14138] = i[27];
  assign o[14139] = i[27];
  assign o[14140] = i[27];
  assign o[14141] = i[27];
  assign o[14142] = i[27];
  assign o[14143] = i[27];
  assign o[14144] = i[27];
  assign o[14145] = i[27];
  assign o[14146] = i[27];
  assign o[14147] = i[27];
  assign o[14148] = i[27];
  assign o[14149] = i[27];
  assign o[14150] = i[27];
  assign o[14151] = i[27];
  assign o[14152] = i[27];
  assign o[14153] = i[27];
  assign o[14154] = i[27];
  assign o[14155] = i[27];
  assign o[14156] = i[27];
  assign o[14157] = i[27];
  assign o[14158] = i[27];
  assign o[14159] = i[27];
  assign o[14160] = i[27];
  assign o[14161] = i[27];
  assign o[14162] = i[27];
  assign o[14163] = i[27];
  assign o[14164] = i[27];
  assign o[14165] = i[27];
  assign o[14166] = i[27];
  assign o[14167] = i[27];
  assign o[14168] = i[27];
  assign o[14169] = i[27];
  assign o[14170] = i[27];
  assign o[14171] = i[27];
  assign o[14172] = i[27];
  assign o[14173] = i[27];
  assign o[14174] = i[27];
  assign o[14175] = i[27];
  assign o[14176] = i[27];
  assign o[14177] = i[27];
  assign o[14178] = i[27];
  assign o[14179] = i[27];
  assign o[14180] = i[27];
  assign o[14181] = i[27];
  assign o[14182] = i[27];
  assign o[14183] = i[27];
  assign o[14184] = i[27];
  assign o[14185] = i[27];
  assign o[14186] = i[27];
  assign o[14187] = i[27];
  assign o[14188] = i[27];
  assign o[14189] = i[27];
  assign o[14190] = i[27];
  assign o[14191] = i[27];
  assign o[14192] = i[27];
  assign o[14193] = i[27];
  assign o[14194] = i[27];
  assign o[14195] = i[27];
  assign o[14196] = i[27];
  assign o[14197] = i[27];
  assign o[14198] = i[27];
  assign o[14199] = i[27];
  assign o[14200] = i[27];
  assign o[14201] = i[27];
  assign o[14202] = i[27];
  assign o[14203] = i[27];
  assign o[14204] = i[27];
  assign o[14205] = i[27];
  assign o[14206] = i[27];
  assign o[14207] = i[27];
  assign o[14208] = i[27];
  assign o[14209] = i[27];
  assign o[14210] = i[27];
  assign o[14211] = i[27];
  assign o[14212] = i[27];
  assign o[14213] = i[27];
  assign o[14214] = i[27];
  assign o[14215] = i[27];
  assign o[14216] = i[27];
  assign o[14217] = i[27];
  assign o[14218] = i[27];
  assign o[14219] = i[27];
  assign o[14220] = i[27];
  assign o[14221] = i[27];
  assign o[14222] = i[27];
  assign o[14223] = i[27];
  assign o[14224] = i[27];
  assign o[14225] = i[27];
  assign o[14226] = i[27];
  assign o[14227] = i[27];
  assign o[14228] = i[27];
  assign o[14229] = i[27];
  assign o[14230] = i[27];
  assign o[14231] = i[27];
  assign o[14232] = i[27];
  assign o[14233] = i[27];
  assign o[14234] = i[27];
  assign o[14235] = i[27];
  assign o[14236] = i[27];
  assign o[14237] = i[27];
  assign o[14238] = i[27];
  assign o[14239] = i[27];
  assign o[14240] = i[27];
  assign o[14241] = i[27];
  assign o[14242] = i[27];
  assign o[14243] = i[27];
  assign o[14244] = i[27];
  assign o[14245] = i[27];
  assign o[14246] = i[27];
  assign o[14247] = i[27];
  assign o[14248] = i[27];
  assign o[14249] = i[27];
  assign o[14250] = i[27];
  assign o[14251] = i[27];
  assign o[14252] = i[27];
  assign o[14253] = i[27];
  assign o[14254] = i[27];
  assign o[14255] = i[27];
  assign o[14256] = i[27];
  assign o[14257] = i[27];
  assign o[14258] = i[27];
  assign o[14259] = i[27];
  assign o[14260] = i[27];
  assign o[14261] = i[27];
  assign o[14262] = i[27];
  assign o[14263] = i[27];
  assign o[14264] = i[27];
  assign o[14265] = i[27];
  assign o[14266] = i[27];
  assign o[14267] = i[27];
  assign o[14268] = i[27];
  assign o[14269] = i[27];
  assign o[14270] = i[27];
  assign o[14271] = i[27];
  assign o[14272] = i[27];
  assign o[14273] = i[27];
  assign o[14274] = i[27];
  assign o[14275] = i[27];
  assign o[14276] = i[27];
  assign o[14277] = i[27];
  assign o[14278] = i[27];
  assign o[14279] = i[27];
  assign o[14280] = i[27];
  assign o[14281] = i[27];
  assign o[14282] = i[27];
  assign o[14283] = i[27];
  assign o[14284] = i[27];
  assign o[14285] = i[27];
  assign o[14286] = i[27];
  assign o[14287] = i[27];
  assign o[14288] = i[27];
  assign o[14289] = i[27];
  assign o[14290] = i[27];
  assign o[14291] = i[27];
  assign o[14292] = i[27];
  assign o[14293] = i[27];
  assign o[14294] = i[27];
  assign o[14295] = i[27];
  assign o[14296] = i[27];
  assign o[14297] = i[27];
  assign o[14298] = i[27];
  assign o[14299] = i[27];
  assign o[14300] = i[27];
  assign o[14301] = i[27];
  assign o[14302] = i[27];
  assign o[14303] = i[27];
  assign o[14304] = i[27];
  assign o[14305] = i[27];
  assign o[14306] = i[27];
  assign o[14307] = i[27];
  assign o[14308] = i[27];
  assign o[14309] = i[27];
  assign o[14310] = i[27];
  assign o[14311] = i[27];
  assign o[14312] = i[27];
  assign o[14313] = i[27];
  assign o[14314] = i[27];
  assign o[14315] = i[27];
  assign o[14316] = i[27];
  assign o[14317] = i[27];
  assign o[14318] = i[27];
  assign o[14319] = i[27];
  assign o[14320] = i[27];
  assign o[14321] = i[27];
  assign o[14322] = i[27];
  assign o[14323] = i[27];
  assign o[14324] = i[27];
  assign o[14325] = i[27];
  assign o[14326] = i[27];
  assign o[14327] = i[27];
  assign o[14328] = i[27];
  assign o[14329] = i[27];
  assign o[14330] = i[27];
  assign o[14331] = i[27];
  assign o[14332] = i[27];
  assign o[14333] = i[27];
  assign o[14334] = i[27];
  assign o[14335] = i[27];
  assign o[13312] = i[26];
  assign o[13313] = i[26];
  assign o[13314] = i[26];
  assign o[13315] = i[26];
  assign o[13316] = i[26];
  assign o[13317] = i[26];
  assign o[13318] = i[26];
  assign o[13319] = i[26];
  assign o[13320] = i[26];
  assign o[13321] = i[26];
  assign o[13322] = i[26];
  assign o[13323] = i[26];
  assign o[13324] = i[26];
  assign o[13325] = i[26];
  assign o[13326] = i[26];
  assign o[13327] = i[26];
  assign o[13328] = i[26];
  assign o[13329] = i[26];
  assign o[13330] = i[26];
  assign o[13331] = i[26];
  assign o[13332] = i[26];
  assign o[13333] = i[26];
  assign o[13334] = i[26];
  assign o[13335] = i[26];
  assign o[13336] = i[26];
  assign o[13337] = i[26];
  assign o[13338] = i[26];
  assign o[13339] = i[26];
  assign o[13340] = i[26];
  assign o[13341] = i[26];
  assign o[13342] = i[26];
  assign o[13343] = i[26];
  assign o[13344] = i[26];
  assign o[13345] = i[26];
  assign o[13346] = i[26];
  assign o[13347] = i[26];
  assign o[13348] = i[26];
  assign o[13349] = i[26];
  assign o[13350] = i[26];
  assign o[13351] = i[26];
  assign o[13352] = i[26];
  assign o[13353] = i[26];
  assign o[13354] = i[26];
  assign o[13355] = i[26];
  assign o[13356] = i[26];
  assign o[13357] = i[26];
  assign o[13358] = i[26];
  assign o[13359] = i[26];
  assign o[13360] = i[26];
  assign o[13361] = i[26];
  assign o[13362] = i[26];
  assign o[13363] = i[26];
  assign o[13364] = i[26];
  assign o[13365] = i[26];
  assign o[13366] = i[26];
  assign o[13367] = i[26];
  assign o[13368] = i[26];
  assign o[13369] = i[26];
  assign o[13370] = i[26];
  assign o[13371] = i[26];
  assign o[13372] = i[26];
  assign o[13373] = i[26];
  assign o[13374] = i[26];
  assign o[13375] = i[26];
  assign o[13376] = i[26];
  assign o[13377] = i[26];
  assign o[13378] = i[26];
  assign o[13379] = i[26];
  assign o[13380] = i[26];
  assign o[13381] = i[26];
  assign o[13382] = i[26];
  assign o[13383] = i[26];
  assign o[13384] = i[26];
  assign o[13385] = i[26];
  assign o[13386] = i[26];
  assign o[13387] = i[26];
  assign o[13388] = i[26];
  assign o[13389] = i[26];
  assign o[13390] = i[26];
  assign o[13391] = i[26];
  assign o[13392] = i[26];
  assign o[13393] = i[26];
  assign o[13394] = i[26];
  assign o[13395] = i[26];
  assign o[13396] = i[26];
  assign o[13397] = i[26];
  assign o[13398] = i[26];
  assign o[13399] = i[26];
  assign o[13400] = i[26];
  assign o[13401] = i[26];
  assign o[13402] = i[26];
  assign o[13403] = i[26];
  assign o[13404] = i[26];
  assign o[13405] = i[26];
  assign o[13406] = i[26];
  assign o[13407] = i[26];
  assign o[13408] = i[26];
  assign o[13409] = i[26];
  assign o[13410] = i[26];
  assign o[13411] = i[26];
  assign o[13412] = i[26];
  assign o[13413] = i[26];
  assign o[13414] = i[26];
  assign o[13415] = i[26];
  assign o[13416] = i[26];
  assign o[13417] = i[26];
  assign o[13418] = i[26];
  assign o[13419] = i[26];
  assign o[13420] = i[26];
  assign o[13421] = i[26];
  assign o[13422] = i[26];
  assign o[13423] = i[26];
  assign o[13424] = i[26];
  assign o[13425] = i[26];
  assign o[13426] = i[26];
  assign o[13427] = i[26];
  assign o[13428] = i[26];
  assign o[13429] = i[26];
  assign o[13430] = i[26];
  assign o[13431] = i[26];
  assign o[13432] = i[26];
  assign o[13433] = i[26];
  assign o[13434] = i[26];
  assign o[13435] = i[26];
  assign o[13436] = i[26];
  assign o[13437] = i[26];
  assign o[13438] = i[26];
  assign o[13439] = i[26];
  assign o[13440] = i[26];
  assign o[13441] = i[26];
  assign o[13442] = i[26];
  assign o[13443] = i[26];
  assign o[13444] = i[26];
  assign o[13445] = i[26];
  assign o[13446] = i[26];
  assign o[13447] = i[26];
  assign o[13448] = i[26];
  assign o[13449] = i[26];
  assign o[13450] = i[26];
  assign o[13451] = i[26];
  assign o[13452] = i[26];
  assign o[13453] = i[26];
  assign o[13454] = i[26];
  assign o[13455] = i[26];
  assign o[13456] = i[26];
  assign o[13457] = i[26];
  assign o[13458] = i[26];
  assign o[13459] = i[26];
  assign o[13460] = i[26];
  assign o[13461] = i[26];
  assign o[13462] = i[26];
  assign o[13463] = i[26];
  assign o[13464] = i[26];
  assign o[13465] = i[26];
  assign o[13466] = i[26];
  assign o[13467] = i[26];
  assign o[13468] = i[26];
  assign o[13469] = i[26];
  assign o[13470] = i[26];
  assign o[13471] = i[26];
  assign o[13472] = i[26];
  assign o[13473] = i[26];
  assign o[13474] = i[26];
  assign o[13475] = i[26];
  assign o[13476] = i[26];
  assign o[13477] = i[26];
  assign o[13478] = i[26];
  assign o[13479] = i[26];
  assign o[13480] = i[26];
  assign o[13481] = i[26];
  assign o[13482] = i[26];
  assign o[13483] = i[26];
  assign o[13484] = i[26];
  assign o[13485] = i[26];
  assign o[13486] = i[26];
  assign o[13487] = i[26];
  assign o[13488] = i[26];
  assign o[13489] = i[26];
  assign o[13490] = i[26];
  assign o[13491] = i[26];
  assign o[13492] = i[26];
  assign o[13493] = i[26];
  assign o[13494] = i[26];
  assign o[13495] = i[26];
  assign o[13496] = i[26];
  assign o[13497] = i[26];
  assign o[13498] = i[26];
  assign o[13499] = i[26];
  assign o[13500] = i[26];
  assign o[13501] = i[26];
  assign o[13502] = i[26];
  assign o[13503] = i[26];
  assign o[13504] = i[26];
  assign o[13505] = i[26];
  assign o[13506] = i[26];
  assign o[13507] = i[26];
  assign o[13508] = i[26];
  assign o[13509] = i[26];
  assign o[13510] = i[26];
  assign o[13511] = i[26];
  assign o[13512] = i[26];
  assign o[13513] = i[26];
  assign o[13514] = i[26];
  assign o[13515] = i[26];
  assign o[13516] = i[26];
  assign o[13517] = i[26];
  assign o[13518] = i[26];
  assign o[13519] = i[26];
  assign o[13520] = i[26];
  assign o[13521] = i[26];
  assign o[13522] = i[26];
  assign o[13523] = i[26];
  assign o[13524] = i[26];
  assign o[13525] = i[26];
  assign o[13526] = i[26];
  assign o[13527] = i[26];
  assign o[13528] = i[26];
  assign o[13529] = i[26];
  assign o[13530] = i[26];
  assign o[13531] = i[26];
  assign o[13532] = i[26];
  assign o[13533] = i[26];
  assign o[13534] = i[26];
  assign o[13535] = i[26];
  assign o[13536] = i[26];
  assign o[13537] = i[26];
  assign o[13538] = i[26];
  assign o[13539] = i[26];
  assign o[13540] = i[26];
  assign o[13541] = i[26];
  assign o[13542] = i[26];
  assign o[13543] = i[26];
  assign o[13544] = i[26];
  assign o[13545] = i[26];
  assign o[13546] = i[26];
  assign o[13547] = i[26];
  assign o[13548] = i[26];
  assign o[13549] = i[26];
  assign o[13550] = i[26];
  assign o[13551] = i[26];
  assign o[13552] = i[26];
  assign o[13553] = i[26];
  assign o[13554] = i[26];
  assign o[13555] = i[26];
  assign o[13556] = i[26];
  assign o[13557] = i[26];
  assign o[13558] = i[26];
  assign o[13559] = i[26];
  assign o[13560] = i[26];
  assign o[13561] = i[26];
  assign o[13562] = i[26];
  assign o[13563] = i[26];
  assign o[13564] = i[26];
  assign o[13565] = i[26];
  assign o[13566] = i[26];
  assign o[13567] = i[26];
  assign o[13568] = i[26];
  assign o[13569] = i[26];
  assign o[13570] = i[26];
  assign o[13571] = i[26];
  assign o[13572] = i[26];
  assign o[13573] = i[26];
  assign o[13574] = i[26];
  assign o[13575] = i[26];
  assign o[13576] = i[26];
  assign o[13577] = i[26];
  assign o[13578] = i[26];
  assign o[13579] = i[26];
  assign o[13580] = i[26];
  assign o[13581] = i[26];
  assign o[13582] = i[26];
  assign o[13583] = i[26];
  assign o[13584] = i[26];
  assign o[13585] = i[26];
  assign o[13586] = i[26];
  assign o[13587] = i[26];
  assign o[13588] = i[26];
  assign o[13589] = i[26];
  assign o[13590] = i[26];
  assign o[13591] = i[26];
  assign o[13592] = i[26];
  assign o[13593] = i[26];
  assign o[13594] = i[26];
  assign o[13595] = i[26];
  assign o[13596] = i[26];
  assign o[13597] = i[26];
  assign o[13598] = i[26];
  assign o[13599] = i[26];
  assign o[13600] = i[26];
  assign o[13601] = i[26];
  assign o[13602] = i[26];
  assign o[13603] = i[26];
  assign o[13604] = i[26];
  assign o[13605] = i[26];
  assign o[13606] = i[26];
  assign o[13607] = i[26];
  assign o[13608] = i[26];
  assign o[13609] = i[26];
  assign o[13610] = i[26];
  assign o[13611] = i[26];
  assign o[13612] = i[26];
  assign o[13613] = i[26];
  assign o[13614] = i[26];
  assign o[13615] = i[26];
  assign o[13616] = i[26];
  assign o[13617] = i[26];
  assign o[13618] = i[26];
  assign o[13619] = i[26];
  assign o[13620] = i[26];
  assign o[13621] = i[26];
  assign o[13622] = i[26];
  assign o[13623] = i[26];
  assign o[13624] = i[26];
  assign o[13625] = i[26];
  assign o[13626] = i[26];
  assign o[13627] = i[26];
  assign o[13628] = i[26];
  assign o[13629] = i[26];
  assign o[13630] = i[26];
  assign o[13631] = i[26];
  assign o[13632] = i[26];
  assign o[13633] = i[26];
  assign o[13634] = i[26];
  assign o[13635] = i[26];
  assign o[13636] = i[26];
  assign o[13637] = i[26];
  assign o[13638] = i[26];
  assign o[13639] = i[26];
  assign o[13640] = i[26];
  assign o[13641] = i[26];
  assign o[13642] = i[26];
  assign o[13643] = i[26];
  assign o[13644] = i[26];
  assign o[13645] = i[26];
  assign o[13646] = i[26];
  assign o[13647] = i[26];
  assign o[13648] = i[26];
  assign o[13649] = i[26];
  assign o[13650] = i[26];
  assign o[13651] = i[26];
  assign o[13652] = i[26];
  assign o[13653] = i[26];
  assign o[13654] = i[26];
  assign o[13655] = i[26];
  assign o[13656] = i[26];
  assign o[13657] = i[26];
  assign o[13658] = i[26];
  assign o[13659] = i[26];
  assign o[13660] = i[26];
  assign o[13661] = i[26];
  assign o[13662] = i[26];
  assign o[13663] = i[26];
  assign o[13664] = i[26];
  assign o[13665] = i[26];
  assign o[13666] = i[26];
  assign o[13667] = i[26];
  assign o[13668] = i[26];
  assign o[13669] = i[26];
  assign o[13670] = i[26];
  assign o[13671] = i[26];
  assign o[13672] = i[26];
  assign o[13673] = i[26];
  assign o[13674] = i[26];
  assign o[13675] = i[26];
  assign o[13676] = i[26];
  assign o[13677] = i[26];
  assign o[13678] = i[26];
  assign o[13679] = i[26];
  assign o[13680] = i[26];
  assign o[13681] = i[26];
  assign o[13682] = i[26];
  assign o[13683] = i[26];
  assign o[13684] = i[26];
  assign o[13685] = i[26];
  assign o[13686] = i[26];
  assign o[13687] = i[26];
  assign o[13688] = i[26];
  assign o[13689] = i[26];
  assign o[13690] = i[26];
  assign o[13691] = i[26];
  assign o[13692] = i[26];
  assign o[13693] = i[26];
  assign o[13694] = i[26];
  assign o[13695] = i[26];
  assign o[13696] = i[26];
  assign o[13697] = i[26];
  assign o[13698] = i[26];
  assign o[13699] = i[26];
  assign o[13700] = i[26];
  assign o[13701] = i[26];
  assign o[13702] = i[26];
  assign o[13703] = i[26];
  assign o[13704] = i[26];
  assign o[13705] = i[26];
  assign o[13706] = i[26];
  assign o[13707] = i[26];
  assign o[13708] = i[26];
  assign o[13709] = i[26];
  assign o[13710] = i[26];
  assign o[13711] = i[26];
  assign o[13712] = i[26];
  assign o[13713] = i[26];
  assign o[13714] = i[26];
  assign o[13715] = i[26];
  assign o[13716] = i[26];
  assign o[13717] = i[26];
  assign o[13718] = i[26];
  assign o[13719] = i[26];
  assign o[13720] = i[26];
  assign o[13721] = i[26];
  assign o[13722] = i[26];
  assign o[13723] = i[26];
  assign o[13724] = i[26];
  assign o[13725] = i[26];
  assign o[13726] = i[26];
  assign o[13727] = i[26];
  assign o[13728] = i[26];
  assign o[13729] = i[26];
  assign o[13730] = i[26];
  assign o[13731] = i[26];
  assign o[13732] = i[26];
  assign o[13733] = i[26];
  assign o[13734] = i[26];
  assign o[13735] = i[26];
  assign o[13736] = i[26];
  assign o[13737] = i[26];
  assign o[13738] = i[26];
  assign o[13739] = i[26];
  assign o[13740] = i[26];
  assign o[13741] = i[26];
  assign o[13742] = i[26];
  assign o[13743] = i[26];
  assign o[13744] = i[26];
  assign o[13745] = i[26];
  assign o[13746] = i[26];
  assign o[13747] = i[26];
  assign o[13748] = i[26];
  assign o[13749] = i[26];
  assign o[13750] = i[26];
  assign o[13751] = i[26];
  assign o[13752] = i[26];
  assign o[13753] = i[26];
  assign o[13754] = i[26];
  assign o[13755] = i[26];
  assign o[13756] = i[26];
  assign o[13757] = i[26];
  assign o[13758] = i[26];
  assign o[13759] = i[26];
  assign o[13760] = i[26];
  assign o[13761] = i[26];
  assign o[13762] = i[26];
  assign o[13763] = i[26];
  assign o[13764] = i[26];
  assign o[13765] = i[26];
  assign o[13766] = i[26];
  assign o[13767] = i[26];
  assign o[13768] = i[26];
  assign o[13769] = i[26];
  assign o[13770] = i[26];
  assign o[13771] = i[26];
  assign o[13772] = i[26];
  assign o[13773] = i[26];
  assign o[13774] = i[26];
  assign o[13775] = i[26];
  assign o[13776] = i[26];
  assign o[13777] = i[26];
  assign o[13778] = i[26];
  assign o[13779] = i[26];
  assign o[13780] = i[26];
  assign o[13781] = i[26];
  assign o[13782] = i[26];
  assign o[13783] = i[26];
  assign o[13784] = i[26];
  assign o[13785] = i[26];
  assign o[13786] = i[26];
  assign o[13787] = i[26];
  assign o[13788] = i[26];
  assign o[13789] = i[26];
  assign o[13790] = i[26];
  assign o[13791] = i[26];
  assign o[13792] = i[26];
  assign o[13793] = i[26];
  assign o[13794] = i[26];
  assign o[13795] = i[26];
  assign o[13796] = i[26];
  assign o[13797] = i[26];
  assign o[13798] = i[26];
  assign o[13799] = i[26];
  assign o[13800] = i[26];
  assign o[13801] = i[26];
  assign o[13802] = i[26];
  assign o[13803] = i[26];
  assign o[13804] = i[26];
  assign o[13805] = i[26];
  assign o[13806] = i[26];
  assign o[13807] = i[26];
  assign o[13808] = i[26];
  assign o[13809] = i[26];
  assign o[13810] = i[26];
  assign o[13811] = i[26];
  assign o[13812] = i[26];
  assign o[13813] = i[26];
  assign o[13814] = i[26];
  assign o[13815] = i[26];
  assign o[13816] = i[26];
  assign o[13817] = i[26];
  assign o[13818] = i[26];
  assign o[13819] = i[26];
  assign o[13820] = i[26];
  assign o[13821] = i[26];
  assign o[13822] = i[26];
  assign o[13823] = i[26];
  assign o[12800] = i[25];
  assign o[12801] = i[25];
  assign o[12802] = i[25];
  assign o[12803] = i[25];
  assign o[12804] = i[25];
  assign o[12805] = i[25];
  assign o[12806] = i[25];
  assign o[12807] = i[25];
  assign o[12808] = i[25];
  assign o[12809] = i[25];
  assign o[12810] = i[25];
  assign o[12811] = i[25];
  assign o[12812] = i[25];
  assign o[12813] = i[25];
  assign o[12814] = i[25];
  assign o[12815] = i[25];
  assign o[12816] = i[25];
  assign o[12817] = i[25];
  assign o[12818] = i[25];
  assign o[12819] = i[25];
  assign o[12820] = i[25];
  assign o[12821] = i[25];
  assign o[12822] = i[25];
  assign o[12823] = i[25];
  assign o[12824] = i[25];
  assign o[12825] = i[25];
  assign o[12826] = i[25];
  assign o[12827] = i[25];
  assign o[12828] = i[25];
  assign o[12829] = i[25];
  assign o[12830] = i[25];
  assign o[12831] = i[25];
  assign o[12832] = i[25];
  assign o[12833] = i[25];
  assign o[12834] = i[25];
  assign o[12835] = i[25];
  assign o[12836] = i[25];
  assign o[12837] = i[25];
  assign o[12838] = i[25];
  assign o[12839] = i[25];
  assign o[12840] = i[25];
  assign o[12841] = i[25];
  assign o[12842] = i[25];
  assign o[12843] = i[25];
  assign o[12844] = i[25];
  assign o[12845] = i[25];
  assign o[12846] = i[25];
  assign o[12847] = i[25];
  assign o[12848] = i[25];
  assign o[12849] = i[25];
  assign o[12850] = i[25];
  assign o[12851] = i[25];
  assign o[12852] = i[25];
  assign o[12853] = i[25];
  assign o[12854] = i[25];
  assign o[12855] = i[25];
  assign o[12856] = i[25];
  assign o[12857] = i[25];
  assign o[12858] = i[25];
  assign o[12859] = i[25];
  assign o[12860] = i[25];
  assign o[12861] = i[25];
  assign o[12862] = i[25];
  assign o[12863] = i[25];
  assign o[12864] = i[25];
  assign o[12865] = i[25];
  assign o[12866] = i[25];
  assign o[12867] = i[25];
  assign o[12868] = i[25];
  assign o[12869] = i[25];
  assign o[12870] = i[25];
  assign o[12871] = i[25];
  assign o[12872] = i[25];
  assign o[12873] = i[25];
  assign o[12874] = i[25];
  assign o[12875] = i[25];
  assign o[12876] = i[25];
  assign o[12877] = i[25];
  assign o[12878] = i[25];
  assign o[12879] = i[25];
  assign o[12880] = i[25];
  assign o[12881] = i[25];
  assign o[12882] = i[25];
  assign o[12883] = i[25];
  assign o[12884] = i[25];
  assign o[12885] = i[25];
  assign o[12886] = i[25];
  assign o[12887] = i[25];
  assign o[12888] = i[25];
  assign o[12889] = i[25];
  assign o[12890] = i[25];
  assign o[12891] = i[25];
  assign o[12892] = i[25];
  assign o[12893] = i[25];
  assign o[12894] = i[25];
  assign o[12895] = i[25];
  assign o[12896] = i[25];
  assign o[12897] = i[25];
  assign o[12898] = i[25];
  assign o[12899] = i[25];
  assign o[12900] = i[25];
  assign o[12901] = i[25];
  assign o[12902] = i[25];
  assign o[12903] = i[25];
  assign o[12904] = i[25];
  assign o[12905] = i[25];
  assign o[12906] = i[25];
  assign o[12907] = i[25];
  assign o[12908] = i[25];
  assign o[12909] = i[25];
  assign o[12910] = i[25];
  assign o[12911] = i[25];
  assign o[12912] = i[25];
  assign o[12913] = i[25];
  assign o[12914] = i[25];
  assign o[12915] = i[25];
  assign o[12916] = i[25];
  assign o[12917] = i[25];
  assign o[12918] = i[25];
  assign o[12919] = i[25];
  assign o[12920] = i[25];
  assign o[12921] = i[25];
  assign o[12922] = i[25];
  assign o[12923] = i[25];
  assign o[12924] = i[25];
  assign o[12925] = i[25];
  assign o[12926] = i[25];
  assign o[12927] = i[25];
  assign o[12928] = i[25];
  assign o[12929] = i[25];
  assign o[12930] = i[25];
  assign o[12931] = i[25];
  assign o[12932] = i[25];
  assign o[12933] = i[25];
  assign o[12934] = i[25];
  assign o[12935] = i[25];
  assign o[12936] = i[25];
  assign o[12937] = i[25];
  assign o[12938] = i[25];
  assign o[12939] = i[25];
  assign o[12940] = i[25];
  assign o[12941] = i[25];
  assign o[12942] = i[25];
  assign o[12943] = i[25];
  assign o[12944] = i[25];
  assign o[12945] = i[25];
  assign o[12946] = i[25];
  assign o[12947] = i[25];
  assign o[12948] = i[25];
  assign o[12949] = i[25];
  assign o[12950] = i[25];
  assign o[12951] = i[25];
  assign o[12952] = i[25];
  assign o[12953] = i[25];
  assign o[12954] = i[25];
  assign o[12955] = i[25];
  assign o[12956] = i[25];
  assign o[12957] = i[25];
  assign o[12958] = i[25];
  assign o[12959] = i[25];
  assign o[12960] = i[25];
  assign o[12961] = i[25];
  assign o[12962] = i[25];
  assign o[12963] = i[25];
  assign o[12964] = i[25];
  assign o[12965] = i[25];
  assign o[12966] = i[25];
  assign o[12967] = i[25];
  assign o[12968] = i[25];
  assign o[12969] = i[25];
  assign o[12970] = i[25];
  assign o[12971] = i[25];
  assign o[12972] = i[25];
  assign o[12973] = i[25];
  assign o[12974] = i[25];
  assign o[12975] = i[25];
  assign o[12976] = i[25];
  assign o[12977] = i[25];
  assign o[12978] = i[25];
  assign o[12979] = i[25];
  assign o[12980] = i[25];
  assign o[12981] = i[25];
  assign o[12982] = i[25];
  assign o[12983] = i[25];
  assign o[12984] = i[25];
  assign o[12985] = i[25];
  assign o[12986] = i[25];
  assign o[12987] = i[25];
  assign o[12988] = i[25];
  assign o[12989] = i[25];
  assign o[12990] = i[25];
  assign o[12991] = i[25];
  assign o[12992] = i[25];
  assign o[12993] = i[25];
  assign o[12994] = i[25];
  assign o[12995] = i[25];
  assign o[12996] = i[25];
  assign o[12997] = i[25];
  assign o[12998] = i[25];
  assign o[12999] = i[25];
  assign o[13000] = i[25];
  assign o[13001] = i[25];
  assign o[13002] = i[25];
  assign o[13003] = i[25];
  assign o[13004] = i[25];
  assign o[13005] = i[25];
  assign o[13006] = i[25];
  assign o[13007] = i[25];
  assign o[13008] = i[25];
  assign o[13009] = i[25];
  assign o[13010] = i[25];
  assign o[13011] = i[25];
  assign o[13012] = i[25];
  assign o[13013] = i[25];
  assign o[13014] = i[25];
  assign o[13015] = i[25];
  assign o[13016] = i[25];
  assign o[13017] = i[25];
  assign o[13018] = i[25];
  assign o[13019] = i[25];
  assign o[13020] = i[25];
  assign o[13021] = i[25];
  assign o[13022] = i[25];
  assign o[13023] = i[25];
  assign o[13024] = i[25];
  assign o[13025] = i[25];
  assign o[13026] = i[25];
  assign o[13027] = i[25];
  assign o[13028] = i[25];
  assign o[13029] = i[25];
  assign o[13030] = i[25];
  assign o[13031] = i[25];
  assign o[13032] = i[25];
  assign o[13033] = i[25];
  assign o[13034] = i[25];
  assign o[13035] = i[25];
  assign o[13036] = i[25];
  assign o[13037] = i[25];
  assign o[13038] = i[25];
  assign o[13039] = i[25];
  assign o[13040] = i[25];
  assign o[13041] = i[25];
  assign o[13042] = i[25];
  assign o[13043] = i[25];
  assign o[13044] = i[25];
  assign o[13045] = i[25];
  assign o[13046] = i[25];
  assign o[13047] = i[25];
  assign o[13048] = i[25];
  assign o[13049] = i[25];
  assign o[13050] = i[25];
  assign o[13051] = i[25];
  assign o[13052] = i[25];
  assign o[13053] = i[25];
  assign o[13054] = i[25];
  assign o[13055] = i[25];
  assign o[13056] = i[25];
  assign o[13057] = i[25];
  assign o[13058] = i[25];
  assign o[13059] = i[25];
  assign o[13060] = i[25];
  assign o[13061] = i[25];
  assign o[13062] = i[25];
  assign o[13063] = i[25];
  assign o[13064] = i[25];
  assign o[13065] = i[25];
  assign o[13066] = i[25];
  assign o[13067] = i[25];
  assign o[13068] = i[25];
  assign o[13069] = i[25];
  assign o[13070] = i[25];
  assign o[13071] = i[25];
  assign o[13072] = i[25];
  assign o[13073] = i[25];
  assign o[13074] = i[25];
  assign o[13075] = i[25];
  assign o[13076] = i[25];
  assign o[13077] = i[25];
  assign o[13078] = i[25];
  assign o[13079] = i[25];
  assign o[13080] = i[25];
  assign o[13081] = i[25];
  assign o[13082] = i[25];
  assign o[13083] = i[25];
  assign o[13084] = i[25];
  assign o[13085] = i[25];
  assign o[13086] = i[25];
  assign o[13087] = i[25];
  assign o[13088] = i[25];
  assign o[13089] = i[25];
  assign o[13090] = i[25];
  assign o[13091] = i[25];
  assign o[13092] = i[25];
  assign o[13093] = i[25];
  assign o[13094] = i[25];
  assign o[13095] = i[25];
  assign o[13096] = i[25];
  assign o[13097] = i[25];
  assign o[13098] = i[25];
  assign o[13099] = i[25];
  assign o[13100] = i[25];
  assign o[13101] = i[25];
  assign o[13102] = i[25];
  assign o[13103] = i[25];
  assign o[13104] = i[25];
  assign o[13105] = i[25];
  assign o[13106] = i[25];
  assign o[13107] = i[25];
  assign o[13108] = i[25];
  assign o[13109] = i[25];
  assign o[13110] = i[25];
  assign o[13111] = i[25];
  assign o[13112] = i[25];
  assign o[13113] = i[25];
  assign o[13114] = i[25];
  assign o[13115] = i[25];
  assign o[13116] = i[25];
  assign o[13117] = i[25];
  assign o[13118] = i[25];
  assign o[13119] = i[25];
  assign o[13120] = i[25];
  assign o[13121] = i[25];
  assign o[13122] = i[25];
  assign o[13123] = i[25];
  assign o[13124] = i[25];
  assign o[13125] = i[25];
  assign o[13126] = i[25];
  assign o[13127] = i[25];
  assign o[13128] = i[25];
  assign o[13129] = i[25];
  assign o[13130] = i[25];
  assign o[13131] = i[25];
  assign o[13132] = i[25];
  assign o[13133] = i[25];
  assign o[13134] = i[25];
  assign o[13135] = i[25];
  assign o[13136] = i[25];
  assign o[13137] = i[25];
  assign o[13138] = i[25];
  assign o[13139] = i[25];
  assign o[13140] = i[25];
  assign o[13141] = i[25];
  assign o[13142] = i[25];
  assign o[13143] = i[25];
  assign o[13144] = i[25];
  assign o[13145] = i[25];
  assign o[13146] = i[25];
  assign o[13147] = i[25];
  assign o[13148] = i[25];
  assign o[13149] = i[25];
  assign o[13150] = i[25];
  assign o[13151] = i[25];
  assign o[13152] = i[25];
  assign o[13153] = i[25];
  assign o[13154] = i[25];
  assign o[13155] = i[25];
  assign o[13156] = i[25];
  assign o[13157] = i[25];
  assign o[13158] = i[25];
  assign o[13159] = i[25];
  assign o[13160] = i[25];
  assign o[13161] = i[25];
  assign o[13162] = i[25];
  assign o[13163] = i[25];
  assign o[13164] = i[25];
  assign o[13165] = i[25];
  assign o[13166] = i[25];
  assign o[13167] = i[25];
  assign o[13168] = i[25];
  assign o[13169] = i[25];
  assign o[13170] = i[25];
  assign o[13171] = i[25];
  assign o[13172] = i[25];
  assign o[13173] = i[25];
  assign o[13174] = i[25];
  assign o[13175] = i[25];
  assign o[13176] = i[25];
  assign o[13177] = i[25];
  assign o[13178] = i[25];
  assign o[13179] = i[25];
  assign o[13180] = i[25];
  assign o[13181] = i[25];
  assign o[13182] = i[25];
  assign o[13183] = i[25];
  assign o[13184] = i[25];
  assign o[13185] = i[25];
  assign o[13186] = i[25];
  assign o[13187] = i[25];
  assign o[13188] = i[25];
  assign o[13189] = i[25];
  assign o[13190] = i[25];
  assign o[13191] = i[25];
  assign o[13192] = i[25];
  assign o[13193] = i[25];
  assign o[13194] = i[25];
  assign o[13195] = i[25];
  assign o[13196] = i[25];
  assign o[13197] = i[25];
  assign o[13198] = i[25];
  assign o[13199] = i[25];
  assign o[13200] = i[25];
  assign o[13201] = i[25];
  assign o[13202] = i[25];
  assign o[13203] = i[25];
  assign o[13204] = i[25];
  assign o[13205] = i[25];
  assign o[13206] = i[25];
  assign o[13207] = i[25];
  assign o[13208] = i[25];
  assign o[13209] = i[25];
  assign o[13210] = i[25];
  assign o[13211] = i[25];
  assign o[13212] = i[25];
  assign o[13213] = i[25];
  assign o[13214] = i[25];
  assign o[13215] = i[25];
  assign o[13216] = i[25];
  assign o[13217] = i[25];
  assign o[13218] = i[25];
  assign o[13219] = i[25];
  assign o[13220] = i[25];
  assign o[13221] = i[25];
  assign o[13222] = i[25];
  assign o[13223] = i[25];
  assign o[13224] = i[25];
  assign o[13225] = i[25];
  assign o[13226] = i[25];
  assign o[13227] = i[25];
  assign o[13228] = i[25];
  assign o[13229] = i[25];
  assign o[13230] = i[25];
  assign o[13231] = i[25];
  assign o[13232] = i[25];
  assign o[13233] = i[25];
  assign o[13234] = i[25];
  assign o[13235] = i[25];
  assign o[13236] = i[25];
  assign o[13237] = i[25];
  assign o[13238] = i[25];
  assign o[13239] = i[25];
  assign o[13240] = i[25];
  assign o[13241] = i[25];
  assign o[13242] = i[25];
  assign o[13243] = i[25];
  assign o[13244] = i[25];
  assign o[13245] = i[25];
  assign o[13246] = i[25];
  assign o[13247] = i[25];
  assign o[13248] = i[25];
  assign o[13249] = i[25];
  assign o[13250] = i[25];
  assign o[13251] = i[25];
  assign o[13252] = i[25];
  assign o[13253] = i[25];
  assign o[13254] = i[25];
  assign o[13255] = i[25];
  assign o[13256] = i[25];
  assign o[13257] = i[25];
  assign o[13258] = i[25];
  assign o[13259] = i[25];
  assign o[13260] = i[25];
  assign o[13261] = i[25];
  assign o[13262] = i[25];
  assign o[13263] = i[25];
  assign o[13264] = i[25];
  assign o[13265] = i[25];
  assign o[13266] = i[25];
  assign o[13267] = i[25];
  assign o[13268] = i[25];
  assign o[13269] = i[25];
  assign o[13270] = i[25];
  assign o[13271] = i[25];
  assign o[13272] = i[25];
  assign o[13273] = i[25];
  assign o[13274] = i[25];
  assign o[13275] = i[25];
  assign o[13276] = i[25];
  assign o[13277] = i[25];
  assign o[13278] = i[25];
  assign o[13279] = i[25];
  assign o[13280] = i[25];
  assign o[13281] = i[25];
  assign o[13282] = i[25];
  assign o[13283] = i[25];
  assign o[13284] = i[25];
  assign o[13285] = i[25];
  assign o[13286] = i[25];
  assign o[13287] = i[25];
  assign o[13288] = i[25];
  assign o[13289] = i[25];
  assign o[13290] = i[25];
  assign o[13291] = i[25];
  assign o[13292] = i[25];
  assign o[13293] = i[25];
  assign o[13294] = i[25];
  assign o[13295] = i[25];
  assign o[13296] = i[25];
  assign o[13297] = i[25];
  assign o[13298] = i[25];
  assign o[13299] = i[25];
  assign o[13300] = i[25];
  assign o[13301] = i[25];
  assign o[13302] = i[25];
  assign o[13303] = i[25];
  assign o[13304] = i[25];
  assign o[13305] = i[25];
  assign o[13306] = i[25];
  assign o[13307] = i[25];
  assign o[13308] = i[25];
  assign o[13309] = i[25];
  assign o[13310] = i[25];
  assign o[13311] = i[25];
  assign o[12288] = i[24];
  assign o[12289] = i[24];
  assign o[12290] = i[24];
  assign o[12291] = i[24];
  assign o[12292] = i[24];
  assign o[12293] = i[24];
  assign o[12294] = i[24];
  assign o[12295] = i[24];
  assign o[12296] = i[24];
  assign o[12297] = i[24];
  assign o[12298] = i[24];
  assign o[12299] = i[24];
  assign o[12300] = i[24];
  assign o[12301] = i[24];
  assign o[12302] = i[24];
  assign o[12303] = i[24];
  assign o[12304] = i[24];
  assign o[12305] = i[24];
  assign o[12306] = i[24];
  assign o[12307] = i[24];
  assign o[12308] = i[24];
  assign o[12309] = i[24];
  assign o[12310] = i[24];
  assign o[12311] = i[24];
  assign o[12312] = i[24];
  assign o[12313] = i[24];
  assign o[12314] = i[24];
  assign o[12315] = i[24];
  assign o[12316] = i[24];
  assign o[12317] = i[24];
  assign o[12318] = i[24];
  assign o[12319] = i[24];
  assign o[12320] = i[24];
  assign o[12321] = i[24];
  assign o[12322] = i[24];
  assign o[12323] = i[24];
  assign o[12324] = i[24];
  assign o[12325] = i[24];
  assign o[12326] = i[24];
  assign o[12327] = i[24];
  assign o[12328] = i[24];
  assign o[12329] = i[24];
  assign o[12330] = i[24];
  assign o[12331] = i[24];
  assign o[12332] = i[24];
  assign o[12333] = i[24];
  assign o[12334] = i[24];
  assign o[12335] = i[24];
  assign o[12336] = i[24];
  assign o[12337] = i[24];
  assign o[12338] = i[24];
  assign o[12339] = i[24];
  assign o[12340] = i[24];
  assign o[12341] = i[24];
  assign o[12342] = i[24];
  assign o[12343] = i[24];
  assign o[12344] = i[24];
  assign o[12345] = i[24];
  assign o[12346] = i[24];
  assign o[12347] = i[24];
  assign o[12348] = i[24];
  assign o[12349] = i[24];
  assign o[12350] = i[24];
  assign o[12351] = i[24];
  assign o[12352] = i[24];
  assign o[12353] = i[24];
  assign o[12354] = i[24];
  assign o[12355] = i[24];
  assign o[12356] = i[24];
  assign o[12357] = i[24];
  assign o[12358] = i[24];
  assign o[12359] = i[24];
  assign o[12360] = i[24];
  assign o[12361] = i[24];
  assign o[12362] = i[24];
  assign o[12363] = i[24];
  assign o[12364] = i[24];
  assign o[12365] = i[24];
  assign o[12366] = i[24];
  assign o[12367] = i[24];
  assign o[12368] = i[24];
  assign o[12369] = i[24];
  assign o[12370] = i[24];
  assign o[12371] = i[24];
  assign o[12372] = i[24];
  assign o[12373] = i[24];
  assign o[12374] = i[24];
  assign o[12375] = i[24];
  assign o[12376] = i[24];
  assign o[12377] = i[24];
  assign o[12378] = i[24];
  assign o[12379] = i[24];
  assign o[12380] = i[24];
  assign o[12381] = i[24];
  assign o[12382] = i[24];
  assign o[12383] = i[24];
  assign o[12384] = i[24];
  assign o[12385] = i[24];
  assign o[12386] = i[24];
  assign o[12387] = i[24];
  assign o[12388] = i[24];
  assign o[12389] = i[24];
  assign o[12390] = i[24];
  assign o[12391] = i[24];
  assign o[12392] = i[24];
  assign o[12393] = i[24];
  assign o[12394] = i[24];
  assign o[12395] = i[24];
  assign o[12396] = i[24];
  assign o[12397] = i[24];
  assign o[12398] = i[24];
  assign o[12399] = i[24];
  assign o[12400] = i[24];
  assign o[12401] = i[24];
  assign o[12402] = i[24];
  assign o[12403] = i[24];
  assign o[12404] = i[24];
  assign o[12405] = i[24];
  assign o[12406] = i[24];
  assign o[12407] = i[24];
  assign o[12408] = i[24];
  assign o[12409] = i[24];
  assign o[12410] = i[24];
  assign o[12411] = i[24];
  assign o[12412] = i[24];
  assign o[12413] = i[24];
  assign o[12414] = i[24];
  assign o[12415] = i[24];
  assign o[12416] = i[24];
  assign o[12417] = i[24];
  assign o[12418] = i[24];
  assign o[12419] = i[24];
  assign o[12420] = i[24];
  assign o[12421] = i[24];
  assign o[12422] = i[24];
  assign o[12423] = i[24];
  assign o[12424] = i[24];
  assign o[12425] = i[24];
  assign o[12426] = i[24];
  assign o[12427] = i[24];
  assign o[12428] = i[24];
  assign o[12429] = i[24];
  assign o[12430] = i[24];
  assign o[12431] = i[24];
  assign o[12432] = i[24];
  assign o[12433] = i[24];
  assign o[12434] = i[24];
  assign o[12435] = i[24];
  assign o[12436] = i[24];
  assign o[12437] = i[24];
  assign o[12438] = i[24];
  assign o[12439] = i[24];
  assign o[12440] = i[24];
  assign o[12441] = i[24];
  assign o[12442] = i[24];
  assign o[12443] = i[24];
  assign o[12444] = i[24];
  assign o[12445] = i[24];
  assign o[12446] = i[24];
  assign o[12447] = i[24];
  assign o[12448] = i[24];
  assign o[12449] = i[24];
  assign o[12450] = i[24];
  assign o[12451] = i[24];
  assign o[12452] = i[24];
  assign o[12453] = i[24];
  assign o[12454] = i[24];
  assign o[12455] = i[24];
  assign o[12456] = i[24];
  assign o[12457] = i[24];
  assign o[12458] = i[24];
  assign o[12459] = i[24];
  assign o[12460] = i[24];
  assign o[12461] = i[24];
  assign o[12462] = i[24];
  assign o[12463] = i[24];
  assign o[12464] = i[24];
  assign o[12465] = i[24];
  assign o[12466] = i[24];
  assign o[12467] = i[24];
  assign o[12468] = i[24];
  assign o[12469] = i[24];
  assign o[12470] = i[24];
  assign o[12471] = i[24];
  assign o[12472] = i[24];
  assign o[12473] = i[24];
  assign o[12474] = i[24];
  assign o[12475] = i[24];
  assign o[12476] = i[24];
  assign o[12477] = i[24];
  assign o[12478] = i[24];
  assign o[12479] = i[24];
  assign o[12480] = i[24];
  assign o[12481] = i[24];
  assign o[12482] = i[24];
  assign o[12483] = i[24];
  assign o[12484] = i[24];
  assign o[12485] = i[24];
  assign o[12486] = i[24];
  assign o[12487] = i[24];
  assign o[12488] = i[24];
  assign o[12489] = i[24];
  assign o[12490] = i[24];
  assign o[12491] = i[24];
  assign o[12492] = i[24];
  assign o[12493] = i[24];
  assign o[12494] = i[24];
  assign o[12495] = i[24];
  assign o[12496] = i[24];
  assign o[12497] = i[24];
  assign o[12498] = i[24];
  assign o[12499] = i[24];
  assign o[12500] = i[24];
  assign o[12501] = i[24];
  assign o[12502] = i[24];
  assign o[12503] = i[24];
  assign o[12504] = i[24];
  assign o[12505] = i[24];
  assign o[12506] = i[24];
  assign o[12507] = i[24];
  assign o[12508] = i[24];
  assign o[12509] = i[24];
  assign o[12510] = i[24];
  assign o[12511] = i[24];
  assign o[12512] = i[24];
  assign o[12513] = i[24];
  assign o[12514] = i[24];
  assign o[12515] = i[24];
  assign o[12516] = i[24];
  assign o[12517] = i[24];
  assign o[12518] = i[24];
  assign o[12519] = i[24];
  assign o[12520] = i[24];
  assign o[12521] = i[24];
  assign o[12522] = i[24];
  assign o[12523] = i[24];
  assign o[12524] = i[24];
  assign o[12525] = i[24];
  assign o[12526] = i[24];
  assign o[12527] = i[24];
  assign o[12528] = i[24];
  assign o[12529] = i[24];
  assign o[12530] = i[24];
  assign o[12531] = i[24];
  assign o[12532] = i[24];
  assign o[12533] = i[24];
  assign o[12534] = i[24];
  assign o[12535] = i[24];
  assign o[12536] = i[24];
  assign o[12537] = i[24];
  assign o[12538] = i[24];
  assign o[12539] = i[24];
  assign o[12540] = i[24];
  assign o[12541] = i[24];
  assign o[12542] = i[24];
  assign o[12543] = i[24];
  assign o[12544] = i[24];
  assign o[12545] = i[24];
  assign o[12546] = i[24];
  assign o[12547] = i[24];
  assign o[12548] = i[24];
  assign o[12549] = i[24];
  assign o[12550] = i[24];
  assign o[12551] = i[24];
  assign o[12552] = i[24];
  assign o[12553] = i[24];
  assign o[12554] = i[24];
  assign o[12555] = i[24];
  assign o[12556] = i[24];
  assign o[12557] = i[24];
  assign o[12558] = i[24];
  assign o[12559] = i[24];
  assign o[12560] = i[24];
  assign o[12561] = i[24];
  assign o[12562] = i[24];
  assign o[12563] = i[24];
  assign o[12564] = i[24];
  assign o[12565] = i[24];
  assign o[12566] = i[24];
  assign o[12567] = i[24];
  assign o[12568] = i[24];
  assign o[12569] = i[24];
  assign o[12570] = i[24];
  assign o[12571] = i[24];
  assign o[12572] = i[24];
  assign o[12573] = i[24];
  assign o[12574] = i[24];
  assign o[12575] = i[24];
  assign o[12576] = i[24];
  assign o[12577] = i[24];
  assign o[12578] = i[24];
  assign o[12579] = i[24];
  assign o[12580] = i[24];
  assign o[12581] = i[24];
  assign o[12582] = i[24];
  assign o[12583] = i[24];
  assign o[12584] = i[24];
  assign o[12585] = i[24];
  assign o[12586] = i[24];
  assign o[12587] = i[24];
  assign o[12588] = i[24];
  assign o[12589] = i[24];
  assign o[12590] = i[24];
  assign o[12591] = i[24];
  assign o[12592] = i[24];
  assign o[12593] = i[24];
  assign o[12594] = i[24];
  assign o[12595] = i[24];
  assign o[12596] = i[24];
  assign o[12597] = i[24];
  assign o[12598] = i[24];
  assign o[12599] = i[24];
  assign o[12600] = i[24];
  assign o[12601] = i[24];
  assign o[12602] = i[24];
  assign o[12603] = i[24];
  assign o[12604] = i[24];
  assign o[12605] = i[24];
  assign o[12606] = i[24];
  assign o[12607] = i[24];
  assign o[12608] = i[24];
  assign o[12609] = i[24];
  assign o[12610] = i[24];
  assign o[12611] = i[24];
  assign o[12612] = i[24];
  assign o[12613] = i[24];
  assign o[12614] = i[24];
  assign o[12615] = i[24];
  assign o[12616] = i[24];
  assign o[12617] = i[24];
  assign o[12618] = i[24];
  assign o[12619] = i[24];
  assign o[12620] = i[24];
  assign o[12621] = i[24];
  assign o[12622] = i[24];
  assign o[12623] = i[24];
  assign o[12624] = i[24];
  assign o[12625] = i[24];
  assign o[12626] = i[24];
  assign o[12627] = i[24];
  assign o[12628] = i[24];
  assign o[12629] = i[24];
  assign o[12630] = i[24];
  assign o[12631] = i[24];
  assign o[12632] = i[24];
  assign o[12633] = i[24];
  assign o[12634] = i[24];
  assign o[12635] = i[24];
  assign o[12636] = i[24];
  assign o[12637] = i[24];
  assign o[12638] = i[24];
  assign o[12639] = i[24];
  assign o[12640] = i[24];
  assign o[12641] = i[24];
  assign o[12642] = i[24];
  assign o[12643] = i[24];
  assign o[12644] = i[24];
  assign o[12645] = i[24];
  assign o[12646] = i[24];
  assign o[12647] = i[24];
  assign o[12648] = i[24];
  assign o[12649] = i[24];
  assign o[12650] = i[24];
  assign o[12651] = i[24];
  assign o[12652] = i[24];
  assign o[12653] = i[24];
  assign o[12654] = i[24];
  assign o[12655] = i[24];
  assign o[12656] = i[24];
  assign o[12657] = i[24];
  assign o[12658] = i[24];
  assign o[12659] = i[24];
  assign o[12660] = i[24];
  assign o[12661] = i[24];
  assign o[12662] = i[24];
  assign o[12663] = i[24];
  assign o[12664] = i[24];
  assign o[12665] = i[24];
  assign o[12666] = i[24];
  assign o[12667] = i[24];
  assign o[12668] = i[24];
  assign o[12669] = i[24];
  assign o[12670] = i[24];
  assign o[12671] = i[24];
  assign o[12672] = i[24];
  assign o[12673] = i[24];
  assign o[12674] = i[24];
  assign o[12675] = i[24];
  assign o[12676] = i[24];
  assign o[12677] = i[24];
  assign o[12678] = i[24];
  assign o[12679] = i[24];
  assign o[12680] = i[24];
  assign o[12681] = i[24];
  assign o[12682] = i[24];
  assign o[12683] = i[24];
  assign o[12684] = i[24];
  assign o[12685] = i[24];
  assign o[12686] = i[24];
  assign o[12687] = i[24];
  assign o[12688] = i[24];
  assign o[12689] = i[24];
  assign o[12690] = i[24];
  assign o[12691] = i[24];
  assign o[12692] = i[24];
  assign o[12693] = i[24];
  assign o[12694] = i[24];
  assign o[12695] = i[24];
  assign o[12696] = i[24];
  assign o[12697] = i[24];
  assign o[12698] = i[24];
  assign o[12699] = i[24];
  assign o[12700] = i[24];
  assign o[12701] = i[24];
  assign o[12702] = i[24];
  assign o[12703] = i[24];
  assign o[12704] = i[24];
  assign o[12705] = i[24];
  assign o[12706] = i[24];
  assign o[12707] = i[24];
  assign o[12708] = i[24];
  assign o[12709] = i[24];
  assign o[12710] = i[24];
  assign o[12711] = i[24];
  assign o[12712] = i[24];
  assign o[12713] = i[24];
  assign o[12714] = i[24];
  assign o[12715] = i[24];
  assign o[12716] = i[24];
  assign o[12717] = i[24];
  assign o[12718] = i[24];
  assign o[12719] = i[24];
  assign o[12720] = i[24];
  assign o[12721] = i[24];
  assign o[12722] = i[24];
  assign o[12723] = i[24];
  assign o[12724] = i[24];
  assign o[12725] = i[24];
  assign o[12726] = i[24];
  assign o[12727] = i[24];
  assign o[12728] = i[24];
  assign o[12729] = i[24];
  assign o[12730] = i[24];
  assign o[12731] = i[24];
  assign o[12732] = i[24];
  assign o[12733] = i[24];
  assign o[12734] = i[24];
  assign o[12735] = i[24];
  assign o[12736] = i[24];
  assign o[12737] = i[24];
  assign o[12738] = i[24];
  assign o[12739] = i[24];
  assign o[12740] = i[24];
  assign o[12741] = i[24];
  assign o[12742] = i[24];
  assign o[12743] = i[24];
  assign o[12744] = i[24];
  assign o[12745] = i[24];
  assign o[12746] = i[24];
  assign o[12747] = i[24];
  assign o[12748] = i[24];
  assign o[12749] = i[24];
  assign o[12750] = i[24];
  assign o[12751] = i[24];
  assign o[12752] = i[24];
  assign o[12753] = i[24];
  assign o[12754] = i[24];
  assign o[12755] = i[24];
  assign o[12756] = i[24];
  assign o[12757] = i[24];
  assign o[12758] = i[24];
  assign o[12759] = i[24];
  assign o[12760] = i[24];
  assign o[12761] = i[24];
  assign o[12762] = i[24];
  assign o[12763] = i[24];
  assign o[12764] = i[24];
  assign o[12765] = i[24];
  assign o[12766] = i[24];
  assign o[12767] = i[24];
  assign o[12768] = i[24];
  assign o[12769] = i[24];
  assign o[12770] = i[24];
  assign o[12771] = i[24];
  assign o[12772] = i[24];
  assign o[12773] = i[24];
  assign o[12774] = i[24];
  assign o[12775] = i[24];
  assign o[12776] = i[24];
  assign o[12777] = i[24];
  assign o[12778] = i[24];
  assign o[12779] = i[24];
  assign o[12780] = i[24];
  assign o[12781] = i[24];
  assign o[12782] = i[24];
  assign o[12783] = i[24];
  assign o[12784] = i[24];
  assign o[12785] = i[24];
  assign o[12786] = i[24];
  assign o[12787] = i[24];
  assign o[12788] = i[24];
  assign o[12789] = i[24];
  assign o[12790] = i[24];
  assign o[12791] = i[24];
  assign o[12792] = i[24];
  assign o[12793] = i[24];
  assign o[12794] = i[24];
  assign o[12795] = i[24];
  assign o[12796] = i[24];
  assign o[12797] = i[24];
  assign o[12798] = i[24];
  assign o[12799] = i[24];
  assign o[11776] = i[23];
  assign o[11777] = i[23];
  assign o[11778] = i[23];
  assign o[11779] = i[23];
  assign o[11780] = i[23];
  assign o[11781] = i[23];
  assign o[11782] = i[23];
  assign o[11783] = i[23];
  assign o[11784] = i[23];
  assign o[11785] = i[23];
  assign o[11786] = i[23];
  assign o[11787] = i[23];
  assign o[11788] = i[23];
  assign o[11789] = i[23];
  assign o[11790] = i[23];
  assign o[11791] = i[23];
  assign o[11792] = i[23];
  assign o[11793] = i[23];
  assign o[11794] = i[23];
  assign o[11795] = i[23];
  assign o[11796] = i[23];
  assign o[11797] = i[23];
  assign o[11798] = i[23];
  assign o[11799] = i[23];
  assign o[11800] = i[23];
  assign o[11801] = i[23];
  assign o[11802] = i[23];
  assign o[11803] = i[23];
  assign o[11804] = i[23];
  assign o[11805] = i[23];
  assign o[11806] = i[23];
  assign o[11807] = i[23];
  assign o[11808] = i[23];
  assign o[11809] = i[23];
  assign o[11810] = i[23];
  assign o[11811] = i[23];
  assign o[11812] = i[23];
  assign o[11813] = i[23];
  assign o[11814] = i[23];
  assign o[11815] = i[23];
  assign o[11816] = i[23];
  assign o[11817] = i[23];
  assign o[11818] = i[23];
  assign o[11819] = i[23];
  assign o[11820] = i[23];
  assign o[11821] = i[23];
  assign o[11822] = i[23];
  assign o[11823] = i[23];
  assign o[11824] = i[23];
  assign o[11825] = i[23];
  assign o[11826] = i[23];
  assign o[11827] = i[23];
  assign o[11828] = i[23];
  assign o[11829] = i[23];
  assign o[11830] = i[23];
  assign o[11831] = i[23];
  assign o[11832] = i[23];
  assign o[11833] = i[23];
  assign o[11834] = i[23];
  assign o[11835] = i[23];
  assign o[11836] = i[23];
  assign o[11837] = i[23];
  assign o[11838] = i[23];
  assign o[11839] = i[23];
  assign o[11840] = i[23];
  assign o[11841] = i[23];
  assign o[11842] = i[23];
  assign o[11843] = i[23];
  assign o[11844] = i[23];
  assign o[11845] = i[23];
  assign o[11846] = i[23];
  assign o[11847] = i[23];
  assign o[11848] = i[23];
  assign o[11849] = i[23];
  assign o[11850] = i[23];
  assign o[11851] = i[23];
  assign o[11852] = i[23];
  assign o[11853] = i[23];
  assign o[11854] = i[23];
  assign o[11855] = i[23];
  assign o[11856] = i[23];
  assign o[11857] = i[23];
  assign o[11858] = i[23];
  assign o[11859] = i[23];
  assign o[11860] = i[23];
  assign o[11861] = i[23];
  assign o[11862] = i[23];
  assign o[11863] = i[23];
  assign o[11864] = i[23];
  assign o[11865] = i[23];
  assign o[11866] = i[23];
  assign o[11867] = i[23];
  assign o[11868] = i[23];
  assign o[11869] = i[23];
  assign o[11870] = i[23];
  assign o[11871] = i[23];
  assign o[11872] = i[23];
  assign o[11873] = i[23];
  assign o[11874] = i[23];
  assign o[11875] = i[23];
  assign o[11876] = i[23];
  assign o[11877] = i[23];
  assign o[11878] = i[23];
  assign o[11879] = i[23];
  assign o[11880] = i[23];
  assign o[11881] = i[23];
  assign o[11882] = i[23];
  assign o[11883] = i[23];
  assign o[11884] = i[23];
  assign o[11885] = i[23];
  assign o[11886] = i[23];
  assign o[11887] = i[23];
  assign o[11888] = i[23];
  assign o[11889] = i[23];
  assign o[11890] = i[23];
  assign o[11891] = i[23];
  assign o[11892] = i[23];
  assign o[11893] = i[23];
  assign o[11894] = i[23];
  assign o[11895] = i[23];
  assign o[11896] = i[23];
  assign o[11897] = i[23];
  assign o[11898] = i[23];
  assign o[11899] = i[23];
  assign o[11900] = i[23];
  assign o[11901] = i[23];
  assign o[11902] = i[23];
  assign o[11903] = i[23];
  assign o[11904] = i[23];
  assign o[11905] = i[23];
  assign o[11906] = i[23];
  assign o[11907] = i[23];
  assign o[11908] = i[23];
  assign o[11909] = i[23];
  assign o[11910] = i[23];
  assign o[11911] = i[23];
  assign o[11912] = i[23];
  assign o[11913] = i[23];
  assign o[11914] = i[23];
  assign o[11915] = i[23];
  assign o[11916] = i[23];
  assign o[11917] = i[23];
  assign o[11918] = i[23];
  assign o[11919] = i[23];
  assign o[11920] = i[23];
  assign o[11921] = i[23];
  assign o[11922] = i[23];
  assign o[11923] = i[23];
  assign o[11924] = i[23];
  assign o[11925] = i[23];
  assign o[11926] = i[23];
  assign o[11927] = i[23];
  assign o[11928] = i[23];
  assign o[11929] = i[23];
  assign o[11930] = i[23];
  assign o[11931] = i[23];
  assign o[11932] = i[23];
  assign o[11933] = i[23];
  assign o[11934] = i[23];
  assign o[11935] = i[23];
  assign o[11936] = i[23];
  assign o[11937] = i[23];
  assign o[11938] = i[23];
  assign o[11939] = i[23];
  assign o[11940] = i[23];
  assign o[11941] = i[23];
  assign o[11942] = i[23];
  assign o[11943] = i[23];
  assign o[11944] = i[23];
  assign o[11945] = i[23];
  assign o[11946] = i[23];
  assign o[11947] = i[23];
  assign o[11948] = i[23];
  assign o[11949] = i[23];
  assign o[11950] = i[23];
  assign o[11951] = i[23];
  assign o[11952] = i[23];
  assign o[11953] = i[23];
  assign o[11954] = i[23];
  assign o[11955] = i[23];
  assign o[11956] = i[23];
  assign o[11957] = i[23];
  assign o[11958] = i[23];
  assign o[11959] = i[23];
  assign o[11960] = i[23];
  assign o[11961] = i[23];
  assign o[11962] = i[23];
  assign o[11963] = i[23];
  assign o[11964] = i[23];
  assign o[11965] = i[23];
  assign o[11966] = i[23];
  assign o[11967] = i[23];
  assign o[11968] = i[23];
  assign o[11969] = i[23];
  assign o[11970] = i[23];
  assign o[11971] = i[23];
  assign o[11972] = i[23];
  assign o[11973] = i[23];
  assign o[11974] = i[23];
  assign o[11975] = i[23];
  assign o[11976] = i[23];
  assign o[11977] = i[23];
  assign o[11978] = i[23];
  assign o[11979] = i[23];
  assign o[11980] = i[23];
  assign o[11981] = i[23];
  assign o[11982] = i[23];
  assign o[11983] = i[23];
  assign o[11984] = i[23];
  assign o[11985] = i[23];
  assign o[11986] = i[23];
  assign o[11987] = i[23];
  assign o[11988] = i[23];
  assign o[11989] = i[23];
  assign o[11990] = i[23];
  assign o[11991] = i[23];
  assign o[11992] = i[23];
  assign o[11993] = i[23];
  assign o[11994] = i[23];
  assign o[11995] = i[23];
  assign o[11996] = i[23];
  assign o[11997] = i[23];
  assign o[11998] = i[23];
  assign o[11999] = i[23];
  assign o[12000] = i[23];
  assign o[12001] = i[23];
  assign o[12002] = i[23];
  assign o[12003] = i[23];
  assign o[12004] = i[23];
  assign o[12005] = i[23];
  assign o[12006] = i[23];
  assign o[12007] = i[23];
  assign o[12008] = i[23];
  assign o[12009] = i[23];
  assign o[12010] = i[23];
  assign o[12011] = i[23];
  assign o[12012] = i[23];
  assign o[12013] = i[23];
  assign o[12014] = i[23];
  assign o[12015] = i[23];
  assign o[12016] = i[23];
  assign o[12017] = i[23];
  assign o[12018] = i[23];
  assign o[12019] = i[23];
  assign o[12020] = i[23];
  assign o[12021] = i[23];
  assign o[12022] = i[23];
  assign o[12023] = i[23];
  assign o[12024] = i[23];
  assign o[12025] = i[23];
  assign o[12026] = i[23];
  assign o[12027] = i[23];
  assign o[12028] = i[23];
  assign o[12029] = i[23];
  assign o[12030] = i[23];
  assign o[12031] = i[23];
  assign o[12032] = i[23];
  assign o[12033] = i[23];
  assign o[12034] = i[23];
  assign o[12035] = i[23];
  assign o[12036] = i[23];
  assign o[12037] = i[23];
  assign o[12038] = i[23];
  assign o[12039] = i[23];
  assign o[12040] = i[23];
  assign o[12041] = i[23];
  assign o[12042] = i[23];
  assign o[12043] = i[23];
  assign o[12044] = i[23];
  assign o[12045] = i[23];
  assign o[12046] = i[23];
  assign o[12047] = i[23];
  assign o[12048] = i[23];
  assign o[12049] = i[23];
  assign o[12050] = i[23];
  assign o[12051] = i[23];
  assign o[12052] = i[23];
  assign o[12053] = i[23];
  assign o[12054] = i[23];
  assign o[12055] = i[23];
  assign o[12056] = i[23];
  assign o[12057] = i[23];
  assign o[12058] = i[23];
  assign o[12059] = i[23];
  assign o[12060] = i[23];
  assign o[12061] = i[23];
  assign o[12062] = i[23];
  assign o[12063] = i[23];
  assign o[12064] = i[23];
  assign o[12065] = i[23];
  assign o[12066] = i[23];
  assign o[12067] = i[23];
  assign o[12068] = i[23];
  assign o[12069] = i[23];
  assign o[12070] = i[23];
  assign o[12071] = i[23];
  assign o[12072] = i[23];
  assign o[12073] = i[23];
  assign o[12074] = i[23];
  assign o[12075] = i[23];
  assign o[12076] = i[23];
  assign o[12077] = i[23];
  assign o[12078] = i[23];
  assign o[12079] = i[23];
  assign o[12080] = i[23];
  assign o[12081] = i[23];
  assign o[12082] = i[23];
  assign o[12083] = i[23];
  assign o[12084] = i[23];
  assign o[12085] = i[23];
  assign o[12086] = i[23];
  assign o[12087] = i[23];
  assign o[12088] = i[23];
  assign o[12089] = i[23];
  assign o[12090] = i[23];
  assign o[12091] = i[23];
  assign o[12092] = i[23];
  assign o[12093] = i[23];
  assign o[12094] = i[23];
  assign o[12095] = i[23];
  assign o[12096] = i[23];
  assign o[12097] = i[23];
  assign o[12098] = i[23];
  assign o[12099] = i[23];
  assign o[12100] = i[23];
  assign o[12101] = i[23];
  assign o[12102] = i[23];
  assign o[12103] = i[23];
  assign o[12104] = i[23];
  assign o[12105] = i[23];
  assign o[12106] = i[23];
  assign o[12107] = i[23];
  assign o[12108] = i[23];
  assign o[12109] = i[23];
  assign o[12110] = i[23];
  assign o[12111] = i[23];
  assign o[12112] = i[23];
  assign o[12113] = i[23];
  assign o[12114] = i[23];
  assign o[12115] = i[23];
  assign o[12116] = i[23];
  assign o[12117] = i[23];
  assign o[12118] = i[23];
  assign o[12119] = i[23];
  assign o[12120] = i[23];
  assign o[12121] = i[23];
  assign o[12122] = i[23];
  assign o[12123] = i[23];
  assign o[12124] = i[23];
  assign o[12125] = i[23];
  assign o[12126] = i[23];
  assign o[12127] = i[23];
  assign o[12128] = i[23];
  assign o[12129] = i[23];
  assign o[12130] = i[23];
  assign o[12131] = i[23];
  assign o[12132] = i[23];
  assign o[12133] = i[23];
  assign o[12134] = i[23];
  assign o[12135] = i[23];
  assign o[12136] = i[23];
  assign o[12137] = i[23];
  assign o[12138] = i[23];
  assign o[12139] = i[23];
  assign o[12140] = i[23];
  assign o[12141] = i[23];
  assign o[12142] = i[23];
  assign o[12143] = i[23];
  assign o[12144] = i[23];
  assign o[12145] = i[23];
  assign o[12146] = i[23];
  assign o[12147] = i[23];
  assign o[12148] = i[23];
  assign o[12149] = i[23];
  assign o[12150] = i[23];
  assign o[12151] = i[23];
  assign o[12152] = i[23];
  assign o[12153] = i[23];
  assign o[12154] = i[23];
  assign o[12155] = i[23];
  assign o[12156] = i[23];
  assign o[12157] = i[23];
  assign o[12158] = i[23];
  assign o[12159] = i[23];
  assign o[12160] = i[23];
  assign o[12161] = i[23];
  assign o[12162] = i[23];
  assign o[12163] = i[23];
  assign o[12164] = i[23];
  assign o[12165] = i[23];
  assign o[12166] = i[23];
  assign o[12167] = i[23];
  assign o[12168] = i[23];
  assign o[12169] = i[23];
  assign o[12170] = i[23];
  assign o[12171] = i[23];
  assign o[12172] = i[23];
  assign o[12173] = i[23];
  assign o[12174] = i[23];
  assign o[12175] = i[23];
  assign o[12176] = i[23];
  assign o[12177] = i[23];
  assign o[12178] = i[23];
  assign o[12179] = i[23];
  assign o[12180] = i[23];
  assign o[12181] = i[23];
  assign o[12182] = i[23];
  assign o[12183] = i[23];
  assign o[12184] = i[23];
  assign o[12185] = i[23];
  assign o[12186] = i[23];
  assign o[12187] = i[23];
  assign o[12188] = i[23];
  assign o[12189] = i[23];
  assign o[12190] = i[23];
  assign o[12191] = i[23];
  assign o[12192] = i[23];
  assign o[12193] = i[23];
  assign o[12194] = i[23];
  assign o[12195] = i[23];
  assign o[12196] = i[23];
  assign o[12197] = i[23];
  assign o[12198] = i[23];
  assign o[12199] = i[23];
  assign o[12200] = i[23];
  assign o[12201] = i[23];
  assign o[12202] = i[23];
  assign o[12203] = i[23];
  assign o[12204] = i[23];
  assign o[12205] = i[23];
  assign o[12206] = i[23];
  assign o[12207] = i[23];
  assign o[12208] = i[23];
  assign o[12209] = i[23];
  assign o[12210] = i[23];
  assign o[12211] = i[23];
  assign o[12212] = i[23];
  assign o[12213] = i[23];
  assign o[12214] = i[23];
  assign o[12215] = i[23];
  assign o[12216] = i[23];
  assign o[12217] = i[23];
  assign o[12218] = i[23];
  assign o[12219] = i[23];
  assign o[12220] = i[23];
  assign o[12221] = i[23];
  assign o[12222] = i[23];
  assign o[12223] = i[23];
  assign o[12224] = i[23];
  assign o[12225] = i[23];
  assign o[12226] = i[23];
  assign o[12227] = i[23];
  assign o[12228] = i[23];
  assign o[12229] = i[23];
  assign o[12230] = i[23];
  assign o[12231] = i[23];
  assign o[12232] = i[23];
  assign o[12233] = i[23];
  assign o[12234] = i[23];
  assign o[12235] = i[23];
  assign o[12236] = i[23];
  assign o[12237] = i[23];
  assign o[12238] = i[23];
  assign o[12239] = i[23];
  assign o[12240] = i[23];
  assign o[12241] = i[23];
  assign o[12242] = i[23];
  assign o[12243] = i[23];
  assign o[12244] = i[23];
  assign o[12245] = i[23];
  assign o[12246] = i[23];
  assign o[12247] = i[23];
  assign o[12248] = i[23];
  assign o[12249] = i[23];
  assign o[12250] = i[23];
  assign o[12251] = i[23];
  assign o[12252] = i[23];
  assign o[12253] = i[23];
  assign o[12254] = i[23];
  assign o[12255] = i[23];
  assign o[12256] = i[23];
  assign o[12257] = i[23];
  assign o[12258] = i[23];
  assign o[12259] = i[23];
  assign o[12260] = i[23];
  assign o[12261] = i[23];
  assign o[12262] = i[23];
  assign o[12263] = i[23];
  assign o[12264] = i[23];
  assign o[12265] = i[23];
  assign o[12266] = i[23];
  assign o[12267] = i[23];
  assign o[12268] = i[23];
  assign o[12269] = i[23];
  assign o[12270] = i[23];
  assign o[12271] = i[23];
  assign o[12272] = i[23];
  assign o[12273] = i[23];
  assign o[12274] = i[23];
  assign o[12275] = i[23];
  assign o[12276] = i[23];
  assign o[12277] = i[23];
  assign o[12278] = i[23];
  assign o[12279] = i[23];
  assign o[12280] = i[23];
  assign o[12281] = i[23];
  assign o[12282] = i[23];
  assign o[12283] = i[23];
  assign o[12284] = i[23];
  assign o[12285] = i[23];
  assign o[12286] = i[23];
  assign o[12287] = i[23];
  assign o[11264] = i[22];
  assign o[11265] = i[22];
  assign o[11266] = i[22];
  assign o[11267] = i[22];
  assign o[11268] = i[22];
  assign o[11269] = i[22];
  assign o[11270] = i[22];
  assign o[11271] = i[22];
  assign o[11272] = i[22];
  assign o[11273] = i[22];
  assign o[11274] = i[22];
  assign o[11275] = i[22];
  assign o[11276] = i[22];
  assign o[11277] = i[22];
  assign o[11278] = i[22];
  assign o[11279] = i[22];
  assign o[11280] = i[22];
  assign o[11281] = i[22];
  assign o[11282] = i[22];
  assign o[11283] = i[22];
  assign o[11284] = i[22];
  assign o[11285] = i[22];
  assign o[11286] = i[22];
  assign o[11287] = i[22];
  assign o[11288] = i[22];
  assign o[11289] = i[22];
  assign o[11290] = i[22];
  assign o[11291] = i[22];
  assign o[11292] = i[22];
  assign o[11293] = i[22];
  assign o[11294] = i[22];
  assign o[11295] = i[22];
  assign o[11296] = i[22];
  assign o[11297] = i[22];
  assign o[11298] = i[22];
  assign o[11299] = i[22];
  assign o[11300] = i[22];
  assign o[11301] = i[22];
  assign o[11302] = i[22];
  assign o[11303] = i[22];
  assign o[11304] = i[22];
  assign o[11305] = i[22];
  assign o[11306] = i[22];
  assign o[11307] = i[22];
  assign o[11308] = i[22];
  assign o[11309] = i[22];
  assign o[11310] = i[22];
  assign o[11311] = i[22];
  assign o[11312] = i[22];
  assign o[11313] = i[22];
  assign o[11314] = i[22];
  assign o[11315] = i[22];
  assign o[11316] = i[22];
  assign o[11317] = i[22];
  assign o[11318] = i[22];
  assign o[11319] = i[22];
  assign o[11320] = i[22];
  assign o[11321] = i[22];
  assign o[11322] = i[22];
  assign o[11323] = i[22];
  assign o[11324] = i[22];
  assign o[11325] = i[22];
  assign o[11326] = i[22];
  assign o[11327] = i[22];
  assign o[11328] = i[22];
  assign o[11329] = i[22];
  assign o[11330] = i[22];
  assign o[11331] = i[22];
  assign o[11332] = i[22];
  assign o[11333] = i[22];
  assign o[11334] = i[22];
  assign o[11335] = i[22];
  assign o[11336] = i[22];
  assign o[11337] = i[22];
  assign o[11338] = i[22];
  assign o[11339] = i[22];
  assign o[11340] = i[22];
  assign o[11341] = i[22];
  assign o[11342] = i[22];
  assign o[11343] = i[22];
  assign o[11344] = i[22];
  assign o[11345] = i[22];
  assign o[11346] = i[22];
  assign o[11347] = i[22];
  assign o[11348] = i[22];
  assign o[11349] = i[22];
  assign o[11350] = i[22];
  assign o[11351] = i[22];
  assign o[11352] = i[22];
  assign o[11353] = i[22];
  assign o[11354] = i[22];
  assign o[11355] = i[22];
  assign o[11356] = i[22];
  assign o[11357] = i[22];
  assign o[11358] = i[22];
  assign o[11359] = i[22];
  assign o[11360] = i[22];
  assign o[11361] = i[22];
  assign o[11362] = i[22];
  assign o[11363] = i[22];
  assign o[11364] = i[22];
  assign o[11365] = i[22];
  assign o[11366] = i[22];
  assign o[11367] = i[22];
  assign o[11368] = i[22];
  assign o[11369] = i[22];
  assign o[11370] = i[22];
  assign o[11371] = i[22];
  assign o[11372] = i[22];
  assign o[11373] = i[22];
  assign o[11374] = i[22];
  assign o[11375] = i[22];
  assign o[11376] = i[22];
  assign o[11377] = i[22];
  assign o[11378] = i[22];
  assign o[11379] = i[22];
  assign o[11380] = i[22];
  assign o[11381] = i[22];
  assign o[11382] = i[22];
  assign o[11383] = i[22];
  assign o[11384] = i[22];
  assign o[11385] = i[22];
  assign o[11386] = i[22];
  assign o[11387] = i[22];
  assign o[11388] = i[22];
  assign o[11389] = i[22];
  assign o[11390] = i[22];
  assign o[11391] = i[22];
  assign o[11392] = i[22];
  assign o[11393] = i[22];
  assign o[11394] = i[22];
  assign o[11395] = i[22];
  assign o[11396] = i[22];
  assign o[11397] = i[22];
  assign o[11398] = i[22];
  assign o[11399] = i[22];
  assign o[11400] = i[22];
  assign o[11401] = i[22];
  assign o[11402] = i[22];
  assign o[11403] = i[22];
  assign o[11404] = i[22];
  assign o[11405] = i[22];
  assign o[11406] = i[22];
  assign o[11407] = i[22];
  assign o[11408] = i[22];
  assign o[11409] = i[22];
  assign o[11410] = i[22];
  assign o[11411] = i[22];
  assign o[11412] = i[22];
  assign o[11413] = i[22];
  assign o[11414] = i[22];
  assign o[11415] = i[22];
  assign o[11416] = i[22];
  assign o[11417] = i[22];
  assign o[11418] = i[22];
  assign o[11419] = i[22];
  assign o[11420] = i[22];
  assign o[11421] = i[22];
  assign o[11422] = i[22];
  assign o[11423] = i[22];
  assign o[11424] = i[22];
  assign o[11425] = i[22];
  assign o[11426] = i[22];
  assign o[11427] = i[22];
  assign o[11428] = i[22];
  assign o[11429] = i[22];
  assign o[11430] = i[22];
  assign o[11431] = i[22];
  assign o[11432] = i[22];
  assign o[11433] = i[22];
  assign o[11434] = i[22];
  assign o[11435] = i[22];
  assign o[11436] = i[22];
  assign o[11437] = i[22];
  assign o[11438] = i[22];
  assign o[11439] = i[22];
  assign o[11440] = i[22];
  assign o[11441] = i[22];
  assign o[11442] = i[22];
  assign o[11443] = i[22];
  assign o[11444] = i[22];
  assign o[11445] = i[22];
  assign o[11446] = i[22];
  assign o[11447] = i[22];
  assign o[11448] = i[22];
  assign o[11449] = i[22];
  assign o[11450] = i[22];
  assign o[11451] = i[22];
  assign o[11452] = i[22];
  assign o[11453] = i[22];
  assign o[11454] = i[22];
  assign o[11455] = i[22];
  assign o[11456] = i[22];
  assign o[11457] = i[22];
  assign o[11458] = i[22];
  assign o[11459] = i[22];
  assign o[11460] = i[22];
  assign o[11461] = i[22];
  assign o[11462] = i[22];
  assign o[11463] = i[22];
  assign o[11464] = i[22];
  assign o[11465] = i[22];
  assign o[11466] = i[22];
  assign o[11467] = i[22];
  assign o[11468] = i[22];
  assign o[11469] = i[22];
  assign o[11470] = i[22];
  assign o[11471] = i[22];
  assign o[11472] = i[22];
  assign o[11473] = i[22];
  assign o[11474] = i[22];
  assign o[11475] = i[22];
  assign o[11476] = i[22];
  assign o[11477] = i[22];
  assign o[11478] = i[22];
  assign o[11479] = i[22];
  assign o[11480] = i[22];
  assign o[11481] = i[22];
  assign o[11482] = i[22];
  assign o[11483] = i[22];
  assign o[11484] = i[22];
  assign o[11485] = i[22];
  assign o[11486] = i[22];
  assign o[11487] = i[22];
  assign o[11488] = i[22];
  assign o[11489] = i[22];
  assign o[11490] = i[22];
  assign o[11491] = i[22];
  assign o[11492] = i[22];
  assign o[11493] = i[22];
  assign o[11494] = i[22];
  assign o[11495] = i[22];
  assign o[11496] = i[22];
  assign o[11497] = i[22];
  assign o[11498] = i[22];
  assign o[11499] = i[22];
  assign o[11500] = i[22];
  assign o[11501] = i[22];
  assign o[11502] = i[22];
  assign o[11503] = i[22];
  assign o[11504] = i[22];
  assign o[11505] = i[22];
  assign o[11506] = i[22];
  assign o[11507] = i[22];
  assign o[11508] = i[22];
  assign o[11509] = i[22];
  assign o[11510] = i[22];
  assign o[11511] = i[22];
  assign o[11512] = i[22];
  assign o[11513] = i[22];
  assign o[11514] = i[22];
  assign o[11515] = i[22];
  assign o[11516] = i[22];
  assign o[11517] = i[22];
  assign o[11518] = i[22];
  assign o[11519] = i[22];
  assign o[11520] = i[22];
  assign o[11521] = i[22];
  assign o[11522] = i[22];
  assign o[11523] = i[22];
  assign o[11524] = i[22];
  assign o[11525] = i[22];
  assign o[11526] = i[22];
  assign o[11527] = i[22];
  assign o[11528] = i[22];
  assign o[11529] = i[22];
  assign o[11530] = i[22];
  assign o[11531] = i[22];
  assign o[11532] = i[22];
  assign o[11533] = i[22];
  assign o[11534] = i[22];
  assign o[11535] = i[22];
  assign o[11536] = i[22];
  assign o[11537] = i[22];
  assign o[11538] = i[22];
  assign o[11539] = i[22];
  assign o[11540] = i[22];
  assign o[11541] = i[22];
  assign o[11542] = i[22];
  assign o[11543] = i[22];
  assign o[11544] = i[22];
  assign o[11545] = i[22];
  assign o[11546] = i[22];
  assign o[11547] = i[22];
  assign o[11548] = i[22];
  assign o[11549] = i[22];
  assign o[11550] = i[22];
  assign o[11551] = i[22];
  assign o[11552] = i[22];
  assign o[11553] = i[22];
  assign o[11554] = i[22];
  assign o[11555] = i[22];
  assign o[11556] = i[22];
  assign o[11557] = i[22];
  assign o[11558] = i[22];
  assign o[11559] = i[22];
  assign o[11560] = i[22];
  assign o[11561] = i[22];
  assign o[11562] = i[22];
  assign o[11563] = i[22];
  assign o[11564] = i[22];
  assign o[11565] = i[22];
  assign o[11566] = i[22];
  assign o[11567] = i[22];
  assign o[11568] = i[22];
  assign o[11569] = i[22];
  assign o[11570] = i[22];
  assign o[11571] = i[22];
  assign o[11572] = i[22];
  assign o[11573] = i[22];
  assign o[11574] = i[22];
  assign o[11575] = i[22];
  assign o[11576] = i[22];
  assign o[11577] = i[22];
  assign o[11578] = i[22];
  assign o[11579] = i[22];
  assign o[11580] = i[22];
  assign o[11581] = i[22];
  assign o[11582] = i[22];
  assign o[11583] = i[22];
  assign o[11584] = i[22];
  assign o[11585] = i[22];
  assign o[11586] = i[22];
  assign o[11587] = i[22];
  assign o[11588] = i[22];
  assign o[11589] = i[22];
  assign o[11590] = i[22];
  assign o[11591] = i[22];
  assign o[11592] = i[22];
  assign o[11593] = i[22];
  assign o[11594] = i[22];
  assign o[11595] = i[22];
  assign o[11596] = i[22];
  assign o[11597] = i[22];
  assign o[11598] = i[22];
  assign o[11599] = i[22];
  assign o[11600] = i[22];
  assign o[11601] = i[22];
  assign o[11602] = i[22];
  assign o[11603] = i[22];
  assign o[11604] = i[22];
  assign o[11605] = i[22];
  assign o[11606] = i[22];
  assign o[11607] = i[22];
  assign o[11608] = i[22];
  assign o[11609] = i[22];
  assign o[11610] = i[22];
  assign o[11611] = i[22];
  assign o[11612] = i[22];
  assign o[11613] = i[22];
  assign o[11614] = i[22];
  assign o[11615] = i[22];
  assign o[11616] = i[22];
  assign o[11617] = i[22];
  assign o[11618] = i[22];
  assign o[11619] = i[22];
  assign o[11620] = i[22];
  assign o[11621] = i[22];
  assign o[11622] = i[22];
  assign o[11623] = i[22];
  assign o[11624] = i[22];
  assign o[11625] = i[22];
  assign o[11626] = i[22];
  assign o[11627] = i[22];
  assign o[11628] = i[22];
  assign o[11629] = i[22];
  assign o[11630] = i[22];
  assign o[11631] = i[22];
  assign o[11632] = i[22];
  assign o[11633] = i[22];
  assign o[11634] = i[22];
  assign o[11635] = i[22];
  assign o[11636] = i[22];
  assign o[11637] = i[22];
  assign o[11638] = i[22];
  assign o[11639] = i[22];
  assign o[11640] = i[22];
  assign o[11641] = i[22];
  assign o[11642] = i[22];
  assign o[11643] = i[22];
  assign o[11644] = i[22];
  assign o[11645] = i[22];
  assign o[11646] = i[22];
  assign o[11647] = i[22];
  assign o[11648] = i[22];
  assign o[11649] = i[22];
  assign o[11650] = i[22];
  assign o[11651] = i[22];
  assign o[11652] = i[22];
  assign o[11653] = i[22];
  assign o[11654] = i[22];
  assign o[11655] = i[22];
  assign o[11656] = i[22];
  assign o[11657] = i[22];
  assign o[11658] = i[22];
  assign o[11659] = i[22];
  assign o[11660] = i[22];
  assign o[11661] = i[22];
  assign o[11662] = i[22];
  assign o[11663] = i[22];
  assign o[11664] = i[22];
  assign o[11665] = i[22];
  assign o[11666] = i[22];
  assign o[11667] = i[22];
  assign o[11668] = i[22];
  assign o[11669] = i[22];
  assign o[11670] = i[22];
  assign o[11671] = i[22];
  assign o[11672] = i[22];
  assign o[11673] = i[22];
  assign o[11674] = i[22];
  assign o[11675] = i[22];
  assign o[11676] = i[22];
  assign o[11677] = i[22];
  assign o[11678] = i[22];
  assign o[11679] = i[22];
  assign o[11680] = i[22];
  assign o[11681] = i[22];
  assign o[11682] = i[22];
  assign o[11683] = i[22];
  assign o[11684] = i[22];
  assign o[11685] = i[22];
  assign o[11686] = i[22];
  assign o[11687] = i[22];
  assign o[11688] = i[22];
  assign o[11689] = i[22];
  assign o[11690] = i[22];
  assign o[11691] = i[22];
  assign o[11692] = i[22];
  assign o[11693] = i[22];
  assign o[11694] = i[22];
  assign o[11695] = i[22];
  assign o[11696] = i[22];
  assign o[11697] = i[22];
  assign o[11698] = i[22];
  assign o[11699] = i[22];
  assign o[11700] = i[22];
  assign o[11701] = i[22];
  assign o[11702] = i[22];
  assign o[11703] = i[22];
  assign o[11704] = i[22];
  assign o[11705] = i[22];
  assign o[11706] = i[22];
  assign o[11707] = i[22];
  assign o[11708] = i[22];
  assign o[11709] = i[22];
  assign o[11710] = i[22];
  assign o[11711] = i[22];
  assign o[11712] = i[22];
  assign o[11713] = i[22];
  assign o[11714] = i[22];
  assign o[11715] = i[22];
  assign o[11716] = i[22];
  assign o[11717] = i[22];
  assign o[11718] = i[22];
  assign o[11719] = i[22];
  assign o[11720] = i[22];
  assign o[11721] = i[22];
  assign o[11722] = i[22];
  assign o[11723] = i[22];
  assign o[11724] = i[22];
  assign o[11725] = i[22];
  assign o[11726] = i[22];
  assign o[11727] = i[22];
  assign o[11728] = i[22];
  assign o[11729] = i[22];
  assign o[11730] = i[22];
  assign o[11731] = i[22];
  assign o[11732] = i[22];
  assign o[11733] = i[22];
  assign o[11734] = i[22];
  assign o[11735] = i[22];
  assign o[11736] = i[22];
  assign o[11737] = i[22];
  assign o[11738] = i[22];
  assign o[11739] = i[22];
  assign o[11740] = i[22];
  assign o[11741] = i[22];
  assign o[11742] = i[22];
  assign o[11743] = i[22];
  assign o[11744] = i[22];
  assign o[11745] = i[22];
  assign o[11746] = i[22];
  assign o[11747] = i[22];
  assign o[11748] = i[22];
  assign o[11749] = i[22];
  assign o[11750] = i[22];
  assign o[11751] = i[22];
  assign o[11752] = i[22];
  assign o[11753] = i[22];
  assign o[11754] = i[22];
  assign o[11755] = i[22];
  assign o[11756] = i[22];
  assign o[11757] = i[22];
  assign o[11758] = i[22];
  assign o[11759] = i[22];
  assign o[11760] = i[22];
  assign o[11761] = i[22];
  assign o[11762] = i[22];
  assign o[11763] = i[22];
  assign o[11764] = i[22];
  assign o[11765] = i[22];
  assign o[11766] = i[22];
  assign o[11767] = i[22];
  assign o[11768] = i[22];
  assign o[11769] = i[22];
  assign o[11770] = i[22];
  assign o[11771] = i[22];
  assign o[11772] = i[22];
  assign o[11773] = i[22];
  assign o[11774] = i[22];
  assign o[11775] = i[22];
  assign o[10752] = i[21];
  assign o[10753] = i[21];
  assign o[10754] = i[21];
  assign o[10755] = i[21];
  assign o[10756] = i[21];
  assign o[10757] = i[21];
  assign o[10758] = i[21];
  assign o[10759] = i[21];
  assign o[10760] = i[21];
  assign o[10761] = i[21];
  assign o[10762] = i[21];
  assign o[10763] = i[21];
  assign o[10764] = i[21];
  assign o[10765] = i[21];
  assign o[10766] = i[21];
  assign o[10767] = i[21];
  assign o[10768] = i[21];
  assign o[10769] = i[21];
  assign o[10770] = i[21];
  assign o[10771] = i[21];
  assign o[10772] = i[21];
  assign o[10773] = i[21];
  assign o[10774] = i[21];
  assign o[10775] = i[21];
  assign o[10776] = i[21];
  assign o[10777] = i[21];
  assign o[10778] = i[21];
  assign o[10779] = i[21];
  assign o[10780] = i[21];
  assign o[10781] = i[21];
  assign o[10782] = i[21];
  assign o[10783] = i[21];
  assign o[10784] = i[21];
  assign o[10785] = i[21];
  assign o[10786] = i[21];
  assign o[10787] = i[21];
  assign o[10788] = i[21];
  assign o[10789] = i[21];
  assign o[10790] = i[21];
  assign o[10791] = i[21];
  assign o[10792] = i[21];
  assign o[10793] = i[21];
  assign o[10794] = i[21];
  assign o[10795] = i[21];
  assign o[10796] = i[21];
  assign o[10797] = i[21];
  assign o[10798] = i[21];
  assign o[10799] = i[21];
  assign o[10800] = i[21];
  assign o[10801] = i[21];
  assign o[10802] = i[21];
  assign o[10803] = i[21];
  assign o[10804] = i[21];
  assign o[10805] = i[21];
  assign o[10806] = i[21];
  assign o[10807] = i[21];
  assign o[10808] = i[21];
  assign o[10809] = i[21];
  assign o[10810] = i[21];
  assign o[10811] = i[21];
  assign o[10812] = i[21];
  assign o[10813] = i[21];
  assign o[10814] = i[21];
  assign o[10815] = i[21];
  assign o[10816] = i[21];
  assign o[10817] = i[21];
  assign o[10818] = i[21];
  assign o[10819] = i[21];
  assign o[10820] = i[21];
  assign o[10821] = i[21];
  assign o[10822] = i[21];
  assign o[10823] = i[21];
  assign o[10824] = i[21];
  assign o[10825] = i[21];
  assign o[10826] = i[21];
  assign o[10827] = i[21];
  assign o[10828] = i[21];
  assign o[10829] = i[21];
  assign o[10830] = i[21];
  assign o[10831] = i[21];
  assign o[10832] = i[21];
  assign o[10833] = i[21];
  assign o[10834] = i[21];
  assign o[10835] = i[21];
  assign o[10836] = i[21];
  assign o[10837] = i[21];
  assign o[10838] = i[21];
  assign o[10839] = i[21];
  assign o[10840] = i[21];
  assign o[10841] = i[21];
  assign o[10842] = i[21];
  assign o[10843] = i[21];
  assign o[10844] = i[21];
  assign o[10845] = i[21];
  assign o[10846] = i[21];
  assign o[10847] = i[21];
  assign o[10848] = i[21];
  assign o[10849] = i[21];
  assign o[10850] = i[21];
  assign o[10851] = i[21];
  assign o[10852] = i[21];
  assign o[10853] = i[21];
  assign o[10854] = i[21];
  assign o[10855] = i[21];
  assign o[10856] = i[21];
  assign o[10857] = i[21];
  assign o[10858] = i[21];
  assign o[10859] = i[21];
  assign o[10860] = i[21];
  assign o[10861] = i[21];
  assign o[10862] = i[21];
  assign o[10863] = i[21];
  assign o[10864] = i[21];
  assign o[10865] = i[21];
  assign o[10866] = i[21];
  assign o[10867] = i[21];
  assign o[10868] = i[21];
  assign o[10869] = i[21];
  assign o[10870] = i[21];
  assign o[10871] = i[21];
  assign o[10872] = i[21];
  assign o[10873] = i[21];
  assign o[10874] = i[21];
  assign o[10875] = i[21];
  assign o[10876] = i[21];
  assign o[10877] = i[21];
  assign o[10878] = i[21];
  assign o[10879] = i[21];
  assign o[10880] = i[21];
  assign o[10881] = i[21];
  assign o[10882] = i[21];
  assign o[10883] = i[21];
  assign o[10884] = i[21];
  assign o[10885] = i[21];
  assign o[10886] = i[21];
  assign o[10887] = i[21];
  assign o[10888] = i[21];
  assign o[10889] = i[21];
  assign o[10890] = i[21];
  assign o[10891] = i[21];
  assign o[10892] = i[21];
  assign o[10893] = i[21];
  assign o[10894] = i[21];
  assign o[10895] = i[21];
  assign o[10896] = i[21];
  assign o[10897] = i[21];
  assign o[10898] = i[21];
  assign o[10899] = i[21];
  assign o[10900] = i[21];
  assign o[10901] = i[21];
  assign o[10902] = i[21];
  assign o[10903] = i[21];
  assign o[10904] = i[21];
  assign o[10905] = i[21];
  assign o[10906] = i[21];
  assign o[10907] = i[21];
  assign o[10908] = i[21];
  assign o[10909] = i[21];
  assign o[10910] = i[21];
  assign o[10911] = i[21];
  assign o[10912] = i[21];
  assign o[10913] = i[21];
  assign o[10914] = i[21];
  assign o[10915] = i[21];
  assign o[10916] = i[21];
  assign o[10917] = i[21];
  assign o[10918] = i[21];
  assign o[10919] = i[21];
  assign o[10920] = i[21];
  assign o[10921] = i[21];
  assign o[10922] = i[21];
  assign o[10923] = i[21];
  assign o[10924] = i[21];
  assign o[10925] = i[21];
  assign o[10926] = i[21];
  assign o[10927] = i[21];
  assign o[10928] = i[21];
  assign o[10929] = i[21];
  assign o[10930] = i[21];
  assign o[10931] = i[21];
  assign o[10932] = i[21];
  assign o[10933] = i[21];
  assign o[10934] = i[21];
  assign o[10935] = i[21];
  assign o[10936] = i[21];
  assign o[10937] = i[21];
  assign o[10938] = i[21];
  assign o[10939] = i[21];
  assign o[10940] = i[21];
  assign o[10941] = i[21];
  assign o[10942] = i[21];
  assign o[10943] = i[21];
  assign o[10944] = i[21];
  assign o[10945] = i[21];
  assign o[10946] = i[21];
  assign o[10947] = i[21];
  assign o[10948] = i[21];
  assign o[10949] = i[21];
  assign o[10950] = i[21];
  assign o[10951] = i[21];
  assign o[10952] = i[21];
  assign o[10953] = i[21];
  assign o[10954] = i[21];
  assign o[10955] = i[21];
  assign o[10956] = i[21];
  assign o[10957] = i[21];
  assign o[10958] = i[21];
  assign o[10959] = i[21];
  assign o[10960] = i[21];
  assign o[10961] = i[21];
  assign o[10962] = i[21];
  assign o[10963] = i[21];
  assign o[10964] = i[21];
  assign o[10965] = i[21];
  assign o[10966] = i[21];
  assign o[10967] = i[21];
  assign o[10968] = i[21];
  assign o[10969] = i[21];
  assign o[10970] = i[21];
  assign o[10971] = i[21];
  assign o[10972] = i[21];
  assign o[10973] = i[21];
  assign o[10974] = i[21];
  assign o[10975] = i[21];
  assign o[10976] = i[21];
  assign o[10977] = i[21];
  assign o[10978] = i[21];
  assign o[10979] = i[21];
  assign o[10980] = i[21];
  assign o[10981] = i[21];
  assign o[10982] = i[21];
  assign o[10983] = i[21];
  assign o[10984] = i[21];
  assign o[10985] = i[21];
  assign o[10986] = i[21];
  assign o[10987] = i[21];
  assign o[10988] = i[21];
  assign o[10989] = i[21];
  assign o[10990] = i[21];
  assign o[10991] = i[21];
  assign o[10992] = i[21];
  assign o[10993] = i[21];
  assign o[10994] = i[21];
  assign o[10995] = i[21];
  assign o[10996] = i[21];
  assign o[10997] = i[21];
  assign o[10998] = i[21];
  assign o[10999] = i[21];
  assign o[11000] = i[21];
  assign o[11001] = i[21];
  assign o[11002] = i[21];
  assign o[11003] = i[21];
  assign o[11004] = i[21];
  assign o[11005] = i[21];
  assign o[11006] = i[21];
  assign o[11007] = i[21];
  assign o[11008] = i[21];
  assign o[11009] = i[21];
  assign o[11010] = i[21];
  assign o[11011] = i[21];
  assign o[11012] = i[21];
  assign o[11013] = i[21];
  assign o[11014] = i[21];
  assign o[11015] = i[21];
  assign o[11016] = i[21];
  assign o[11017] = i[21];
  assign o[11018] = i[21];
  assign o[11019] = i[21];
  assign o[11020] = i[21];
  assign o[11021] = i[21];
  assign o[11022] = i[21];
  assign o[11023] = i[21];
  assign o[11024] = i[21];
  assign o[11025] = i[21];
  assign o[11026] = i[21];
  assign o[11027] = i[21];
  assign o[11028] = i[21];
  assign o[11029] = i[21];
  assign o[11030] = i[21];
  assign o[11031] = i[21];
  assign o[11032] = i[21];
  assign o[11033] = i[21];
  assign o[11034] = i[21];
  assign o[11035] = i[21];
  assign o[11036] = i[21];
  assign o[11037] = i[21];
  assign o[11038] = i[21];
  assign o[11039] = i[21];
  assign o[11040] = i[21];
  assign o[11041] = i[21];
  assign o[11042] = i[21];
  assign o[11043] = i[21];
  assign o[11044] = i[21];
  assign o[11045] = i[21];
  assign o[11046] = i[21];
  assign o[11047] = i[21];
  assign o[11048] = i[21];
  assign o[11049] = i[21];
  assign o[11050] = i[21];
  assign o[11051] = i[21];
  assign o[11052] = i[21];
  assign o[11053] = i[21];
  assign o[11054] = i[21];
  assign o[11055] = i[21];
  assign o[11056] = i[21];
  assign o[11057] = i[21];
  assign o[11058] = i[21];
  assign o[11059] = i[21];
  assign o[11060] = i[21];
  assign o[11061] = i[21];
  assign o[11062] = i[21];
  assign o[11063] = i[21];
  assign o[11064] = i[21];
  assign o[11065] = i[21];
  assign o[11066] = i[21];
  assign o[11067] = i[21];
  assign o[11068] = i[21];
  assign o[11069] = i[21];
  assign o[11070] = i[21];
  assign o[11071] = i[21];
  assign o[11072] = i[21];
  assign o[11073] = i[21];
  assign o[11074] = i[21];
  assign o[11075] = i[21];
  assign o[11076] = i[21];
  assign o[11077] = i[21];
  assign o[11078] = i[21];
  assign o[11079] = i[21];
  assign o[11080] = i[21];
  assign o[11081] = i[21];
  assign o[11082] = i[21];
  assign o[11083] = i[21];
  assign o[11084] = i[21];
  assign o[11085] = i[21];
  assign o[11086] = i[21];
  assign o[11087] = i[21];
  assign o[11088] = i[21];
  assign o[11089] = i[21];
  assign o[11090] = i[21];
  assign o[11091] = i[21];
  assign o[11092] = i[21];
  assign o[11093] = i[21];
  assign o[11094] = i[21];
  assign o[11095] = i[21];
  assign o[11096] = i[21];
  assign o[11097] = i[21];
  assign o[11098] = i[21];
  assign o[11099] = i[21];
  assign o[11100] = i[21];
  assign o[11101] = i[21];
  assign o[11102] = i[21];
  assign o[11103] = i[21];
  assign o[11104] = i[21];
  assign o[11105] = i[21];
  assign o[11106] = i[21];
  assign o[11107] = i[21];
  assign o[11108] = i[21];
  assign o[11109] = i[21];
  assign o[11110] = i[21];
  assign o[11111] = i[21];
  assign o[11112] = i[21];
  assign o[11113] = i[21];
  assign o[11114] = i[21];
  assign o[11115] = i[21];
  assign o[11116] = i[21];
  assign o[11117] = i[21];
  assign o[11118] = i[21];
  assign o[11119] = i[21];
  assign o[11120] = i[21];
  assign o[11121] = i[21];
  assign o[11122] = i[21];
  assign o[11123] = i[21];
  assign o[11124] = i[21];
  assign o[11125] = i[21];
  assign o[11126] = i[21];
  assign o[11127] = i[21];
  assign o[11128] = i[21];
  assign o[11129] = i[21];
  assign o[11130] = i[21];
  assign o[11131] = i[21];
  assign o[11132] = i[21];
  assign o[11133] = i[21];
  assign o[11134] = i[21];
  assign o[11135] = i[21];
  assign o[11136] = i[21];
  assign o[11137] = i[21];
  assign o[11138] = i[21];
  assign o[11139] = i[21];
  assign o[11140] = i[21];
  assign o[11141] = i[21];
  assign o[11142] = i[21];
  assign o[11143] = i[21];
  assign o[11144] = i[21];
  assign o[11145] = i[21];
  assign o[11146] = i[21];
  assign o[11147] = i[21];
  assign o[11148] = i[21];
  assign o[11149] = i[21];
  assign o[11150] = i[21];
  assign o[11151] = i[21];
  assign o[11152] = i[21];
  assign o[11153] = i[21];
  assign o[11154] = i[21];
  assign o[11155] = i[21];
  assign o[11156] = i[21];
  assign o[11157] = i[21];
  assign o[11158] = i[21];
  assign o[11159] = i[21];
  assign o[11160] = i[21];
  assign o[11161] = i[21];
  assign o[11162] = i[21];
  assign o[11163] = i[21];
  assign o[11164] = i[21];
  assign o[11165] = i[21];
  assign o[11166] = i[21];
  assign o[11167] = i[21];
  assign o[11168] = i[21];
  assign o[11169] = i[21];
  assign o[11170] = i[21];
  assign o[11171] = i[21];
  assign o[11172] = i[21];
  assign o[11173] = i[21];
  assign o[11174] = i[21];
  assign o[11175] = i[21];
  assign o[11176] = i[21];
  assign o[11177] = i[21];
  assign o[11178] = i[21];
  assign o[11179] = i[21];
  assign o[11180] = i[21];
  assign o[11181] = i[21];
  assign o[11182] = i[21];
  assign o[11183] = i[21];
  assign o[11184] = i[21];
  assign o[11185] = i[21];
  assign o[11186] = i[21];
  assign o[11187] = i[21];
  assign o[11188] = i[21];
  assign o[11189] = i[21];
  assign o[11190] = i[21];
  assign o[11191] = i[21];
  assign o[11192] = i[21];
  assign o[11193] = i[21];
  assign o[11194] = i[21];
  assign o[11195] = i[21];
  assign o[11196] = i[21];
  assign o[11197] = i[21];
  assign o[11198] = i[21];
  assign o[11199] = i[21];
  assign o[11200] = i[21];
  assign o[11201] = i[21];
  assign o[11202] = i[21];
  assign o[11203] = i[21];
  assign o[11204] = i[21];
  assign o[11205] = i[21];
  assign o[11206] = i[21];
  assign o[11207] = i[21];
  assign o[11208] = i[21];
  assign o[11209] = i[21];
  assign o[11210] = i[21];
  assign o[11211] = i[21];
  assign o[11212] = i[21];
  assign o[11213] = i[21];
  assign o[11214] = i[21];
  assign o[11215] = i[21];
  assign o[11216] = i[21];
  assign o[11217] = i[21];
  assign o[11218] = i[21];
  assign o[11219] = i[21];
  assign o[11220] = i[21];
  assign o[11221] = i[21];
  assign o[11222] = i[21];
  assign o[11223] = i[21];
  assign o[11224] = i[21];
  assign o[11225] = i[21];
  assign o[11226] = i[21];
  assign o[11227] = i[21];
  assign o[11228] = i[21];
  assign o[11229] = i[21];
  assign o[11230] = i[21];
  assign o[11231] = i[21];
  assign o[11232] = i[21];
  assign o[11233] = i[21];
  assign o[11234] = i[21];
  assign o[11235] = i[21];
  assign o[11236] = i[21];
  assign o[11237] = i[21];
  assign o[11238] = i[21];
  assign o[11239] = i[21];
  assign o[11240] = i[21];
  assign o[11241] = i[21];
  assign o[11242] = i[21];
  assign o[11243] = i[21];
  assign o[11244] = i[21];
  assign o[11245] = i[21];
  assign o[11246] = i[21];
  assign o[11247] = i[21];
  assign o[11248] = i[21];
  assign o[11249] = i[21];
  assign o[11250] = i[21];
  assign o[11251] = i[21];
  assign o[11252] = i[21];
  assign o[11253] = i[21];
  assign o[11254] = i[21];
  assign o[11255] = i[21];
  assign o[11256] = i[21];
  assign o[11257] = i[21];
  assign o[11258] = i[21];
  assign o[11259] = i[21];
  assign o[11260] = i[21];
  assign o[11261] = i[21];
  assign o[11262] = i[21];
  assign o[11263] = i[21];
  assign o[10240] = i[20];
  assign o[10241] = i[20];
  assign o[10242] = i[20];
  assign o[10243] = i[20];
  assign o[10244] = i[20];
  assign o[10245] = i[20];
  assign o[10246] = i[20];
  assign o[10247] = i[20];
  assign o[10248] = i[20];
  assign o[10249] = i[20];
  assign o[10250] = i[20];
  assign o[10251] = i[20];
  assign o[10252] = i[20];
  assign o[10253] = i[20];
  assign o[10254] = i[20];
  assign o[10255] = i[20];
  assign o[10256] = i[20];
  assign o[10257] = i[20];
  assign o[10258] = i[20];
  assign o[10259] = i[20];
  assign o[10260] = i[20];
  assign o[10261] = i[20];
  assign o[10262] = i[20];
  assign o[10263] = i[20];
  assign o[10264] = i[20];
  assign o[10265] = i[20];
  assign o[10266] = i[20];
  assign o[10267] = i[20];
  assign o[10268] = i[20];
  assign o[10269] = i[20];
  assign o[10270] = i[20];
  assign o[10271] = i[20];
  assign o[10272] = i[20];
  assign o[10273] = i[20];
  assign o[10274] = i[20];
  assign o[10275] = i[20];
  assign o[10276] = i[20];
  assign o[10277] = i[20];
  assign o[10278] = i[20];
  assign o[10279] = i[20];
  assign o[10280] = i[20];
  assign o[10281] = i[20];
  assign o[10282] = i[20];
  assign o[10283] = i[20];
  assign o[10284] = i[20];
  assign o[10285] = i[20];
  assign o[10286] = i[20];
  assign o[10287] = i[20];
  assign o[10288] = i[20];
  assign o[10289] = i[20];
  assign o[10290] = i[20];
  assign o[10291] = i[20];
  assign o[10292] = i[20];
  assign o[10293] = i[20];
  assign o[10294] = i[20];
  assign o[10295] = i[20];
  assign o[10296] = i[20];
  assign o[10297] = i[20];
  assign o[10298] = i[20];
  assign o[10299] = i[20];
  assign o[10300] = i[20];
  assign o[10301] = i[20];
  assign o[10302] = i[20];
  assign o[10303] = i[20];
  assign o[10304] = i[20];
  assign o[10305] = i[20];
  assign o[10306] = i[20];
  assign o[10307] = i[20];
  assign o[10308] = i[20];
  assign o[10309] = i[20];
  assign o[10310] = i[20];
  assign o[10311] = i[20];
  assign o[10312] = i[20];
  assign o[10313] = i[20];
  assign o[10314] = i[20];
  assign o[10315] = i[20];
  assign o[10316] = i[20];
  assign o[10317] = i[20];
  assign o[10318] = i[20];
  assign o[10319] = i[20];
  assign o[10320] = i[20];
  assign o[10321] = i[20];
  assign o[10322] = i[20];
  assign o[10323] = i[20];
  assign o[10324] = i[20];
  assign o[10325] = i[20];
  assign o[10326] = i[20];
  assign o[10327] = i[20];
  assign o[10328] = i[20];
  assign o[10329] = i[20];
  assign o[10330] = i[20];
  assign o[10331] = i[20];
  assign o[10332] = i[20];
  assign o[10333] = i[20];
  assign o[10334] = i[20];
  assign o[10335] = i[20];
  assign o[10336] = i[20];
  assign o[10337] = i[20];
  assign o[10338] = i[20];
  assign o[10339] = i[20];
  assign o[10340] = i[20];
  assign o[10341] = i[20];
  assign o[10342] = i[20];
  assign o[10343] = i[20];
  assign o[10344] = i[20];
  assign o[10345] = i[20];
  assign o[10346] = i[20];
  assign o[10347] = i[20];
  assign o[10348] = i[20];
  assign o[10349] = i[20];
  assign o[10350] = i[20];
  assign o[10351] = i[20];
  assign o[10352] = i[20];
  assign o[10353] = i[20];
  assign o[10354] = i[20];
  assign o[10355] = i[20];
  assign o[10356] = i[20];
  assign o[10357] = i[20];
  assign o[10358] = i[20];
  assign o[10359] = i[20];
  assign o[10360] = i[20];
  assign o[10361] = i[20];
  assign o[10362] = i[20];
  assign o[10363] = i[20];
  assign o[10364] = i[20];
  assign o[10365] = i[20];
  assign o[10366] = i[20];
  assign o[10367] = i[20];
  assign o[10368] = i[20];
  assign o[10369] = i[20];
  assign o[10370] = i[20];
  assign o[10371] = i[20];
  assign o[10372] = i[20];
  assign o[10373] = i[20];
  assign o[10374] = i[20];
  assign o[10375] = i[20];
  assign o[10376] = i[20];
  assign o[10377] = i[20];
  assign o[10378] = i[20];
  assign o[10379] = i[20];
  assign o[10380] = i[20];
  assign o[10381] = i[20];
  assign o[10382] = i[20];
  assign o[10383] = i[20];
  assign o[10384] = i[20];
  assign o[10385] = i[20];
  assign o[10386] = i[20];
  assign o[10387] = i[20];
  assign o[10388] = i[20];
  assign o[10389] = i[20];
  assign o[10390] = i[20];
  assign o[10391] = i[20];
  assign o[10392] = i[20];
  assign o[10393] = i[20];
  assign o[10394] = i[20];
  assign o[10395] = i[20];
  assign o[10396] = i[20];
  assign o[10397] = i[20];
  assign o[10398] = i[20];
  assign o[10399] = i[20];
  assign o[10400] = i[20];
  assign o[10401] = i[20];
  assign o[10402] = i[20];
  assign o[10403] = i[20];
  assign o[10404] = i[20];
  assign o[10405] = i[20];
  assign o[10406] = i[20];
  assign o[10407] = i[20];
  assign o[10408] = i[20];
  assign o[10409] = i[20];
  assign o[10410] = i[20];
  assign o[10411] = i[20];
  assign o[10412] = i[20];
  assign o[10413] = i[20];
  assign o[10414] = i[20];
  assign o[10415] = i[20];
  assign o[10416] = i[20];
  assign o[10417] = i[20];
  assign o[10418] = i[20];
  assign o[10419] = i[20];
  assign o[10420] = i[20];
  assign o[10421] = i[20];
  assign o[10422] = i[20];
  assign o[10423] = i[20];
  assign o[10424] = i[20];
  assign o[10425] = i[20];
  assign o[10426] = i[20];
  assign o[10427] = i[20];
  assign o[10428] = i[20];
  assign o[10429] = i[20];
  assign o[10430] = i[20];
  assign o[10431] = i[20];
  assign o[10432] = i[20];
  assign o[10433] = i[20];
  assign o[10434] = i[20];
  assign o[10435] = i[20];
  assign o[10436] = i[20];
  assign o[10437] = i[20];
  assign o[10438] = i[20];
  assign o[10439] = i[20];
  assign o[10440] = i[20];
  assign o[10441] = i[20];
  assign o[10442] = i[20];
  assign o[10443] = i[20];
  assign o[10444] = i[20];
  assign o[10445] = i[20];
  assign o[10446] = i[20];
  assign o[10447] = i[20];
  assign o[10448] = i[20];
  assign o[10449] = i[20];
  assign o[10450] = i[20];
  assign o[10451] = i[20];
  assign o[10452] = i[20];
  assign o[10453] = i[20];
  assign o[10454] = i[20];
  assign o[10455] = i[20];
  assign o[10456] = i[20];
  assign o[10457] = i[20];
  assign o[10458] = i[20];
  assign o[10459] = i[20];
  assign o[10460] = i[20];
  assign o[10461] = i[20];
  assign o[10462] = i[20];
  assign o[10463] = i[20];
  assign o[10464] = i[20];
  assign o[10465] = i[20];
  assign o[10466] = i[20];
  assign o[10467] = i[20];
  assign o[10468] = i[20];
  assign o[10469] = i[20];
  assign o[10470] = i[20];
  assign o[10471] = i[20];
  assign o[10472] = i[20];
  assign o[10473] = i[20];
  assign o[10474] = i[20];
  assign o[10475] = i[20];
  assign o[10476] = i[20];
  assign o[10477] = i[20];
  assign o[10478] = i[20];
  assign o[10479] = i[20];
  assign o[10480] = i[20];
  assign o[10481] = i[20];
  assign o[10482] = i[20];
  assign o[10483] = i[20];
  assign o[10484] = i[20];
  assign o[10485] = i[20];
  assign o[10486] = i[20];
  assign o[10487] = i[20];
  assign o[10488] = i[20];
  assign o[10489] = i[20];
  assign o[10490] = i[20];
  assign o[10491] = i[20];
  assign o[10492] = i[20];
  assign o[10493] = i[20];
  assign o[10494] = i[20];
  assign o[10495] = i[20];
  assign o[10496] = i[20];
  assign o[10497] = i[20];
  assign o[10498] = i[20];
  assign o[10499] = i[20];
  assign o[10500] = i[20];
  assign o[10501] = i[20];
  assign o[10502] = i[20];
  assign o[10503] = i[20];
  assign o[10504] = i[20];
  assign o[10505] = i[20];
  assign o[10506] = i[20];
  assign o[10507] = i[20];
  assign o[10508] = i[20];
  assign o[10509] = i[20];
  assign o[10510] = i[20];
  assign o[10511] = i[20];
  assign o[10512] = i[20];
  assign o[10513] = i[20];
  assign o[10514] = i[20];
  assign o[10515] = i[20];
  assign o[10516] = i[20];
  assign o[10517] = i[20];
  assign o[10518] = i[20];
  assign o[10519] = i[20];
  assign o[10520] = i[20];
  assign o[10521] = i[20];
  assign o[10522] = i[20];
  assign o[10523] = i[20];
  assign o[10524] = i[20];
  assign o[10525] = i[20];
  assign o[10526] = i[20];
  assign o[10527] = i[20];
  assign o[10528] = i[20];
  assign o[10529] = i[20];
  assign o[10530] = i[20];
  assign o[10531] = i[20];
  assign o[10532] = i[20];
  assign o[10533] = i[20];
  assign o[10534] = i[20];
  assign o[10535] = i[20];
  assign o[10536] = i[20];
  assign o[10537] = i[20];
  assign o[10538] = i[20];
  assign o[10539] = i[20];
  assign o[10540] = i[20];
  assign o[10541] = i[20];
  assign o[10542] = i[20];
  assign o[10543] = i[20];
  assign o[10544] = i[20];
  assign o[10545] = i[20];
  assign o[10546] = i[20];
  assign o[10547] = i[20];
  assign o[10548] = i[20];
  assign o[10549] = i[20];
  assign o[10550] = i[20];
  assign o[10551] = i[20];
  assign o[10552] = i[20];
  assign o[10553] = i[20];
  assign o[10554] = i[20];
  assign o[10555] = i[20];
  assign o[10556] = i[20];
  assign o[10557] = i[20];
  assign o[10558] = i[20];
  assign o[10559] = i[20];
  assign o[10560] = i[20];
  assign o[10561] = i[20];
  assign o[10562] = i[20];
  assign o[10563] = i[20];
  assign o[10564] = i[20];
  assign o[10565] = i[20];
  assign o[10566] = i[20];
  assign o[10567] = i[20];
  assign o[10568] = i[20];
  assign o[10569] = i[20];
  assign o[10570] = i[20];
  assign o[10571] = i[20];
  assign o[10572] = i[20];
  assign o[10573] = i[20];
  assign o[10574] = i[20];
  assign o[10575] = i[20];
  assign o[10576] = i[20];
  assign o[10577] = i[20];
  assign o[10578] = i[20];
  assign o[10579] = i[20];
  assign o[10580] = i[20];
  assign o[10581] = i[20];
  assign o[10582] = i[20];
  assign o[10583] = i[20];
  assign o[10584] = i[20];
  assign o[10585] = i[20];
  assign o[10586] = i[20];
  assign o[10587] = i[20];
  assign o[10588] = i[20];
  assign o[10589] = i[20];
  assign o[10590] = i[20];
  assign o[10591] = i[20];
  assign o[10592] = i[20];
  assign o[10593] = i[20];
  assign o[10594] = i[20];
  assign o[10595] = i[20];
  assign o[10596] = i[20];
  assign o[10597] = i[20];
  assign o[10598] = i[20];
  assign o[10599] = i[20];
  assign o[10600] = i[20];
  assign o[10601] = i[20];
  assign o[10602] = i[20];
  assign o[10603] = i[20];
  assign o[10604] = i[20];
  assign o[10605] = i[20];
  assign o[10606] = i[20];
  assign o[10607] = i[20];
  assign o[10608] = i[20];
  assign o[10609] = i[20];
  assign o[10610] = i[20];
  assign o[10611] = i[20];
  assign o[10612] = i[20];
  assign o[10613] = i[20];
  assign o[10614] = i[20];
  assign o[10615] = i[20];
  assign o[10616] = i[20];
  assign o[10617] = i[20];
  assign o[10618] = i[20];
  assign o[10619] = i[20];
  assign o[10620] = i[20];
  assign o[10621] = i[20];
  assign o[10622] = i[20];
  assign o[10623] = i[20];
  assign o[10624] = i[20];
  assign o[10625] = i[20];
  assign o[10626] = i[20];
  assign o[10627] = i[20];
  assign o[10628] = i[20];
  assign o[10629] = i[20];
  assign o[10630] = i[20];
  assign o[10631] = i[20];
  assign o[10632] = i[20];
  assign o[10633] = i[20];
  assign o[10634] = i[20];
  assign o[10635] = i[20];
  assign o[10636] = i[20];
  assign o[10637] = i[20];
  assign o[10638] = i[20];
  assign o[10639] = i[20];
  assign o[10640] = i[20];
  assign o[10641] = i[20];
  assign o[10642] = i[20];
  assign o[10643] = i[20];
  assign o[10644] = i[20];
  assign o[10645] = i[20];
  assign o[10646] = i[20];
  assign o[10647] = i[20];
  assign o[10648] = i[20];
  assign o[10649] = i[20];
  assign o[10650] = i[20];
  assign o[10651] = i[20];
  assign o[10652] = i[20];
  assign o[10653] = i[20];
  assign o[10654] = i[20];
  assign o[10655] = i[20];
  assign o[10656] = i[20];
  assign o[10657] = i[20];
  assign o[10658] = i[20];
  assign o[10659] = i[20];
  assign o[10660] = i[20];
  assign o[10661] = i[20];
  assign o[10662] = i[20];
  assign o[10663] = i[20];
  assign o[10664] = i[20];
  assign o[10665] = i[20];
  assign o[10666] = i[20];
  assign o[10667] = i[20];
  assign o[10668] = i[20];
  assign o[10669] = i[20];
  assign o[10670] = i[20];
  assign o[10671] = i[20];
  assign o[10672] = i[20];
  assign o[10673] = i[20];
  assign o[10674] = i[20];
  assign o[10675] = i[20];
  assign o[10676] = i[20];
  assign o[10677] = i[20];
  assign o[10678] = i[20];
  assign o[10679] = i[20];
  assign o[10680] = i[20];
  assign o[10681] = i[20];
  assign o[10682] = i[20];
  assign o[10683] = i[20];
  assign o[10684] = i[20];
  assign o[10685] = i[20];
  assign o[10686] = i[20];
  assign o[10687] = i[20];
  assign o[10688] = i[20];
  assign o[10689] = i[20];
  assign o[10690] = i[20];
  assign o[10691] = i[20];
  assign o[10692] = i[20];
  assign o[10693] = i[20];
  assign o[10694] = i[20];
  assign o[10695] = i[20];
  assign o[10696] = i[20];
  assign o[10697] = i[20];
  assign o[10698] = i[20];
  assign o[10699] = i[20];
  assign o[10700] = i[20];
  assign o[10701] = i[20];
  assign o[10702] = i[20];
  assign o[10703] = i[20];
  assign o[10704] = i[20];
  assign o[10705] = i[20];
  assign o[10706] = i[20];
  assign o[10707] = i[20];
  assign o[10708] = i[20];
  assign o[10709] = i[20];
  assign o[10710] = i[20];
  assign o[10711] = i[20];
  assign o[10712] = i[20];
  assign o[10713] = i[20];
  assign o[10714] = i[20];
  assign o[10715] = i[20];
  assign o[10716] = i[20];
  assign o[10717] = i[20];
  assign o[10718] = i[20];
  assign o[10719] = i[20];
  assign o[10720] = i[20];
  assign o[10721] = i[20];
  assign o[10722] = i[20];
  assign o[10723] = i[20];
  assign o[10724] = i[20];
  assign o[10725] = i[20];
  assign o[10726] = i[20];
  assign o[10727] = i[20];
  assign o[10728] = i[20];
  assign o[10729] = i[20];
  assign o[10730] = i[20];
  assign o[10731] = i[20];
  assign o[10732] = i[20];
  assign o[10733] = i[20];
  assign o[10734] = i[20];
  assign o[10735] = i[20];
  assign o[10736] = i[20];
  assign o[10737] = i[20];
  assign o[10738] = i[20];
  assign o[10739] = i[20];
  assign o[10740] = i[20];
  assign o[10741] = i[20];
  assign o[10742] = i[20];
  assign o[10743] = i[20];
  assign o[10744] = i[20];
  assign o[10745] = i[20];
  assign o[10746] = i[20];
  assign o[10747] = i[20];
  assign o[10748] = i[20];
  assign o[10749] = i[20];
  assign o[10750] = i[20];
  assign o[10751] = i[20];
  assign o[9728] = i[19];
  assign o[9729] = i[19];
  assign o[9730] = i[19];
  assign o[9731] = i[19];
  assign o[9732] = i[19];
  assign o[9733] = i[19];
  assign o[9734] = i[19];
  assign o[9735] = i[19];
  assign o[9736] = i[19];
  assign o[9737] = i[19];
  assign o[9738] = i[19];
  assign o[9739] = i[19];
  assign o[9740] = i[19];
  assign o[9741] = i[19];
  assign o[9742] = i[19];
  assign o[9743] = i[19];
  assign o[9744] = i[19];
  assign o[9745] = i[19];
  assign o[9746] = i[19];
  assign o[9747] = i[19];
  assign o[9748] = i[19];
  assign o[9749] = i[19];
  assign o[9750] = i[19];
  assign o[9751] = i[19];
  assign o[9752] = i[19];
  assign o[9753] = i[19];
  assign o[9754] = i[19];
  assign o[9755] = i[19];
  assign o[9756] = i[19];
  assign o[9757] = i[19];
  assign o[9758] = i[19];
  assign o[9759] = i[19];
  assign o[9760] = i[19];
  assign o[9761] = i[19];
  assign o[9762] = i[19];
  assign o[9763] = i[19];
  assign o[9764] = i[19];
  assign o[9765] = i[19];
  assign o[9766] = i[19];
  assign o[9767] = i[19];
  assign o[9768] = i[19];
  assign o[9769] = i[19];
  assign o[9770] = i[19];
  assign o[9771] = i[19];
  assign o[9772] = i[19];
  assign o[9773] = i[19];
  assign o[9774] = i[19];
  assign o[9775] = i[19];
  assign o[9776] = i[19];
  assign o[9777] = i[19];
  assign o[9778] = i[19];
  assign o[9779] = i[19];
  assign o[9780] = i[19];
  assign o[9781] = i[19];
  assign o[9782] = i[19];
  assign o[9783] = i[19];
  assign o[9784] = i[19];
  assign o[9785] = i[19];
  assign o[9786] = i[19];
  assign o[9787] = i[19];
  assign o[9788] = i[19];
  assign o[9789] = i[19];
  assign o[9790] = i[19];
  assign o[9791] = i[19];
  assign o[9792] = i[19];
  assign o[9793] = i[19];
  assign o[9794] = i[19];
  assign o[9795] = i[19];
  assign o[9796] = i[19];
  assign o[9797] = i[19];
  assign o[9798] = i[19];
  assign o[9799] = i[19];
  assign o[9800] = i[19];
  assign o[9801] = i[19];
  assign o[9802] = i[19];
  assign o[9803] = i[19];
  assign o[9804] = i[19];
  assign o[9805] = i[19];
  assign o[9806] = i[19];
  assign o[9807] = i[19];
  assign o[9808] = i[19];
  assign o[9809] = i[19];
  assign o[9810] = i[19];
  assign o[9811] = i[19];
  assign o[9812] = i[19];
  assign o[9813] = i[19];
  assign o[9814] = i[19];
  assign o[9815] = i[19];
  assign o[9816] = i[19];
  assign o[9817] = i[19];
  assign o[9818] = i[19];
  assign o[9819] = i[19];
  assign o[9820] = i[19];
  assign o[9821] = i[19];
  assign o[9822] = i[19];
  assign o[9823] = i[19];
  assign o[9824] = i[19];
  assign o[9825] = i[19];
  assign o[9826] = i[19];
  assign o[9827] = i[19];
  assign o[9828] = i[19];
  assign o[9829] = i[19];
  assign o[9830] = i[19];
  assign o[9831] = i[19];
  assign o[9832] = i[19];
  assign o[9833] = i[19];
  assign o[9834] = i[19];
  assign o[9835] = i[19];
  assign o[9836] = i[19];
  assign o[9837] = i[19];
  assign o[9838] = i[19];
  assign o[9839] = i[19];
  assign o[9840] = i[19];
  assign o[9841] = i[19];
  assign o[9842] = i[19];
  assign o[9843] = i[19];
  assign o[9844] = i[19];
  assign o[9845] = i[19];
  assign o[9846] = i[19];
  assign o[9847] = i[19];
  assign o[9848] = i[19];
  assign o[9849] = i[19];
  assign o[9850] = i[19];
  assign o[9851] = i[19];
  assign o[9852] = i[19];
  assign o[9853] = i[19];
  assign o[9854] = i[19];
  assign o[9855] = i[19];
  assign o[9856] = i[19];
  assign o[9857] = i[19];
  assign o[9858] = i[19];
  assign o[9859] = i[19];
  assign o[9860] = i[19];
  assign o[9861] = i[19];
  assign o[9862] = i[19];
  assign o[9863] = i[19];
  assign o[9864] = i[19];
  assign o[9865] = i[19];
  assign o[9866] = i[19];
  assign o[9867] = i[19];
  assign o[9868] = i[19];
  assign o[9869] = i[19];
  assign o[9870] = i[19];
  assign o[9871] = i[19];
  assign o[9872] = i[19];
  assign o[9873] = i[19];
  assign o[9874] = i[19];
  assign o[9875] = i[19];
  assign o[9876] = i[19];
  assign o[9877] = i[19];
  assign o[9878] = i[19];
  assign o[9879] = i[19];
  assign o[9880] = i[19];
  assign o[9881] = i[19];
  assign o[9882] = i[19];
  assign o[9883] = i[19];
  assign o[9884] = i[19];
  assign o[9885] = i[19];
  assign o[9886] = i[19];
  assign o[9887] = i[19];
  assign o[9888] = i[19];
  assign o[9889] = i[19];
  assign o[9890] = i[19];
  assign o[9891] = i[19];
  assign o[9892] = i[19];
  assign o[9893] = i[19];
  assign o[9894] = i[19];
  assign o[9895] = i[19];
  assign o[9896] = i[19];
  assign o[9897] = i[19];
  assign o[9898] = i[19];
  assign o[9899] = i[19];
  assign o[9900] = i[19];
  assign o[9901] = i[19];
  assign o[9902] = i[19];
  assign o[9903] = i[19];
  assign o[9904] = i[19];
  assign o[9905] = i[19];
  assign o[9906] = i[19];
  assign o[9907] = i[19];
  assign o[9908] = i[19];
  assign o[9909] = i[19];
  assign o[9910] = i[19];
  assign o[9911] = i[19];
  assign o[9912] = i[19];
  assign o[9913] = i[19];
  assign o[9914] = i[19];
  assign o[9915] = i[19];
  assign o[9916] = i[19];
  assign o[9917] = i[19];
  assign o[9918] = i[19];
  assign o[9919] = i[19];
  assign o[9920] = i[19];
  assign o[9921] = i[19];
  assign o[9922] = i[19];
  assign o[9923] = i[19];
  assign o[9924] = i[19];
  assign o[9925] = i[19];
  assign o[9926] = i[19];
  assign o[9927] = i[19];
  assign o[9928] = i[19];
  assign o[9929] = i[19];
  assign o[9930] = i[19];
  assign o[9931] = i[19];
  assign o[9932] = i[19];
  assign o[9933] = i[19];
  assign o[9934] = i[19];
  assign o[9935] = i[19];
  assign o[9936] = i[19];
  assign o[9937] = i[19];
  assign o[9938] = i[19];
  assign o[9939] = i[19];
  assign o[9940] = i[19];
  assign o[9941] = i[19];
  assign o[9942] = i[19];
  assign o[9943] = i[19];
  assign o[9944] = i[19];
  assign o[9945] = i[19];
  assign o[9946] = i[19];
  assign o[9947] = i[19];
  assign o[9948] = i[19];
  assign o[9949] = i[19];
  assign o[9950] = i[19];
  assign o[9951] = i[19];
  assign o[9952] = i[19];
  assign o[9953] = i[19];
  assign o[9954] = i[19];
  assign o[9955] = i[19];
  assign o[9956] = i[19];
  assign o[9957] = i[19];
  assign o[9958] = i[19];
  assign o[9959] = i[19];
  assign o[9960] = i[19];
  assign o[9961] = i[19];
  assign o[9962] = i[19];
  assign o[9963] = i[19];
  assign o[9964] = i[19];
  assign o[9965] = i[19];
  assign o[9966] = i[19];
  assign o[9967] = i[19];
  assign o[9968] = i[19];
  assign o[9969] = i[19];
  assign o[9970] = i[19];
  assign o[9971] = i[19];
  assign o[9972] = i[19];
  assign o[9973] = i[19];
  assign o[9974] = i[19];
  assign o[9975] = i[19];
  assign o[9976] = i[19];
  assign o[9977] = i[19];
  assign o[9978] = i[19];
  assign o[9979] = i[19];
  assign o[9980] = i[19];
  assign o[9981] = i[19];
  assign o[9982] = i[19];
  assign o[9983] = i[19];
  assign o[9984] = i[19];
  assign o[9985] = i[19];
  assign o[9986] = i[19];
  assign o[9987] = i[19];
  assign o[9988] = i[19];
  assign o[9989] = i[19];
  assign o[9990] = i[19];
  assign o[9991] = i[19];
  assign o[9992] = i[19];
  assign o[9993] = i[19];
  assign o[9994] = i[19];
  assign o[9995] = i[19];
  assign o[9996] = i[19];
  assign o[9997] = i[19];
  assign o[9998] = i[19];
  assign o[9999] = i[19];
  assign o[10000] = i[19];
  assign o[10001] = i[19];
  assign o[10002] = i[19];
  assign o[10003] = i[19];
  assign o[10004] = i[19];
  assign o[10005] = i[19];
  assign o[10006] = i[19];
  assign o[10007] = i[19];
  assign o[10008] = i[19];
  assign o[10009] = i[19];
  assign o[10010] = i[19];
  assign o[10011] = i[19];
  assign o[10012] = i[19];
  assign o[10013] = i[19];
  assign o[10014] = i[19];
  assign o[10015] = i[19];
  assign o[10016] = i[19];
  assign o[10017] = i[19];
  assign o[10018] = i[19];
  assign o[10019] = i[19];
  assign o[10020] = i[19];
  assign o[10021] = i[19];
  assign o[10022] = i[19];
  assign o[10023] = i[19];
  assign o[10024] = i[19];
  assign o[10025] = i[19];
  assign o[10026] = i[19];
  assign o[10027] = i[19];
  assign o[10028] = i[19];
  assign o[10029] = i[19];
  assign o[10030] = i[19];
  assign o[10031] = i[19];
  assign o[10032] = i[19];
  assign o[10033] = i[19];
  assign o[10034] = i[19];
  assign o[10035] = i[19];
  assign o[10036] = i[19];
  assign o[10037] = i[19];
  assign o[10038] = i[19];
  assign o[10039] = i[19];
  assign o[10040] = i[19];
  assign o[10041] = i[19];
  assign o[10042] = i[19];
  assign o[10043] = i[19];
  assign o[10044] = i[19];
  assign o[10045] = i[19];
  assign o[10046] = i[19];
  assign o[10047] = i[19];
  assign o[10048] = i[19];
  assign o[10049] = i[19];
  assign o[10050] = i[19];
  assign o[10051] = i[19];
  assign o[10052] = i[19];
  assign o[10053] = i[19];
  assign o[10054] = i[19];
  assign o[10055] = i[19];
  assign o[10056] = i[19];
  assign o[10057] = i[19];
  assign o[10058] = i[19];
  assign o[10059] = i[19];
  assign o[10060] = i[19];
  assign o[10061] = i[19];
  assign o[10062] = i[19];
  assign o[10063] = i[19];
  assign o[10064] = i[19];
  assign o[10065] = i[19];
  assign o[10066] = i[19];
  assign o[10067] = i[19];
  assign o[10068] = i[19];
  assign o[10069] = i[19];
  assign o[10070] = i[19];
  assign o[10071] = i[19];
  assign o[10072] = i[19];
  assign o[10073] = i[19];
  assign o[10074] = i[19];
  assign o[10075] = i[19];
  assign o[10076] = i[19];
  assign o[10077] = i[19];
  assign o[10078] = i[19];
  assign o[10079] = i[19];
  assign o[10080] = i[19];
  assign o[10081] = i[19];
  assign o[10082] = i[19];
  assign o[10083] = i[19];
  assign o[10084] = i[19];
  assign o[10085] = i[19];
  assign o[10086] = i[19];
  assign o[10087] = i[19];
  assign o[10088] = i[19];
  assign o[10089] = i[19];
  assign o[10090] = i[19];
  assign o[10091] = i[19];
  assign o[10092] = i[19];
  assign o[10093] = i[19];
  assign o[10094] = i[19];
  assign o[10095] = i[19];
  assign o[10096] = i[19];
  assign o[10097] = i[19];
  assign o[10098] = i[19];
  assign o[10099] = i[19];
  assign o[10100] = i[19];
  assign o[10101] = i[19];
  assign o[10102] = i[19];
  assign o[10103] = i[19];
  assign o[10104] = i[19];
  assign o[10105] = i[19];
  assign o[10106] = i[19];
  assign o[10107] = i[19];
  assign o[10108] = i[19];
  assign o[10109] = i[19];
  assign o[10110] = i[19];
  assign o[10111] = i[19];
  assign o[10112] = i[19];
  assign o[10113] = i[19];
  assign o[10114] = i[19];
  assign o[10115] = i[19];
  assign o[10116] = i[19];
  assign o[10117] = i[19];
  assign o[10118] = i[19];
  assign o[10119] = i[19];
  assign o[10120] = i[19];
  assign o[10121] = i[19];
  assign o[10122] = i[19];
  assign o[10123] = i[19];
  assign o[10124] = i[19];
  assign o[10125] = i[19];
  assign o[10126] = i[19];
  assign o[10127] = i[19];
  assign o[10128] = i[19];
  assign o[10129] = i[19];
  assign o[10130] = i[19];
  assign o[10131] = i[19];
  assign o[10132] = i[19];
  assign o[10133] = i[19];
  assign o[10134] = i[19];
  assign o[10135] = i[19];
  assign o[10136] = i[19];
  assign o[10137] = i[19];
  assign o[10138] = i[19];
  assign o[10139] = i[19];
  assign o[10140] = i[19];
  assign o[10141] = i[19];
  assign o[10142] = i[19];
  assign o[10143] = i[19];
  assign o[10144] = i[19];
  assign o[10145] = i[19];
  assign o[10146] = i[19];
  assign o[10147] = i[19];
  assign o[10148] = i[19];
  assign o[10149] = i[19];
  assign o[10150] = i[19];
  assign o[10151] = i[19];
  assign o[10152] = i[19];
  assign o[10153] = i[19];
  assign o[10154] = i[19];
  assign o[10155] = i[19];
  assign o[10156] = i[19];
  assign o[10157] = i[19];
  assign o[10158] = i[19];
  assign o[10159] = i[19];
  assign o[10160] = i[19];
  assign o[10161] = i[19];
  assign o[10162] = i[19];
  assign o[10163] = i[19];
  assign o[10164] = i[19];
  assign o[10165] = i[19];
  assign o[10166] = i[19];
  assign o[10167] = i[19];
  assign o[10168] = i[19];
  assign o[10169] = i[19];
  assign o[10170] = i[19];
  assign o[10171] = i[19];
  assign o[10172] = i[19];
  assign o[10173] = i[19];
  assign o[10174] = i[19];
  assign o[10175] = i[19];
  assign o[10176] = i[19];
  assign o[10177] = i[19];
  assign o[10178] = i[19];
  assign o[10179] = i[19];
  assign o[10180] = i[19];
  assign o[10181] = i[19];
  assign o[10182] = i[19];
  assign o[10183] = i[19];
  assign o[10184] = i[19];
  assign o[10185] = i[19];
  assign o[10186] = i[19];
  assign o[10187] = i[19];
  assign o[10188] = i[19];
  assign o[10189] = i[19];
  assign o[10190] = i[19];
  assign o[10191] = i[19];
  assign o[10192] = i[19];
  assign o[10193] = i[19];
  assign o[10194] = i[19];
  assign o[10195] = i[19];
  assign o[10196] = i[19];
  assign o[10197] = i[19];
  assign o[10198] = i[19];
  assign o[10199] = i[19];
  assign o[10200] = i[19];
  assign o[10201] = i[19];
  assign o[10202] = i[19];
  assign o[10203] = i[19];
  assign o[10204] = i[19];
  assign o[10205] = i[19];
  assign o[10206] = i[19];
  assign o[10207] = i[19];
  assign o[10208] = i[19];
  assign o[10209] = i[19];
  assign o[10210] = i[19];
  assign o[10211] = i[19];
  assign o[10212] = i[19];
  assign o[10213] = i[19];
  assign o[10214] = i[19];
  assign o[10215] = i[19];
  assign o[10216] = i[19];
  assign o[10217] = i[19];
  assign o[10218] = i[19];
  assign o[10219] = i[19];
  assign o[10220] = i[19];
  assign o[10221] = i[19];
  assign o[10222] = i[19];
  assign o[10223] = i[19];
  assign o[10224] = i[19];
  assign o[10225] = i[19];
  assign o[10226] = i[19];
  assign o[10227] = i[19];
  assign o[10228] = i[19];
  assign o[10229] = i[19];
  assign o[10230] = i[19];
  assign o[10231] = i[19];
  assign o[10232] = i[19];
  assign o[10233] = i[19];
  assign o[10234] = i[19];
  assign o[10235] = i[19];
  assign o[10236] = i[19];
  assign o[10237] = i[19];
  assign o[10238] = i[19];
  assign o[10239] = i[19];
  assign o[9216] = i[18];
  assign o[9217] = i[18];
  assign o[9218] = i[18];
  assign o[9219] = i[18];
  assign o[9220] = i[18];
  assign o[9221] = i[18];
  assign o[9222] = i[18];
  assign o[9223] = i[18];
  assign o[9224] = i[18];
  assign o[9225] = i[18];
  assign o[9226] = i[18];
  assign o[9227] = i[18];
  assign o[9228] = i[18];
  assign o[9229] = i[18];
  assign o[9230] = i[18];
  assign o[9231] = i[18];
  assign o[9232] = i[18];
  assign o[9233] = i[18];
  assign o[9234] = i[18];
  assign o[9235] = i[18];
  assign o[9236] = i[18];
  assign o[9237] = i[18];
  assign o[9238] = i[18];
  assign o[9239] = i[18];
  assign o[9240] = i[18];
  assign o[9241] = i[18];
  assign o[9242] = i[18];
  assign o[9243] = i[18];
  assign o[9244] = i[18];
  assign o[9245] = i[18];
  assign o[9246] = i[18];
  assign o[9247] = i[18];
  assign o[9248] = i[18];
  assign o[9249] = i[18];
  assign o[9250] = i[18];
  assign o[9251] = i[18];
  assign o[9252] = i[18];
  assign o[9253] = i[18];
  assign o[9254] = i[18];
  assign o[9255] = i[18];
  assign o[9256] = i[18];
  assign o[9257] = i[18];
  assign o[9258] = i[18];
  assign o[9259] = i[18];
  assign o[9260] = i[18];
  assign o[9261] = i[18];
  assign o[9262] = i[18];
  assign o[9263] = i[18];
  assign o[9264] = i[18];
  assign o[9265] = i[18];
  assign o[9266] = i[18];
  assign o[9267] = i[18];
  assign o[9268] = i[18];
  assign o[9269] = i[18];
  assign o[9270] = i[18];
  assign o[9271] = i[18];
  assign o[9272] = i[18];
  assign o[9273] = i[18];
  assign o[9274] = i[18];
  assign o[9275] = i[18];
  assign o[9276] = i[18];
  assign o[9277] = i[18];
  assign o[9278] = i[18];
  assign o[9279] = i[18];
  assign o[9280] = i[18];
  assign o[9281] = i[18];
  assign o[9282] = i[18];
  assign o[9283] = i[18];
  assign o[9284] = i[18];
  assign o[9285] = i[18];
  assign o[9286] = i[18];
  assign o[9287] = i[18];
  assign o[9288] = i[18];
  assign o[9289] = i[18];
  assign o[9290] = i[18];
  assign o[9291] = i[18];
  assign o[9292] = i[18];
  assign o[9293] = i[18];
  assign o[9294] = i[18];
  assign o[9295] = i[18];
  assign o[9296] = i[18];
  assign o[9297] = i[18];
  assign o[9298] = i[18];
  assign o[9299] = i[18];
  assign o[9300] = i[18];
  assign o[9301] = i[18];
  assign o[9302] = i[18];
  assign o[9303] = i[18];
  assign o[9304] = i[18];
  assign o[9305] = i[18];
  assign o[9306] = i[18];
  assign o[9307] = i[18];
  assign o[9308] = i[18];
  assign o[9309] = i[18];
  assign o[9310] = i[18];
  assign o[9311] = i[18];
  assign o[9312] = i[18];
  assign o[9313] = i[18];
  assign o[9314] = i[18];
  assign o[9315] = i[18];
  assign o[9316] = i[18];
  assign o[9317] = i[18];
  assign o[9318] = i[18];
  assign o[9319] = i[18];
  assign o[9320] = i[18];
  assign o[9321] = i[18];
  assign o[9322] = i[18];
  assign o[9323] = i[18];
  assign o[9324] = i[18];
  assign o[9325] = i[18];
  assign o[9326] = i[18];
  assign o[9327] = i[18];
  assign o[9328] = i[18];
  assign o[9329] = i[18];
  assign o[9330] = i[18];
  assign o[9331] = i[18];
  assign o[9332] = i[18];
  assign o[9333] = i[18];
  assign o[9334] = i[18];
  assign o[9335] = i[18];
  assign o[9336] = i[18];
  assign o[9337] = i[18];
  assign o[9338] = i[18];
  assign o[9339] = i[18];
  assign o[9340] = i[18];
  assign o[9341] = i[18];
  assign o[9342] = i[18];
  assign o[9343] = i[18];
  assign o[9344] = i[18];
  assign o[9345] = i[18];
  assign o[9346] = i[18];
  assign o[9347] = i[18];
  assign o[9348] = i[18];
  assign o[9349] = i[18];
  assign o[9350] = i[18];
  assign o[9351] = i[18];
  assign o[9352] = i[18];
  assign o[9353] = i[18];
  assign o[9354] = i[18];
  assign o[9355] = i[18];
  assign o[9356] = i[18];
  assign o[9357] = i[18];
  assign o[9358] = i[18];
  assign o[9359] = i[18];
  assign o[9360] = i[18];
  assign o[9361] = i[18];
  assign o[9362] = i[18];
  assign o[9363] = i[18];
  assign o[9364] = i[18];
  assign o[9365] = i[18];
  assign o[9366] = i[18];
  assign o[9367] = i[18];
  assign o[9368] = i[18];
  assign o[9369] = i[18];
  assign o[9370] = i[18];
  assign o[9371] = i[18];
  assign o[9372] = i[18];
  assign o[9373] = i[18];
  assign o[9374] = i[18];
  assign o[9375] = i[18];
  assign o[9376] = i[18];
  assign o[9377] = i[18];
  assign o[9378] = i[18];
  assign o[9379] = i[18];
  assign o[9380] = i[18];
  assign o[9381] = i[18];
  assign o[9382] = i[18];
  assign o[9383] = i[18];
  assign o[9384] = i[18];
  assign o[9385] = i[18];
  assign o[9386] = i[18];
  assign o[9387] = i[18];
  assign o[9388] = i[18];
  assign o[9389] = i[18];
  assign o[9390] = i[18];
  assign o[9391] = i[18];
  assign o[9392] = i[18];
  assign o[9393] = i[18];
  assign o[9394] = i[18];
  assign o[9395] = i[18];
  assign o[9396] = i[18];
  assign o[9397] = i[18];
  assign o[9398] = i[18];
  assign o[9399] = i[18];
  assign o[9400] = i[18];
  assign o[9401] = i[18];
  assign o[9402] = i[18];
  assign o[9403] = i[18];
  assign o[9404] = i[18];
  assign o[9405] = i[18];
  assign o[9406] = i[18];
  assign o[9407] = i[18];
  assign o[9408] = i[18];
  assign o[9409] = i[18];
  assign o[9410] = i[18];
  assign o[9411] = i[18];
  assign o[9412] = i[18];
  assign o[9413] = i[18];
  assign o[9414] = i[18];
  assign o[9415] = i[18];
  assign o[9416] = i[18];
  assign o[9417] = i[18];
  assign o[9418] = i[18];
  assign o[9419] = i[18];
  assign o[9420] = i[18];
  assign o[9421] = i[18];
  assign o[9422] = i[18];
  assign o[9423] = i[18];
  assign o[9424] = i[18];
  assign o[9425] = i[18];
  assign o[9426] = i[18];
  assign o[9427] = i[18];
  assign o[9428] = i[18];
  assign o[9429] = i[18];
  assign o[9430] = i[18];
  assign o[9431] = i[18];
  assign o[9432] = i[18];
  assign o[9433] = i[18];
  assign o[9434] = i[18];
  assign o[9435] = i[18];
  assign o[9436] = i[18];
  assign o[9437] = i[18];
  assign o[9438] = i[18];
  assign o[9439] = i[18];
  assign o[9440] = i[18];
  assign o[9441] = i[18];
  assign o[9442] = i[18];
  assign o[9443] = i[18];
  assign o[9444] = i[18];
  assign o[9445] = i[18];
  assign o[9446] = i[18];
  assign o[9447] = i[18];
  assign o[9448] = i[18];
  assign o[9449] = i[18];
  assign o[9450] = i[18];
  assign o[9451] = i[18];
  assign o[9452] = i[18];
  assign o[9453] = i[18];
  assign o[9454] = i[18];
  assign o[9455] = i[18];
  assign o[9456] = i[18];
  assign o[9457] = i[18];
  assign o[9458] = i[18];
  assign o[9459] = i[18];
  assign o[9460] = i[18];
  assign o[9461] = i[18];
  assign o[9462] = i[18];
  assign o[9463] = i[18];
  assign o[9464] = i[18];
  assign o[9465] = i[18];
  assign o[9466] = i[18];
  assign o[9467] = i[18];
  assign o[9468] = i[18];
  assign o[9469] = i[18];
  assign o[9470] = i[18];
  assign o[9471] = i[18];
  assign o[9472] = i[18];
  assign o[9473] = i[18];
  assign o[9474] = i[18];
  assign o[9475] = i[18];
  assign o[9476] = i[18];
  assign o[9477] = i[18];
  assign o[9478] = i[18];
  assign o[9479] = i[18];
  assign o[9480] = i[18];
  assign o[9481] = i[18];
  assign o[9482] = i[18];
  assign o[9483] = i[18];
  assign o[9484] = i[18];
  assign o[9485] = i[18];
  assign o[9486] = i[18];
  assign o[9487] = i[18];
  assign o[9488] = i[18];
  assign o[9489] = i[18];
  assign o[9490] = i[18];
  assign o[9491] = i[18];
  assign o[9492] = i[18];
  assign o[9493] = i[18];
  assign o[9494] = i[18];
  assign o[9495] = i[18];
  assign o[9496] = i[18];
  assign o[9497] = i[18];
  assign o[9498] = i[18];
  assign o[9499] = i[18];
  assign o[9500] = i[18];
  assign o[9501] = i[18];
  assign o[9502] = i[18];
  assign o[9503] = i[18];
  assign o[9504] = i[18];
  assign o[9505] = i[18];
  assign o[9506] = i[18];
  assign o[9507] = i[18];
  assign o[9508] = i[18];
  assign o[9509] = i[18];
  assign o[9510] = i[18];
  assign o[9511] = i[18];
  assign o[9512] = i[18];
  assign o[9513] = i[18];
  assign o[9514] = i[18];
  assign o[9515] = i[18];
  assign o[9516] = i[18];
  assign o[9517] = i[18];
  assign o[9518] = i[18];
  assign o[9519] = i[18];
  assign o[9520] = i[18];
  assign o[9521] = i[18];
  assign o[9522] = i[18];
  assign o[9523] = i[18];
  assign o[9524] = i[18];
  assign o[9525] = i[18];
  assign o[9526] = i[18];
  assign o[9527] = i[18];
  assign o[9528] = i[18];
  assign o[9529] = i[18];
  assign o[9530] = i[18];
  assign o[9531] = i[18];
  assign o[9532] = i[18];
  assign o[9533] = i[18];
  assign o[9534] = i[18];
  assign o[9535] = i[18];
  assign o[9536] = i[18];
  assign o[9537] = i[18];
  assign o[9538] = i[18];
  assign o[9539] = i[18];
  assign o[9540] = i[18];
  assign o[9541] = i[18];
  assign o[9542] = i[18];
  assign o[9543] = i[18];
  assign o[9544] = i[18];
  assign o[9545] = i[18];
  assign o[9546] = i[18];
  assign o[9547] = i[18];
  assign o[9548] = i[18];
  assign o[9549] = i[18];
  assign o[9550] = i[18];
  assign o[9551] = i[18];
  assign o[9552] = i[18];
  assign o[9553] = i[18];
  assign o[9554] = i[18];
  assign o[9555] = i[18];
  assign o[9556] = i[18];
  assign o[9557] = i[18];
  assign o[9558] = i[18];
  assign o[9559] = i[18];
  assign o[9560] = i[18];
  assign o[9561] = i[18];
  assign o[9562] = i[18];
  assign o[9563] = i[18];
  assign o[9564] = i[18];
  assign o[9565] = i[18];
  assign o[9566] = i[18];
  assign o[9567] = i[18];
  assign o[9568] = i[18];
  assign o[9569] = i[18];
  assign o[9570] = i[18];
  assign o[9571] = i[18];
  assign o[9572] = i[18];
  assign o[9573] = i[18];
  assign o[9574] = i[18];
  assign o[9575] = i[18];
  assign o[9576] = i[18];
  assign o[9577] = i[18];
  assign o[9578] = i[18];
  assign o[9579] = i[18];
  assign o[9580] = i[18];
  assign o[9581] = i[18];
  assign o[9582] = i[18];
  assign o[9583] = i[18];
  assign o[9584] = i[18];
  assign o[9585] = i[18];
  assign o[9586] = i[18];
  assign o[9587] = i[18];
  assign o[9588] = i[18];
  assign o[9589] = i[18];
  assign o[9590] = i[18];
  assign o[9591] = i[18];
  assign o[9592] = i[18];
  assign o[9593] = i[18];
  assign o[9594] = i[18];
  assign o[9595] = i[18];
  assign o[9596] = i[18];
  assign o[9597] = i[18];
  assign o[9598] = i[18];
  assign o[9599] = i[18];
  assign o[9600] = i[18];
  assign o[9601] = i[18];
  assign o[9602] = i[18];
  assign o[9603] = i[18];
  assign o[9604] = i[18];
  assign o[9605] = i[18];
  assign o[9606] = i[18];
  assign o[9607] = i[18];
  assign o[9608] = i[18];
  assign o[9609] = i[18];
  assign o[9610] = i[18];
  assign o[9611] = i[18];
  assign o[9612] = i[18];
  assign o[9613] = i[18];
  assign o[9614] = i[18];
  assign o[9615] = i[18];
  assign o[9616] = i[18];
  assign o[9617] = i[18];
  assign o[9618] = i[18];
  assign o[9619] = i[18];
  assign o[9620] = i[18];
  assign o[9621] = i[18];
  assign o[9622] = i[18];
  assign o[9623] = i[18];
  assign o[9624] = i[18];
  assign o[9625] = i[18];
  assign o[9626] = i[18];
  assign o[9627] = i[18];
  assign o[9628] = i[18];
  assign o[9629] = i[18];
  assign o[9630] = i[18];
  assign o[9631] = i[18];
  assign o[9632] = i[18];
  assign o[9633] = i[18];
  assign o[9634] = i[18];
  assign o[9635] = i[18];
  assign o[9636] = i[18];
  assign o[9637] = i[18];
  assign o[9638] = i[18];
  assign o[9639] = i[18];
  assign o[9640] = i[18];
  assign o[9641] = i[18];
  assign o[9642] = i[18];
  assign o[9643] = i[18];
  assign o[9644] = i[18];
  assign o[9645] = i[18];
  assign o[9646] = i[18];
  assign o[9647] = i[18];
  assign o[9648] = i[18];
  assign o[9649] = i[18];
  assign o[9650] = i[18];
  assign o[9651] = i[18];
  assign o[9652] = i[18];
  assign o[9653] = i[18];
  assign o[9654] = i[18];
  assign o[9655] = i[18];
  assign o[9656] = i[18];
  assign o[9657] = i[18];
  assign o[9658] = i[18];
  assign o[9659] = i[18];
  assign o[9660] = i[18];
  assign o[9661] = i[18];
  assign o[9662] = i[18];
  assign o[9663] = i[18];
  assign o[9664] = i[18];
  assign o[9665] = i[18];
  assign o[9666] = i[18];
  assign o[9667] = i[18];
  assign o[9668] = i[18];
  assign o[9669] = i[18];
  assign o[9670] = i[18];
  assign o[9671] = i[18];
  assign o[9672] = i[18];
  assign o[9673] = i[18];
  assign o[9674] = i[18];
  assign o[9675] = i[18];
  assign o[9676] = i[18];
  assign o[9677] = i[18];
  assign o[9678] = i[18];
  assign o[9679] = i[18];
  assign o[9680] = i[18];
  assign o[9681] = i[18];
  assign o[9682] = i[18];
  assign o[9683] = i[18];
  assign o[9684] = i[18];
  assign o[9685] = i[18];
  assign o[9686] = i[18];
  assign o[9687] = i[18];
  assign o[9688] = i[18];
  assign o[9689] = i[18];
  assign o[9690] = i[18];
  assign o[9691] = i[18];
  assign o[9692] = i[18];
  assign o[9693] = i[18];
  assign o[9694] = i[18];
  assign o[9695] = i[18];
  assign o[9696] = i[18];
  assign o[9697] = i[18];
  assign o[9698] = i[18];
  assign o[9699] = i[18];
  assign o[9700] = i[18];
  assign o[9701] = i[18];
  assign o[9702] = i[18];
  assign o[9703] = i[18];
  assign o[9704] = i[18];
  assign o[9705] = i[18];
  assign o[9706] = i[18];
  assign o[9707] = i[18];
  assign o[9708] = i[18];
  assign o[9709] = i[18];
  assign o[9710] = i[18];
  assign o[9711] = i[18];
  assign o[9712] = i[18];
  assign o[9713] = i[18];
  assign o[9714] = i[18];
  assign o[9715] = i[18];
  assign o[9716] = i[18];
  assign o[9717] = i[18];
  assign o[9718] = i[18];
  assign o[9719] = i[18];
  assign o[9720] = i[18];
  assign o[9721] = i[18];
  assign o[9722] = i[18];
  assign o[9723] = i[18];
  assign o[9724] = i[18];
  assign o[9725] = i[18];
  assign o[9726] = i[18];
  assign o[9727] = i[18];
  assign o[8704] = i[17];
  assign o[8705] = i[17];
  assign o[8706] = i[17];
  assign o[8707] = i[17];
  assign o[8708] = i[17];
  assign o[8709] = i[17];
  assign o[8710] = i[17];
  assign o[8711] = i[17];
  assign o[8712] = i[17];
  assign o[8713] = i[17];
  assign o[8714] = i[17];
  assign o[8715] = i[17];
  assign o[8716] = i[17];
  assign o[8717] = i[17];
  assign o[8718] = i[17];
  assign o[8719] = i[17];
  assign o[8720] = i[17];
  assign o[8721] = i[17];
  assign o[8722] = i[17];
  assign o[8723] = i[17];
  assign o[8724] = i[17];
  assign o[8725] = i[17];
  assign o[8726] = i[17];
  assign o[8727] = i[17];
  assign o[8728] = i[17];
  assign o[8729] = i[17];
  assign o[8730] = i[17];
  assign o[8731] = i[17];
  assign o[8732] = i[17];
  assign o[8733] = i[17];
  assign o[8734] = i[17];
  assign o[8735] = i[17];
  assign o[8736] = i[17];
  assign o[8737] = i[17];
  assign o[8738] = i[17];
  assign o[8739] = i[17];
  assign o[8740] = i[17];
  assign o[8741] = i[17];
  assign o[8742] = i[17];
  assign o[8743] = i[17];
  assign o[8744] = i[17];
  assign o[8745] = i[17];
  assign o[8746] = i[17];
  assign o[8747] = i[17];
  assign o[8748] = i[17];
  assign o[8749] = i[17];
  assign o[8750] = i[17];
  assign o[8751] = i[17];
  assign o[8752] = i[17];
  assign o[8753] = i[17];
  assign o[8754] = i[17];
  assign o[8755] = i[17];
  assign o[8756] = i[17];
  assign o[8757] = i[17];
  assign o[8758] = i[17];
  assign o[8759] = i[17];
  assign o[8760] = i[17];
  assign o[8761] = i[17];
  assign o[8762] = i[17];
  assign o[8763] = i[17];
  assign o[8764] = i[17];
  assign o[8765] = i[17];
  assign o[8766] = i[17];
  assign o[8767] = i[17];
  assign o[8768] = i[17];
  assign o[8769] = i[17];
  assign o[8770] = i[17];
  assign o[8771] = i[17];
  assign o[8772] = i[17];
  assign o[8773] = i[17];
  assign o[8774] = i[17];
  assign o[8775] = i[17];
  assign o[8776] = i[17];
  assign o[8777] = i[17];
  assign o[8778] = i[17];
  assign o[8779] = i[17];
  assign o[8780] = i[17];
  assign o[8781] = i[17];
  assign o[8782] = i[17];
  assign o[8783] = i[17];
  assign o[8784] = i[17];
  assign o[8785] = i[17];
  assign o[8786] = i[17];
  assign o[8787] = i[17];
  assign o[8788] = i[17];
  assign o[8789] = i[17];
  assign o[8790] = i[17];
  assign o[8791] = i[17];
  assign o[8792] = i[17];
  assign o[8793] = i[17];
  assign o[8794] = i[17];
  assign o[8795] = i[17];
  assign o[8796] = i[17];
  assign o[8797] = i[17];
  assign o[8798] = i[17];
  assign o[8799] = i[17];
  assign o[8800] = i[17];
  assign o[8801] = i[17];
  assign o[8802] = i[17];
  assign o[8803] = i[17];
  assign o[8804] = i[17];
  assign o[8805] = i[17];
  assign o[8806] = i[17];
  assign o[8807] = i[17];
  assign o[8808] = i[17];
  assign o[8809] = i[17];
  assign o[8810] = i[17];
  assign o[8811] = i[17];
  assign o[8812] = i[17];
  assign o[8813] = i[17];
  assign o[8814] = i[17];
  assign o[8815] = i[17];
  assign o[8816] = i[17];
  assign o[8817] = i[17];
  assign o[8818] = i[17];
  assign o[8819] = i[17];
  assign o[8820] = i[17];
  assign o[8821] = i[17];
  assign o[8822] = i[17];
  assign o[8823] = i[17];
  assign o[8824] = i[17];
  assign o[8825] = i[17];
  assign o[8826] = i[17];
  assign o[8827] = i[17];
  assign o[8828] = i[17];
  assign o[8829] = i[17];
  assign o[8830] = i[17];
  assign o[8831] = i[17];
  assign o[8832] = i[17];
  assign o[8833] = i[17];
  assign o[8834] = i[17];
  assign o[8835] = i[17];
  assign o[8836] = i[17];
  assign o[8837] = i[17];
  assign o[8838] = i[17];
  assign o[8839] = i[17];
  assign o[8840] = i[17];
  assign o[8841] = i[17];
  assign o[8842] = i[17];
  assign o[8843] = i[17];
  assign o[8844] = i[17];
  assign o[8845] = i[17];
  assign o[8846] = i[17];
  assign o[8847] = i[17];
  assign o[8848] = i[17];
  assign o[8849] = i[17];
  assign o[8850] = i[17];
  assign o[8851] = i[17];
  assign o[8852] = i[17];
  assign o[8853] = i[17];
  assign o[8854] = i[17];
  assign o[8855] = i[17];
  assign o[8856] = i[17];
  assign o[8857] = i[17];
  assign o[8858] = i[17];
  assign o[8859] = i[17];
  assign o[8860] = i[17];
  assign o[8861] = i[17];
  assign o[8862] = i[17];
  assign o[8863] = i[17];
  assign o[8864] = i[17];
  assign o[8865] = i[17];
  assign o[8866] = i[17];
  assign o[8867] = i[17];
  assign o[8868] = i[17];
  assign o[8869] = i[17];
  assign o[8870] = i[17];
  assign o[8871] = i[17];
  assign o[8872] = i[17];
  assign o[8873] = i[17];
  assign o[8874] = i[17];
  assign o[8875] = i[17];
  assign o[8876] = i[17];
  assign o[8877] = i[17];
  assign o[8878] = i[17];
  assign o[8879] = i[17];
  assign o[8880] = i[17];
  assign o[8881] = i[17];
  assign o[8882] = i[17];
  assign o[8883] = i[17];
  assign o[8884] = i[17];
  assign o[8885] = i[17];
  assign o[8886] = i[17];
  assign o[8887] = i[17];
  assign o[8888] = i[17];
  assign o[8889] = i[17];
  assign o[8890] = i[17];
  assign o[8891] = i[17];
  assign o[8892] = i[17];
  assign o[8893] = i[17];
  assign o[8894] = i[17];
  assign o[8895] = i[17];
  assign o[8896] = i[17];
  assign o[8897] = i[17];
  assign o[8898] = i[17];
  assign o[8899] = i[17];
  assign o[8900] = i[17];
  assign o[8901] = i[17];
  assign o[8902] = i[17];
  assign o[8903] = i[17];
  assign o[8904] = i[17];
  assign o[8905] = i[17];
  assign o[8906] = i[17];
  assign o[8907] = i[17];
  assign o[8908] = i[17];
  assign o[8909] = i[17];
  assign o[8910] = i[17];
  assign o[8911] = i[17];
  assign o[8912] = i[17];
  assign o[8913] = i[17];
  assign o[8914] = i[17];
  assign o[8915] = i[17];
  assign o[8916] = i[17];
  assign o[8917] = i[17];
  assign o[8918] = i[17];
  assign o[8919] = i[17];
  assign o[8920] = i[17];
  assign o[8921] = i[17];
  assign o[8922] = i[17];
  assign o[8923] = i[17];
  assign o[8924] = i[17];
  assign o[8925] = i[17];
  assign o[8926] = i[17];
  assign o[8927] = i[17];
  assign o[8928] = i[17];
  assign o[8929] = i[17];
  assign o[8930] = i[17];
  assign o[8931] = i[17];
  assign o[8932] = i[17];
  assign o[8933] = i[17];
  assign o[8934] = i[17];
  assign o[8935] = i[17];
  assign o[8936] = i[17];
  assign o[8937] = i[17];
  assign o[8938] = i[17];
  assign o[8939] = i[17];
  assign o[8940] = i[17];
  assign o[8941] = i[17];
  assign o[8942] = i[17];
  assign o[8943] = i[17];
  assign o[8944] = i[17];
  assign o[8945] = i[17];
  assign o[8946] = i[17];
  assign o[8947] = i[17];
  assign o[8948] = i[17];
  assign o[8949] = i[17];
  assign o[8950] = i[17];
  assign o[8951] = i[17];
  assign o[8952] = i[17];
  assign o[8953] = i[17];
  assign o[8954] = i[17];
  assign o[8955] = i[17];
  assign o[8956] = i[17];
  assign o[8957] = i[17];
  assign o[8958] = i[17];
  assign o[8959] = i[17];
  assign o[8960] = i[17];
  assign o[8961] = i[17];
  assign o[8962] = i[17];
  assign o[8963] = i[17];
  assign o[8964] = i[17];
  assign o[8965] = i[17];
  assign o[8966] = i[17];
  assign o[8967] = i[17];
  assign o[8968] = i[17];
  assign o[8969] = i[17];
  assign o[8970] = i[17];
  assign o[8971] = i[17];
  assign o[8972] = i[17];
  assign o[8973] = i[17];
  assign o[8974] = i[17];
  assign o[8975] = i[17];
  assign o[8976] = i[17];
  assign o[8977] = i[17];
  assign o[8978] = i[17];
  assign o[8979] = i[17];
  assign o[8980] = i[17];
  assign o[8981] = i[17];
  assign o[8982] = i[17];
  assign o[8983] = i[17];
  assign o[8984] = i[17];
  assign o[8985] = i[17];
  assign o[8986] = i[17];
  assign o[8987] = i[17];
  assign o[8988] = i[17];
  assign o[8989] = i[17];
  assign o[8990] = i[17];
  assign o[8991] = i[17];
  assign o[8992] = i[17];
  assign o[8993] = i[17];
  assign o[8994] = i[17];
  assign o[8995] = i[17];
  assign o[8996] = i[17];
  assign o[8997] = i[17];
  assign o[8998] = i[17];
  assign o[8999] = i[17];
  assign o[9000] = i[17];
  assign o[9001] = i[17];
  assign o[9002] = i[17];
  assign o[9003] = i[17];
  assign o[9004] = i[17];
  assign o[9005] = i[17];
  assign o[9006] = i[17];
  assign o[9007] = i[17];
  assign o[9008] = i[17];
  assign o[9009] = i[17];
  assign o[9010] = i[17];
  assign o[9011] = i[17];
  assign o[9012] = i[17];
  assign o[9013] = i[17];
  assign o[9014] = i[17];
  assign o[9015] = i[17];
  assign o[9016] = i[17];
  assign o[9017] = i[17];
  assign o[9018] = i[17];
  assign o[9019] = i[17];
  assign o[9020] = i[17];
  assign o[9021] = i[17];
  assign o[9022] = i[17];
  assign o[9023] = i[17];
  assign o[9024] = i[17];
  assign o[9025] = i[17];
  assign o[9026] = i[17];
  assign o[9027] = i[17];
  assign o[9028] = i[17];
  assign o[9029] = i[17];
  assign o[9030] = i[17];
  assign o[9031] = i[17];
  assign o[9032] = i[17];
  assign o[9033] = i[17];
  assign o[9034] = i[17];
  assign o[9035] = i[17];
  assign o[9036] = i[17];
  assign o[9037] = i[17];
  assign o[9038] = i[17];
  assign o[9039] = i[17];
  assign o[9040] = i[17];
  assign o[9041] = i[17];
  assign o[9042] = i[17];
  assign o[9043] = i[17];
  assign o[9044] = i[17];
  assign o[9045] = i[17];
  assign o[9046] = i[17];
  assign o[9047] = i[17];
  assign o[9048] = i[17];
  assign o[9049] = i[17];
  assign o[9050] = i[17];
  assign o[9051] = i[17];
  assign o[9052] = i[17];
  assign o[9053] = i[17];
  assign o[9054] = i[17];
  assign o[9055] = i[17];
  assign o[9056] = i[17];
  assign o[9057] = i[17];
  assign o[9058] = i[17];
  assign o[9059] = i[17];
  assign o[9060] = i[17];
  assign o[9061] = i[17];
  assign o[9062] = i[17];
  assign o[9063] = i[17];
  assign o[9064] = i[17];
  assign o[9065] = i[17];
  assign o[9066] = i[17];
  assign o[9067] = i[17];
  assign o[9068] = i[17];
  assign o[9069] = i[17];
  assign o[9070] = i[17];
  assign o[9071] = i[17];
  assign o[9072] = i[17];
  assign o[9073] = i[17];
  assign o[9074] = i[17];
  assign o[9075] = i[17];
  assign o[9076] = i[17];
  assign o[9077] = i[17];
  assign o[9078] = i[17];
  assign o[9079] = i[17];
  assign o[9080] = i[17];
  assign o[9081] = i[17];
  assign o[9082] = i[17];
  assign o[9083] = i[17];
  assign o[9084] = i[17];
  assign o[9085] = i[17];
  assign o[9086] = i[17];
  assign o[9087] = i[17];
  assign o[9088] = i[17];
  assign o[9089] = i[17];
  assign o[9090] = i[17];
  assign o[9091] = i[17];
  assign o[9092] = i[17];
  assign o[9093] = i[17];
  assign o[9094] = i[17];
  assign o[9095] = i[17];
  assign o[9096] = i[17];
  assign o[9097] = i[17];
  assign o[9098] = i[17];
  assign o[9099] = i[17];
  assign o[9100] = i[17];
  assign o[9101] = i[17];
  assign o[9102] = i[17];
  assign o[9103] = i[17];
  assign o[9104] = i[17];
  assign o[9105] = i[17];
  assign o[9106] = i[17];
  assign o[9107] = i[17];
  assign o[9108] = i[17];
  assign o[9109] = i[17];
  assign o[9110] = i[17];
  assign o[9111] = i[17];
  assign o[9112] = i[17];
  assign o[9113] = i[17];
  assign o[9114] = i[17];
  assign o[9115] = i[17];
  assign o[9116] = i[17];
  assign o[9117] = i[17];
  assign o[9118] = i[17];
  assign o[9119] = i[17];
  assign o[9120] = i[17];
  assign o[9121] = i[17];
  assign o[9122] = i[17];
  assign o[9123] = i[17];
  assign o[9124] = i[17];
  assign o[9125] = i[17];
  assign o[9126] = i[17];
  assign o[9127] = i[17];
  assign o[9128] = i[17];
  assign o[9129] = i[17];
  assign o[9130] = i[17];
  assign o[9131] = i[17];
  assign o[9132] = i[17];
  assign o[9133] = i[17];
  assign o[9134] = i[17];
  assign o[9135] = i[17];
  assign o[9136] = i[17];
  assign o[9137] = i[17];
  assign o[9138] = i[17];
  assign o[9139] = i[17];
  assign o[9140] = i[17];
  assign o[9141] = i[17];
  assign o[9142] = i[17];
  assign o[9143] = i[17];
  assign o[9144] = i[17];
  assign o[9145] = i[17];
  assign o[9146] = i[17];
  assign o[9147] = i[17];
  assign o[9148] = i[17];
  assign o[9149] = i[17];
  assign o[9150] = i[17];
  assign o[9151] = i[17];
  assign o[9152] = i[17];
  assign o[9153] = i[17];
  assign o[9154] = i[17];
  assign o[9155] = i[17];
  assign o[9156] = i[17];
  assign o[9157] = i[17];
  assign o[9158] = i[17];
  assign o[9159] = i[17];
  assign o[9160] = i[17];
  assign o[9161] = i[17];
  assign o[9162] = i[17];
  assign o[9163] = i[17];
  assign o[9164] = i[17];
  assign o[9165] = i[17];
  assign o[9166] = i[17];
  assign o[9167] = i[17];
  assign o[9168] = i[17];
  assign o[9169] = i[17];
  assign o[9170] = i[17];
  assign o[9171] = i[17];
  assign o[9172] = i[17];
  assign o[9173] = i[17];
  assign o[9174] = i[17];
  assign o[9175] = i[17];
  assign o[9176] = i[17];
  assign o[9177] = i[17];
  assign o[9178] = i[17];
  assign o[9179] = i[17];
  assign o[9180] = i[17];
  assign o[9181] = i[17];
  assign o[9182] = i[17];
  assign o[9183] = i[17];
  assign o[9184] = i[17];
  assign o[9185] = i[17];
  assign o[9186] = i[17];
  assign o[9187] = i[17];
  assign o[9188] = i[17];
  assign o[9189] = i[17];
  assign o[9190] = i[17];
  assign o[9191] = i[17];
  assign o[9192] = i[17];
  assign o[9193] = i[17];
  assign o[9194] = i[17];
  assign o[9195] = i[17];
  assign o[9196] = i[17];
  assign o[9197] = i[17];
  assign o[9198] = i[17];
  assign o[9199] = i[17];
  assign o[9200] = i[17];
  assign o[9201] = i[17];
  assign o[9202] = i[17];
  assign o[9203] = i[17];
  assign o[9204] = i[17];
  assign o[9205] = i[17];
  assign o[9206] = i[17];
  assign o[9207] = i[17];
  assign o[9208] = i[17];
  assign o[9209] = i[17];
  assign o[9210] = i[17];
  assign o[9211] = i[17];
  assign o[9212] = i[17];
  assign o[9213] = i[17];
  assign o[9214] = i[17];
  assign o[9215] = i[17];
  assign o[8192] = i[16];
  assign o[8193] = i[16];
  assign o[8194] = i[16];
  assign o[8195] = i[16];
  assign o[8196] = i[16];
  assign o[8197] = i[16];
  assign o[8198] = i[16];
  assign o[8199] = i[16];
  assign o[8200] = i[16];
  assign o[8201] = i[16];
  assign o[8202] = i[16];
  assign o[8203] = i[16];
  assign o[8204] = i[16];
  assign o[8205] = i[16];
  assign o[8206] = i[16];
  assign o[8207] = i[16];
  assign o[8208] = i[16];
  assign o[8209] = i[16];
  assign o[8210] = i[16];
  assign o[8211] = i[16];
  assign o[8212] = i[16];
  assign o[8213] = i[16];
  assign o[8214] = i[16];
  assign o[8215] = i[16];
  assign o[8216] = i[16];
  assign o[8217] = i[16];
  assign o[8218] = i[16];
  assign o[8219] = i[16];
  assign o[8220] = i[16];
  assign o[8221] = i[16];
  assign o[8222] = i[16];
  assign o[8223] = i[16];
  assign o[8224] = i[16];
  assign o[8225] = i[16];
  assign o[8226] = i[16];
  assign o[8227] = i[16];
  assign o[8228] = i[16];
  assign o[8229] = i[16];
  assign o[8230] = i[16];
  assign o[8231] = i[16];
  assign o[8232] = i[16];
  assign o[8233] = i[16];
  assign o[8234] = i[16];
  assign o[8235] = i[16];
  assign o[8236] = i[16];
  assign o[8237] = i[16];
  assign o[8238] = i[16];
  assign o[8239] = i[16];
  assign o[8240] = i[16];
  assign o[8241] = i[16];
  assign o[8242] = i[16];
  assign o[8243] = i[16];
  assign o[8244] = i[16];
  assign o[8245] = i[16];
  assign o[8246] = i[16];
  assign o[8247] = i[16];
  assign o[8248] = i[16];
  assign o[8249] = i[16];
  assign o[8250] = i[16];
  assign o[8251] = i[16];
  assign o[8252] = i[16];
  assign o[8253] = i[16];
  assign o[8254] = i[16];
  assign o[8255] = i[16];
  assign o[8256] = i[16];
  assign o[8257] = i[16];
  assign o[8258] = i[16];
  assign o[8259] = i[16];
  assign o[8260] = i[16];
  assign o[8261] = i[16];
  assign o[8262] = i[16];
  assign o[8263] = i[16];
  assign o[8264] = i[16];
  assign o[8265] = i[16];
  assign o[8266] = i[16];
  assign o[8267] = i[16];
  assign o[8268] = i[16];
  assign o[8269] = i[16];
  assign o[8270] = i[16];
  assign o[8271] = i[16];
  assign o[8272] = i[16];
  assign o[8273] = i[16];
  assign o[8274] = i[16];
  assign o[8275] = i[16];
  assign o[8276] = i[16];
  assign o[8277] = i[16];
  assign o[8278] = i[16];
  assign o[8279] = i[16];
  assign o[8280] = i[16];
  assign o[8281] = i[16];
  assign o[8282] = i[16];
  assign o[8283] = i[16];
  assign o[8284] = i[16];
  assign o[8285] = i[16];
  assign o[8286] = i[16];
  assign o[8287] = i[16];
  assign o[8288] = i[16];
  assign o[8289] = i[16];
  assign o[8290] = i[16];
  assign o[8291] = i[16];
  assign o[8292] = i[16];
  assign o[8293] = i[16];
  assign o[8294] = i[16];
  assign o[8295] = i[16];
  assign o[8296] = i[16];
  assign o[8297] = i[16];
  assign o[8298] = i[16];
  assign o[8299] = i[16];
  assign o[8300] = i[16];
  assign o[8301] = i[16];
  assign o[8302] = i[16];
  assign o[8303] = i[16];
  assign o[8304] = i[16];
  assign o[8305] = i[16];
  assign o[8306] = i[16];
  assign o[8307] = i[16];
  assign o[8308] = i[16];
  assign o[8309] = i[16];
  assign o[8310] = i[16];
  assign o[8311] = i[16];
  assign o[8312] = i[16];
  assign o[8313] = i[16];
  assign o[8314] = i[16];
  assign o[8315] = i[16];
  assign o[8316] = i[16];
  assign o[8317] = i[16];
  assign o[8318] = i[16];
  assign o[8319] = i[16];
  assign o[8320] = i[16];
  assign o[8321] = i[16];
  assign o[8322] = i[16];
  assign o[8323] = i[16];
  assign o[8324] = i[16];
  assign o[8325] = i[16];
  assign o[8326] = i[16];
  assign o[8327] = i[16];
  assign o[8328] = i[16];
  assign o[8329] = i[16];
  assign o[8330] = i[16];
  assign o[8331] = i[16];
  assign o[8332] = i[16];
  assign o[8333] = i[16];
  assign o[8334] = i[16];
  assign o[8335] = i[16];
  assign o[8336] = i[16];
  assign o[8337] = i[16];
  assign o[8338] = i[16];
  assign o[8339] = i[16];
  assign o[8340] = i[16];
  assign o[8341] = i[16];
  assign o[8342] = i[16];
  assign o[8343] = i[16];
  assign o[8344] = i[16];
  assign o[8345] = i[16];
  assign o[8346] = i[16];
  assign o[8347] = i[16];
  assign o[8348] = i[16];
  assign o[8349] = i[16];
  assign o[8350] = i[16];
  assign o[8351] = i[16];
  assign o[8352] = i[16];
  assign o[8353] = i[16];
  assign o[8354] = i[16];
  assign o[8355] = i[16];
  assign o[8356] = i[16];
  assign o[8357] = i[16];
  assign o[8358] = i[16];
  assign o[8359] = i[16];
  assign o[8360] = i[16];
  assign o[8361] = i[16];
  assign o[8362] = i[16];
  assign o[8363] = i[16];
  assign o[8364] = i[16];
  assign o[8365] = i[16];
  assign o[8366] = i[16];
  assign o[8367] = i[16];
  assign o[8368] = i[16];
  assign o[8369] = i[16];
  assign o[8370] = i[16];
  assign o[8371] = i[16];
  assign o[8372] = i[16];
  assign o[8373] = i[16];
  assign o[8374] = i[16];
  assign o[8375] = i[16];
  assign o[8376] = i[16];
  assign o[8377] = i[16];
  assign o[8378] = i[16];
  assign o[8379] = i[16];
  assign o[8380] = i[16];
  assign o[8381] = i[16];
  assign o[8382] = i[16];
  assign o[8383] = i[16];
  assign o[8384] = i[16];
  assign o[8385] = i[16];
  assign o[8386] = i[16];
  assign o[8387] = i[16];
  assign o[8388] = i[16];
  assign o[8389] = i[16];
  assign o[8390] = i[16];
  assign o[8391] = i[16];
  assign o[8392] = i[16];
  assign o[8393] = i[16];
  assign o[8394] = i[16];
  assign o[8395] = i[16];
  assign o[8396] = i[16];
  assign o[8397] = i[16];
  assign o[8398] = i[16];
  assign o[8399] = i[16];
  assign o[8400] = i[16];
  assign o[8401] = i[16];
  assign o[8402] = i[16];
  assign o[8403] = i[16];
  assign o[8404] = i[16];
  assign o[8405] = i[16];
  assign o[8406] = i[16];
  assign o[8407] = i[16];
  assign o[8408] = i[16];
  assign o[8409] = i[16];
  assign o[8410] = i[16];
  assign o[8411] = i[16];
  assign o[8412] = i[16];
  assign o[8413] = i[16];
  assign o[8414] = i[16];
  assign o[8415] = i[16];
  assign o[8416] = i[16];
  assign o[8417] = i[16];
  assign o[8418] = i[16];
  assign o[8419] = i[16];
  assign o[8420] = i[16];
  assign o[8421] = i[16];
  assign o[8422] = i[16];
  assign o[8423] = i[16];
  assign o[8424] = i[16];
  assign o[8425] = i[16];
  assign o[8426] = i[16];
  assign o[8427] = i[16];
  assign o[8428] = i[16];
  assign o[8429] = i[16];
  assign o[8430] = i[16];
  assign o[8431] = i[16];
  assign o[8432] = i[16];
  assign o[8433] = i[16];
  assign o[8434] = i[16];
  assign o[8435] = i[16];
  assign o[8436] = i[16];
  assign o[8437] = i[16];
  assign o[8438] = i[16];
  assign o[8439] = i[16];
  assign o[8440] = i[16];
  assign o[8441] = i[16];
  assign o[8442] = i[16];
  assign o[8443] = i[16];
  assign o[8444] = i[16];
  assign o[8445] = i[16];
  assign o[8446] = i[16];
  assign o[8447] = i[16];
  assign o[8448] = i[16];
  assign o[8449] = i[16];
  assign o[8450] = i[16];
  assign o[8451] = i[16];
  assign o[8452] = i[16];
  assign o[8453] = i[16];
  assign o[8454] = i[16];
  assign o[8455] = i[16];
  assign o[8456] = i[16];
  assign o[8457] = i[16];
  assign o[8458] = i[16];
  assign o[8459] = i[16];
  assign o[8460] = i[16];
  assign o[8461] = i[16];
  assign o[8462] = i[16];
  assign o[8463] = i[16];
  assign o[8464] = i[16];
  assign o[8465] = i[16];
  assign o[8466] = i[16];
  assign o[8467] = i[16];
  assign o[8468] = i[16];
  assign o[8469] = i[16];
  assign o[8470] = i[16];
  assign o[8471] = i[16];
  assign o[8472] = i[16];
  assign o[8473] = i[16];
  assign o[8474] = i[16];
  assign o[8475] = i[16];
  assign o[8476] = i[16];
  assign o[8477] = i[16];
  assign o[8478] = i[16];
  assign o[8479] = i[16];
  assign o[8480] = i[16];
  assign o[8481] = i[16];
  assign o[8482] = i[16];
  assign o[8483] = i[16];
  assign o[8484] = i[16];
  assign o[8485] = i[16];
  assign o[8486] = i[16];
  assign o[8487] = i[16];
  assign o[8488] = i[16];
  assign o[8489] = i[16];
  assign o[8490] = i[16];
  assign o[8491] = i[16];
  assign o[8492] = i[16];
  assign o[8493] = i[16];
  assign o[8494] = i[16];
  assign o[8495] = i[16];
  assign o[8496] = i[16];
  assign o[8497] = i[16];
  assign o[8498] = i[16];
  assign o[8499] = i[16];
  assign o[8500] = i[16];
  assign o[8501] = i[16];
  assign o[8502] = i[16];
  assign o[8503] = i[16];
  assign o[8504] = i[16];
  assign o[8505] = i[16];
  assign o[8506] = i[16];
  assign o[8507] = i[16];
  assign o[8508] = i[16];
  assign o[8509] = i[16];
  assign o[8510] = i[16];
  assign o[8511] = i[16];
  assign o[8512] = i[16];
  assign o[8513] = i[16];
  assign o[8514] = i[16];
  assign o[8515] = i[16];
  assign o[8516] = i[16];
  assign o[8517] = i[16];
  assign o[8518] = i[16];
  assign o[8519] = i[16];
  assign o[8520] = i[16];
  assign o[8521] = i[16];
  assign o[8522] = i[16];
  assign o[8523] = i[16];
  assign o[8524] = i[16];
  assign o[8525] = i[16];
  assign o[8526] = i[16];
  assign o[8527] = i[16];
  assign o[8528] = i[16];
  assign o[8529] = i[16];
  assign o[8530] = i[16];
  assign o[8531] = i[16];
  assign o[8532] = i[16];
  assign o[8533] = i[16];
  assign o[8534] = i[16];
  assign o[8535] = i[16];
  assign o[8536] = i[16];
  assign o[8537] = i[16];
  assign o[8538] = i[16];
  assign o[8539] = i[16];
  assign o[8540] = i[16];
  assign o[8541] = i[16];
  assign o[8542] = i[16];
  assign o[8543] = i[16];
  assign o[8544] = i[16];
  assign o[8545] = i[16];
  assign o[8546] = i[16];
  assign o[8547] = i[16];
  assign o[8548] = i[16];
  assign o[8549] = i[16];
  assign o[8550] = i[16];
  assign o[8551] = i[16];
  assign o[8552] = i[16];
  assign o[8553] = i[16];
  assign o[8554] = i[16];
  assign o[8555] = i[16];
  assign o[8556] = i[16];
  assign o[8557] = i[16];
  assign o[8558] = i[16];
  assign o[8559] = i[16];
  assign o[8560] = i[16];
  assign o[8561] = i[16];
  assign o[8562] = i[16];
  assign o[8563] = i[16];
  assign o[8564] = i[16];
  assign o[8565] = i[16];
  assign o[8566] = i[16];
  assign o[8567] = i[16];
  assign o[8568] = i[16];
  assign o[8569] = i[16];
  assign o[8570] = i[16];
  assign o[8571] = i[16];
  assign o[8572] = i[16];
  assign o[8573] = i[16];
  assign o[8574] = i[16];
  assign o[8575] = i[16];
  assign o[8576] = i[16];
  assign o[8577] = i[16];
  assign o[8578] = i[16];
  assign o[8579] = i[16];
  assign o[8580] = i[16];
  assign o[8581] = i[16];
  assign o[8582] = i[16];
  assign o[8583] = i[16];
  assign o[8584] = i[16];
  assign o[8585] = i[16];
  assign o[8586] = i[16];
  assign o[8587] = i[16];
  assign o[8588] = i[16];
  assign o[8589] = i[16];
  assign o[8590] = i[16];
  assign o[8591] = i[16];
  assign o[8592] = i[16];
  assign o[8593] = i[16];
  assign o[8594] = i[16];
  assign o[8595] = i[16];
  assign o[8596] = i[16];
  assign o[8597] = i[16];
  assign o[8598] = i[16];
  assign o[8599] = i[16];
  assign o[8600] = i[16];
  assign o[8601] = i[16];
  assign o[8602] = i[16];
  assign o[8603] = i[16];
  assign o[8604] = i[16];
  assign o[8605] = i[16];
  assign o[8606] = i[16];
  assign o[8607] = i[16];
  assign o[8608] = i[16];
  assign o[8609] = i[16];
  assign o[8610] = i[16];
  assign o[8611] = i[16];
  assign o[8612] = i[16];
  assign o[8613] = i[16];
  assign o[8614] = i[16];
  assign o[8615] = i[16];
  assign o[8616] = i[16];
  assign o[8617] = i[16];
  assign o[8618] = i[16];
  assign o[8619] = i[16];
  assign o[8620] = i[16];
  assign o[8621] = i[16];
  assign o[8622] = i[16];
  assign o[8623] = i[16];
  assign o[8624] = i[16];
  assign o[8625] = i[16];
  assign o[8626] = i[16];
  assign o[8627] = i[16];
  assign o[8628] = i[16];
  assign o[8629] = i[16];
  assign o[8630] = i[16];
  assign o[8631] = i[16];
  assign o[8632] = i[16];
  assign o[8633] = i[16];
  assign o[8634] = i[16];
  assign o[8635] = i[16];
  assign o[8636] = i[16];
  assign o[8637] = i[16];
  assign o[8638] = i[16];
  assign o[8639] = i[16];
  assign o[8640] = i[16];
  assign o[8641] = i[16];
  assign o[8642] = i[16];
  assign o[8643] = i[16];
  assign o[8644] = i[16];
  assign o[8645] = i[16];
  assign o[8646] = i[16];
  assign o[8647] = i[16];
  assign o[8648] = i[16];
  assign o[8649] = i[16];
  assign o[8650] = i[16];
  assign o[8651] = i[16];
  assign o[8652] = i[16];
  assign o[8653] = i[16];
  assign o[8654] = i[16];
  assign o[8655] = i[16];
  assign o[8656] = i[16];
  assign o[8657] = i[16];
  assign o[8658] = i[16];
  assign o[8659] = i[16];
  assign o[8660] = i[16];
  assign o[8661] = i[16];
  assign o[8662] = i[16];
  assign o[8663] = i[16];
  assign o[8664] = i[16];
  assign o[8665] = i[16];
  assign o[8666] = i[16];
  assign o[8667] = i[16];
  assign o[8668] = i[16];
  assign o[8669] = i[16];
  assign o[8670] = i[16];
  assign o[8671] = i[16];
  assign o[8672] = i[16];
  assign o[8673] = i[16];
  assign o[8674] = i[16];
  assign o[8675] = i[16];
  assign o[8676] = i[16];
  assign o[8677] = i[16];
  assign o[8678] = i[16];
  assign o[8679] = i[16];
  assign o[8680] = i[16];
  assign o[8681] = i[16];
  assign o[8682] = i[16];
  assign o[8683] = i[16];
  assign o[8684] = i[16];
  assign o[8685] = i[16];
  assign o[8686] = i[16];
  assign o[8687] = i[16];
  assign o[8688] = i[16];
  assign o[8689] = i[16];
  assign o[8690] = i[16];
  assign o[8691] = i[16];
  assign o[8692] = i[16];
  assign o[8693] = i[16];
  assign o[8694] = i[16];
  assign o[8695] = i[16];
  assign o[8696] = i[16];
  assign o[8697] = i[16];
  assign o[8698] = i[16];
  assign o[8699] = i[16];
  assign o[8700] = i[16];
  assign o[8701] = i[16];
  assign o[8702] = i[16];
  assign o[8703] = i[16];
  assign o[7680] = i[15];
  assign o[7681] = i[15];
  assign o[7682] = i[15];
  assign o[7683] = i[15];
  assign o[7684] = i[15];
  assign o[7685] = i[15];
  assign o[7686] = i[15];
  assign o[7687] = i[15];
  assign o[7688] = i[15];
  assign o[7689] = i[15];
  assign o[7690] = i[15];
  assign o[7691] = i[15];
  assign o[7692] = i[15];
  assign o[7693] = i[15];
  assign o[7694] = i[15];
  assign o[7695] = i[15];
  assign o[7696] = i[15];
  assign o[7697] = i[15];
  assign o[7698] = i[15];
  assign o[7699] = i[15];
  assign o[7700] = i[15];
  assign o[7701] = i[15];
  assign o[7702] = i[15];
  assign o[7703] = i[15];
  assign o[7704] = i[15];
  assign o[7705] = i[15];
  assign o[7706] = i[15];
  assign o[7707] = i[15];
  assign o[7708] = i[15];
  assign o[7709] = i[15];
  assign o[7710] = i[15];
  assign o[7711] = i[15];
  assign o[7712] = i[15];
  assign o[7713] = i[15];
  assign o[7714] = i[15];
  assign o[7715] = i[15];
  assign o[7716] = i[15];
  assign o[7717] = i[15];
  assign o[7718] = i[15];
  assign o[7719] = i[15];
  assign o[7720] = i[15];
  assign o[7721] = i[15];
  assign o[7722] = i[15];
  assign o[7723] = i[15];
  assign o[7724] = i[15];
  assign o[7725] = i[15];
  assign o[7726] = i[15];
  assign o[7727] = i[15];
  assign o[7728] = i[15];
  assign o[7729] = i[15];
  assign o[7730] = i[15];
  assign o[7731] = i[15];
  assign o[7732] = i[15];
  assign o[7733] = i[15];
  assign o[7734] = i[15];
  assign o[7735] = i[15];
  assign o[7736] = i[15];
  assign o[7737] = i[15];
  assign o[7738] = i[15];
  assign o[7739] = i[15];
  assign o[7740] = i[15];
  assign o[7741] = i[15];
  assign o[7742] = i[15];
  assign o[7743] = i[15];
  assign o[7744] = i[15];
  assign o[7745] = i[15];
  assign o[7746] = i[15];
  assign o[7747] = i[15];
  assign o[7748] = i[15];
  assign o[7749] = i[15];
  assign o[7750] = i[15];
  assign o[7751] = i[15];
  assign o[7752] = i[15];
  assign o[7753] = i[15];
  assign o[7754] = i[15];
  assign o[7755] = i[15];
  assign o[7756] = i[15];
  assign o[7757] = i[15];
  assign o[7758] = i[15];
  assign o[7759] = i[15];
  assign o[7760] = i[15];
  assign o[7761] = i[15];
  assign o[7762] = i[15];
  assign o[7763] = i[15];
  assign o[7764] = i[15];
  assign o[7765] = i[15];
  assign o[7766] = i[15];
  assign o[7767] = i[15];
  assign o[7768] = i[15];
  assign o[7769] = i[15];
  assign o[7770] = i[15];
  assign o[7771] = i[15];
  assign o[7772] = i[15];
  assign o[7773] = i[15];
  assign o[7774] = i[15];
  assign o[7775] = i[15];
  assign o[7776] = i[15];
  assign o[7777] = i[15];
  assign o[7778] = i[15];
  assign o[7779] = i[15];
  assign o[7780] = i[15];
  assign o[7781] = i[15];
  assign o[7782] = i[15];
  assign o[7783] = i[15];
  assign o[7784] = i[15];
  assign o[7785] = i[15];
  assign o[7786] = i[15];
  assign o[7787] = i[15];
  assign o[7788] = i[15];
  assign o[7789] = i[15];
  assign o[7790] = i[15];
  assign o[7791] = i[15];
  assign o[7792] = i[15];
  assign o[7793] = i[15];
  assign o[7794] = i[15];
  assign o[7795] = i[15];
  assign o[7796] = i[15];
  assign o[7797] = i[15];
  assign o[7798] = i[15];
  assign o[7799] = i[15];
  assign o[7800] = i[15];
  assign o[7801] = i[15];
  assign o[7802] = i[15];
  assign o[7803] = i[15];
  assign o[7804] = i[15];
  assign o[7805] = i[15];
  assign o[7806] = i[15];
  assign o[7807] = i[15];
  assign o[7808] = i[15];
  assign o[7809] = i[15];
  assign o[7810] = i[15];
  assign o[7811] = i[15];
  assign o[7812] = i[15];
  assign o[7813] = i[15];
  assign o[7814] = i[15];
  assign o[7815] = i[15];
  assign o[7816] = i[15];
  assign o[7817] = i[15];
  assign o[7818] = i[15];
  assign o[7819] = i[15];
  assign o[7820] = i[15];
  assign o[7821] = i[15];
  assign o[7822] = i[15];
  assign o[7823] = i[15];
  assign o[7824] = i[15];
  assign o[7825] = i[15];
  assign o[7826] = i[15];
  assign o[7827] = i[15];
  assign o[7828] = i[15];
  assign o[7829] = i[15];
  assign o[7830] = i[15];
  assign o[7831] = i[15];
  assign o[7832] = i[15];
  assign o[7833] = i[15];
  assign o[7834] = i[15];
  assign o[7835] = i[15];
  assign o[7836] = i[15];
  assign o[7837] = i[15];
  assign o[7838] = i[15];
  assign o[7839] = i[15];
  assign o[7840] = i[15];
  assign o[7841] = i[15];
  assign o[7842] = i[15];
  assign o[7843] = i[15];
  assign o[7844] = i[15];
  assign o[7845] = i[15];
  assign o[7846] = i[15];
  assign o[7847] = i[15];
  assign o[7848] = i[15];
  assign o[7849] = i[15];
  assign o[7850] = i[15];
  assign o[7851] = i[15];
  assign o[7852] = i[15];
  assign o[7853] = i[15];
  assign o[7854] = i[15];
  assign o[7855] = i[15];
  assign o[7856] = i[15];
  assign o[7857] = i[15];
  assign o[7858] = i[15];
  assign o[7859] = i[15];
  assign o[7860] = i[15];
  assign o[7861] = i[15];
  assign o[7862] = i[15];
  assign o[7863] = i[15];
  assign o[7864] = i[15];
  assign o[7865] = i[15];
  assign o[7866] = i[15];
  assign o[7867] = i[15];
  assign o[7868] = i[15];
  assign o[7869] = i[15];
  assign o[7870] = i[15];
  assign o[7871] = i[15];
  assign o[7872] = i[15];
  assign o[7873] = i[15];
  assign o[7874] = i[15];
  assign o[7875] = i[15];
  assign o[7876] = i[15];
  assign o[7877] = i[15];
  assign o[7878] = i[15];
  assign o[7879] = i[15];
  assign o[7880] = i[15];
  assign o[7881] = i[15];
  assign o[7882] = i[15];
  assign o[7883] = i[15];
  assign o[7884] = i[15];
  assign o[7885] = i[15];
  assign o[7886] = i[15];
  assign o[7887] = i[15];
  assign o[7888] = i[15];
  assign o[7889] = i[15];
  assign o[7890] = i[15];
  assign o[7891] = i[15];
  assign o[7892] = i[15];
  assign o[7893] = i[15];
  assign o[7894] = i[15];
  assign o[7895] = i[15];
  assign o[7896] = i[15];
  assign o[7897] = i[15];
  assign o[7898] = i[15];
  assign o[7899] = i[15];
  assign o[7900] = i[15];
  assign o[7901] = i[15];
  assign o[7902] = i[15];
  assign o[7903] = i[15];
  assign o[7904] = i[15];
  assign o[7905] = i[15];
  assign o[7906] = i[15];
  assign o[7907] = i[15];
  assign o[7908] = i[15];
  assign o[7909] = i[15];
  assign o[7910] = i[15];
  assign o[7911] = i[15];
  assign o[7912] = i[15];
  assign o[7913] = i[15];
  assign o[7914] = i[15];
  assign o[7915] = i[15];
  assign o[7916] = i[15];
  assign o[7917] = i[15];
  assign o[7918] = i[15];
  assign o[7919] = i[15];
  assign o[7920] = i[15];
  assign o[7921] = i[15];
  assign o[7922] = i[15];
  assign o[7923] = i[15];
  assign o[7924] = i[15];
  assign o[7925] = i[15];
  assign o[7926] = i[15];
  assign o[7927] = i[15];
  assign o[7928] = i[15];
  assign o[7929] = i[15];
  assign o[7930] = i[15];
  assign o[7931] = i[15];
  assign o[7932] = i[15];
  assign o[7933] = i[15];
  assign o[7934] = i[15];
  assign o[7935] = i[15];
  assign o[7936] = i[15];
  assign o[7937] = i[15];
  assign o[7938] = i[15];
  assign o[7939] = i[15];
  assign o[7940] = i[15];
  assign o[7941] = i[15];
  assign o[7942] = i[15];
  assign o[7943] = i[15];
  assign o[7944] = i[15];
  assign o[7945] = i[15];
  assign o[7946] = i[15];
  assign o[7947] = i[15];
  assign o[7948] = i[15];
  assign o[7949] = i[15];
  assign o[7950] = i[15];
  assign o[7951] = i[15];
  assign o[7952] = i[15];
  assign o[7953] = i[15];
  assign o[7954] = i[15];
  assign o[7955] = i[15];
  assign o[7956] = i[15];
  assign o[7957] = i[15];
  assign o[7958] = i[15];
  assign o[7959] = i[15];
  assign o[7960] = i[15];
  assign o[7961] = i[15];
  assign o[7962] = i[15];
  assign o[7963] = i[15];
  assign o[7964] = i[15];
  assign o[7965] = i[15];
  assign o[7966] = i[15];
  assign o[7967] = i[15];
  assign o[7968] = i[15];
  assign o[7969] = i[15];
  assign o[7970] = i[15];
  assign o[7971] = i[15];
  assign o[7972] = i[15];
  assign o[7973] = i[15];
  assign o[7974] = i[15];
  assign o[7975] = i[15];
  assign o[7976] = i[15];
  assign o[7977] = i[15];
  assign o[7978] = i[15];
  assign o[7979] = i[15];
  assign o[7980] = i[15];
  assign o[7981] = i[15];
  assign o[7982] = i[15];
  assign o[7983] = i[15];
  assign o[7984] = i[15];
  assign o[7985] = i[15];
  assign o[7986] = i[15];
  assign o[7987] = i[15];
  assign o[7988] = i[15];
  assign o[7989] = i[15];
  assign o[7990] = i[15];
  assign o[7991] = i[15];
  assign o[7992] = i[15];
  assign o[7993] = i[15];
  assign o[7994] = i[15];
  assign o[7995] = i[15];
  assign o[7996] = i[15];
  assign o[7997] = i[15];
  assign o[7998] = i[15];
  assign o[7999] = i[15];
  assign o[8000] = i[15];
  assign o[8001] = i[15];
  assign o[8002] = i[15];
  assign o[8003] = i[15];
  assign o[8004] = i[15];
  assign o[8005] = i[15];
  assign o[8006] = i[15];
  assign o[8007] = i[15];
  assign o[8008] = i[15];
  assign o[8009] = i[15];
  assign o[8010] = i[15];
  assign o[8011] = i[15];
  assign o[8012] = i[15];
  assign o[8013] = i[15];
  assign o[8014] = i[15];
  assign o[8015] = i[15];
  assign o[8016] = i[15];
  assign o[8017] = i[15];
  assign o[8018] = i[15];
  assign o[8019] = i[15];
  assign o[8020] = i[15];
  assign o[8021] = i[15];
  assign o[8022] = i[15];
  assign o[8023] = i[15];
  assign o[8024] = i[15];
  assign o[8025] = i[15];
  assign o[8026] = i[15];
  assign o[8027] = i[15];
  assign o[8028] = i[15];
  assign o[8029] = i[15];
  assign o[8030] = i[15];
  assign o[8031] = i[15];
  assign o[8032] = i[15];
  assign o[8033] = i[15];
  assign o[8034] = i[15];
  assign o[8035] = i[15];
  assign o[8036] = i[15];
  assign o[8037] = i[15];
  assign o[8038] = i[15];
  assign o[8039] = i[15];
  assign o[8040] = i[15];
  assign o[8041] = i[15];
  assign o[8042] = i[15];
  assign o[8043] = i[15];
  assign o[8044] = i[15];
  assign o[8045] = i[15];
  assign o[8046] = i[15];
  assign o[8047] = i[15];
  assign o[8048] = i[15];
  assign o[8049] = i[15];
  assign o[8050] = i[15];
  assign o[8051] = i[15];
  assign o[8052] = i[15];
  assign o[8053] = i[15];
  assign o[8054] = i[15];
  assign o[8055] = i[15];
  assign o[8056] = i[15];
  assign o[8057] = i[15];
  assign o[8058] = i[15];
  assign o[8059] = i[15];
  assign o[8060] = i[15];
  assign o[8061] = i[15];
  assign o[8062] = i[15];
  assign o[8063] = i[15];
  assign o[8064] = i[15];
  assign o[8065] = i[15];
  assign o[8066] = i[15];
  assign o[8067] = i[15];
  assign o[8068] = i[15];
  assign o[8069] = i[15];
  assign o[8070] = i[15];
  assign o[8071] = i[15];
  assign o[8072] = i[15];
  assign o[8073] = i[15];
  assign o[8074] = i[15];
  assign o[8075] = i[15];
  assign o[8076] = i[15];
  assign o[8077] = i[15];
  assign o[8078] = i[15];
  assign o[8079] = i[15];
  assign o[8080] = i[15];
  assign o[8081] = i[15];
  assign o[8082] = i[15];
  assign o[8083] = i[15];
  assign o[8084] = i[15];
  assign o[8085] = i[15];
  assign o[8086] = i[15];
  assign o[8087] = i[15];
  assign o[8088] = i[15];
  assign o[8089] = i[15];
  assign o[8090] = i[15];
  assign o[8091] = i[15];
  assign o[8092] = i[15];
  assign o[8093] = i[15];
  assign o[8094] = i[15];
  assign o[8095] = i[15];
  assign o[8096] = i[15];
  assign o[8097] = i[15];
  assign o[8098] = i[15];
  assign o[8099] = i[15];
  assign o[8100] = i[15];
  assign o[8101] = i[15];
  assign o[8102] = i[15];
  assign o[8103] = i[15];
  assign o[8104] = i[15];
  assign o[8105] = i[15];
  assign o[8106] = i[15];
  assign o[8107] = i[15];
  assign o[8108] = i[15];
  assign o[8109] = i[15];
  assign o[8110] = i[15];
  assign o[8111] = i[15];
  assign o[8112] = i[15];
  assign o[8113] = i[15];
  assign o[8114] = i[15];
  assign o[8115] = i[15];
  assign o[8116] = i[15];
  assign o[8117] = i[15];
  assign o[8118] = i[15];
  assign o[8119] = i[15];
  assign o[8120] = i[15];
  assign o[8121] = i[15];
  assign o[8122] = i[15];
  assign o[8123] = i[15];
  assign o[8124] = i[15];
  assign o[8125] = i[15];
  assign o[8126] = i[15];
  assign o[8127] = i[15];
  assign o[8128] = i[15];
  assign o[8129] = i[15];
  assign o[8130] = i[15];
  assign o[8131] = i[15];
  assign o[8132] = i[15];
  assign o[8133] = i[15];
  assign o[8134] = i[15];
  assign o[8135] = i[15];
  assign o[8136] = i[15];
  assign o[8137] = i[15];
  assign o[8138] = i[15];
  assign o[8139] = i[15];
  assign o[8140] = i[15];
  assign o[8141] = i[15];
  assign o[8142] = i[15];
  assign o[8143] = i[15];
  assign o[8144] = i[15];
  assign o[8145] = i[15];
  assign o[8146] = i[15];
  assign o[8147] = i[15];
  assign o[8148] = i[15];
  assign o[8149] = i[15];
  assign o[8150] = i[15];
  assign o[8151] = i[15];
  assign o[8152] = i[15];
  assign o[8153] = i[15];
  assign o[8154] = i[15];
  assign o[8155] = i[15];
  assign o[8156] = i[15];
  assign o[8157] = i[15];
  assign o[8158] = i[15];
  assign o[8159] = i[15];
  assign o[8160] = i[15];
  assign o[8161] = i[15];
  assign o[8162] = i[15];
  assign o[8163] = i[15];
  assign o[8164] = i[15];
  assign o[8165] = i[15];
  assign o[8166] = i[15];
  assign o[8167] = i[15];
  assign o[8168] = i[15];
  assign o[8169] = i[15];
  assign o[8170] = i[15];
  assign o[8171] = i[15];
  assign o[8172] = i[15];
  assign o[8173] = i[15];
  assign o[8174] = i[15];
  assign o[8175] = i[15];
  assign o[8176] = i[15];
  assign o[8177] = i[15];
  assign o[8178] = i[15];
  assign o[8179] = i[15];
  assign o[8180] = i[15];
  assign o[8181] = i[15];
  assign o[8182] = i[15];
  assign o[8183] = i[15];
  assign o[8184] = i[15];
  assign o[8185] = i[15];
  assign o[8186] = i[15];
  assign o[8187] = i[15];
  assign o[8188] = i[15];
  assign o[8189] = i[15];
  assign o[8190] = i[15];
  assign o[8191] = i[15];
  assign o[7168] = i[14];
  assign o[7169] = i[14];
  assign o[7170] = i[14];
  assign o[7171] = i[14];
  assign o[7172] = i[14];
  assign o[7173] = i[14];
  assign o[7174] = i[14];
  assign o[7175] = i[14];
  assign o[7176] = i[14];
  assign o[7177] = i[14];
  assign o[7178] = i[14];
  assign o[7179] = i[14];
  assign o[7180] = i[14];
  assign o[7181] = i[14];
  assign o[7182] = i[14];
  assign o[7183] = i[14];
  assign o[7184] = i[14];
  assign o[7185] = i[14];
  assign o[7186] = i[14];
  assign o[7187] = i[14];
  assign o[7188] = i[14];
  assign o[7189] = i[14];
  assign o[7190] = i[14];
  assign o[7191] = i[14];
  assign o[7192] = i[14];
  assign o[7193] = i[14];
  assign o[7194] = i[14];
  assign o[7195] = i[14];
  assign o[7196] = i[14];
  assign o[7197] = i[14];
  assign o[7198] = i[14];
  assign o[7199] = i[14];
  assign o[7200] = i[14];
  assign o[7201] = i[14];
  assign o[7202] = i[14];
  assign o[7203] = i[14];
  assign o[7204] = i[14];
  assign o[7205] = i[14];
  assign o[7206] = i[14];
  assign o[7207] = i[14];
  assign o[7208] = i[14];
  assign o[7209] = i[14];
  assign o[7210] = i[14];
  assign o[7211] = i[14];
  assign o[7212] = i[14];
  assign o[7213] = i[14];
  assign o[7214] = i[14];
  assign o[7215] = i[14];
  assign o[7216] = i[14];
  assign o[7217] = i[14];
  assign o[7218] = i[14];
  assign o[7219] = i[14];
  assign o[7220] = i[14];
  assign o[7221] = i[14];
  assign o[7222] = i[14];
  assign o[7223] = i[14];
  assign o[7224] = i[14];
  assign o[7225] = i[14];
  assign o[7226] = i[14];
  assign o[7227] = i[14];
  assign o[7228] = i[14];
  assign o[7229] = i[14];
  assign o[7230] = i[14];
  assign o[7231] = i[14];
  assign o[7232] = i[14];
  assign o[7233] = i[14];
  assign o[7234] = i[14];
  assign o[7235] = i[14];
  assign o[7236] = i[14];
  assign o[7237] = i[14];
  assign o[7238] = i[14];
  assign o[7239] = i[14];
  assign o[7240] = i[14];
  assign o[7241] = i[14];
  assign o[7242] = i[14];
  assign o[7243] = i[14];
  assign o[7244] = i[14];
  assign o[7245] = i[14];
  assign o[7246] = i[14];
  assign o[7247] = i[14];
  assign o[7248] = i[14];
  assign o[7249] = i[14];
  assign o[7250] = i[14];
  assign o[7251] = i[14];
  assign o[7252] = i[14];
  assign o[7253] = i[14];
  assign o[7254] = i[14];
  assign o[7255] = i[14];
  assign o[7256] = i[14];
  assign o[7257] = i[14];
  assign o[7258] = i[14];
  assign o[7259] = i[14];
  assign o[7260] = i[14];
  assign o[7261] = i[14];
  assign o[7262] = i[14];
  assign o[7263] = i[14];
  assign o[7264] = i[14];
  assign o[7265] = i[14];
  assign o[7266] = i[14];
  assign o[7267] = i[14];
  assign o[7268] = i[14];
  assign o[7269] = i[14];
  assign o[7270] = i[14];
  assign o[7271] = i[14];
  assign o[7272] = i[14];
  assign o[7273] = i[14];
  assign o[7274] = i[14];
  assign o[7275] = i[14];
  assign o[7276] = i[14];
  assign o[7277] = i[14];
  assign o[7278] = i[14];
  assign o[7279] = i[14];
  assign o[7280] = i[14];
  assign o[7281] = i[14];
  assign o[7282] = i[14];
  assign o[7283] = i[14];
  assign o[7284] = i[14];
  assign o[7285] = i[14];
  assign o[7286] = i[14];
  assign o[7287] = i[14];
  assign o[7288] = i[14];
  assign o[7289] = i[14];
  assign o[7290] = i[14];
  assign o[7291] = i[14];
  assign o[7292] = i[14];
  assign o[7293] = i[14];
  assign o[7294] = i[14];
  assign o[7295] = i[14];
  assign o[7296] = i[14];
  assign o[7297] = i[14];
  assign o[7298] = i[14];
  assign o[7299] = i[14];
  assign o[7300] = i[14];
  assign o[7301] = i[14];
  assign o[7302] = i[14];
  assign o[7303] = i[14];
  assign o[7304] = i[14];
  assign o[7305] = i[14];
  assign o[7306] = i[14];
  assign o[7307] = i[14];
  assign o[7308] = i[14];
  assign o[7309] = i[14];
  assign o[7310] = i[14];
  assign o[7311] = i[14];
  assign o[7312] = i[14];
  assign o[7313] = i[14];
  assign o[7314] = i[14];
  assign o[7315] = i[14];
  assign o[7316] = i[14];
  assign o[7317] = i[14];
  assign o[7318] = i[14];
  assign o[7319] = i[14];
  assign o[7320] = i[14];
  assign o[7321] = i[14];
  assign o[7322] = i[14];
  assign o[7323] = i[14];
  assign o[7324] = i[14];
  assign o[7325] = i[14];
  assign o[7326] = i[14];
  assign o[7327] = i[14];
  assign o[7328] = i[14];
  assign o[7329] = i[14];
  assign o[7330] = i[14];
  assign o[7331] = i[14];
  assign o[7332] = i[14];
  assign o[7333] = i[14];
  assign o[7334] = i[14];
  assign o[7335] = i[14];
  assign o[7336] = i[14];
  assign o[7337] = i[14];
  assign o[7338] = i[14];
  assign o[7339] = i[14];
  assign o[7340] = i[14];
  assign o[7341] = i[14];
  assign o[7342] = i[14];
  assign o[7343] = i[14];
  assign o[7344] = i[14];
  assign o[7345] = i[14];
  assign o[7346] = i[14];
  assign o[7347] = i[14];
  assign o[7348] = i[14];
  assign o[7349] = i[14];
  assign o[7350] = i[14];
  assign o[7351] = i[14];
  assign o[7352] = i[14];
  assign o[7353] = i[14];
  assign o[7354] = i[14];
  assign o[7355] = i[14];
  assign o[7356] = i[14];
  assign o[7357] = i[14];
  assign o[7358] = i[14];
  assign o[7359] = i[14];
  assign o[7360] = i[14];
  assign o[7361] = i[14];
  assign o[7362] = i[14];
  assign o[7363] = i[14];
  assign o[7364] = i[14];
  assign o[7365] = i[14];
  assign o[7366] = i[14];
  assign o[7367] = i[14];
  assign o[7368] = i[14];
  assign o[7369] = i[14];
  assign o[7370] = i[14];
  assign o[7371] = i[14];
  assign o[7372] = i[14];
  assign o[7373] = i[14];
  assign o[7374] = i[14];
  assign o[7375] = i[14];
  assign o[7376] = i[14];
  assign o[7377] = i[14];
  assign o[7378] = i[14];
  assign o[7379] = i[14];
  assign o[7380] = i[14];
  assign o[7381] = i[14];
  assign o[7382] = i[14];
  assign o[7383] = i[14];
  assign o[7384] = i[14];
  assign o[7385] = i[14];
  assign o[7386] = i[14];
  assign o[7387] = i[14];
  assign o[7388] = i[14];
  assign o[7389] = i[14];
  assign o[7390] = i[14];
  assign o[7391] = i[14];
  assign o[7392] = i[14];
  assign o[7393] = i[14];
  assign o[7394] = i[14];
  assign o[7395] = i[14];
  assign o[7396] = i[14];
  assign o[7397] = i[14];
  assign o[7398] = i[14];
  assign o[7399] = i[14];
  assign o[7400] = i[14];
  assign o[7401] = i[14];
  assign o[7402] = i[14];
  assign o[7403] = i[14];
  assign o[7404] = i[14];
  assign o[7405] = i[14];
  assign o[7406] = i[14];
  assign o[7407] = i[14];
  assign o[7408] = i[14];
  assign o[7409] = i[14];
  assign o[7410] = i[14];
  assign o[7411] = i[14];
  assign o[7412] = i[14];
  assign o[7413] = i[14];
  assign o[7414] = i[14];
  assign o[7415] = i[14];
  assign o[7416] = i[14];
  assign o[7417] = i[14];
  assign o[7418] = i[14];
  assign o[7419] = i[14];
  assign o[7420] = i[14];
  assign o[7421] = i[14];
  assign o[7422] = i[14];
  assign o[7423] = i[14];
  assign o[7424] = i[14];
  assign o[7425] = i[14];
  assign o[7426] = i[14];
  assign o[7427] = i[14];
  assign o[7428] = i[14];
  assign o[7429] = i[14];
  assign o[7430] = i[14];
  assign o[7431] = i[14];
  assign o[7432] = i[14];
  assign o[7433] = i[14];
  assign o[7434] = i[14];
  assign o[7435] = i[14];
  assign o[7436] = i[14];
  assign o[7437] = i[14];
  assign o[7438] = i[14];
  assign o[7439] = i[14];
  assign o[7440] = i[14];
  assign o[7441] = i[14];
  assign o[7442] = i[14];
  assign o[7443] = i[14];
  assign o[7444] = i[14];
  assign o[7445] = i[14];
  assign o[7446] = i[14];
  assign o[7447] = i[14];
  assign o[7448] = i[14];
  assign o[7449] = i[14];
  assign o[7450] = i[14];
  assign o[7451] = i[14];
  assign o[7452] = i[14];
  assign o[7453] = i[14];
  assign o[7454] = i[14];
  assign o[7455] = i[14];
  assign o[7456] = i[14];
  assign o[7457] = i[14];
  assign o[7458] = i[14];
  assign o[7459] = i[14];
  assign o[7460] = i[14];
  assign o[7461] = i[14];
  assign o[7462] = i[14];
  assign o[7463] = i[14];
  assign o[7464] = i[14];
  assign o[7465] = i[14];
  assign o[7466] = i[14];
  assign o[7467] = i[14];
  assign o[7468] = i[14];
  assign o[7469] = i[14];
  assign o[7470] = i[14];
  assign o[7471] = i[14];
  assign o[7472] = i[14];
  assign o[7473] = i[14];
  assign o[7474] = i[14];
  assign o[7475] = i[14];
  assign o[7476] = i[14];
  assign o[7477] = i[14];
  assign o[7478] = i[14];
  assign o[7479] = i[14];
  assign o[7480] = i[14];
  assign o[7481] = i[14];
  assign o[7482] = i[14];
  assign o[7483] = i[14];
  assign o[7484] = i[14];
  assign o[7485] = i[14];
  assign o[7486] = i[14];
  assign o[7487] = i[14];
  assign o[7488] = i[14];
  assign o[7489] = i[14];
  assign o[7490] = i[14];
  assign o[7491] = i[14];
  assign o[7492] = i[14];
  assign o[7493] = i[14];
  assign o[7494] = i[14];
  assign o[7495] = i[14];
  assign o[7496] = i[14];
  assign o[7497] = i[14];
  assign o[7498] = i[14];
  assign o[7499] = i[14];
  assign o[7500] = i[14];
  assign o[7501] = i[14];
  assign o[7502] = i[14];
  assign o[7503] = i[14];
  assign o[7504] = i[14];
  assign o[7505] = i[14];
  assign o[7506] = i[14];
  assign o[7507] = i[14];
  assign o[7508] = i[14];
  assign o[7509] = i[14];
  assign o[7510] = i[14];
  assign o[7511] = i[14];
  assign o[7512] = i[14];
  assign o[7513] = i[14];
  assign o[7514] = i[14];
  assign o[7515] = i[14];
  assign o[7516] = i[14];
  assign o[7517] = i[14];
  assign o[7518] = i[14];
  assign o[7519] = i[14];
  assign o[7520] = i[14];
  assign o[7521] = i[14];
  assign o[7522] = i[14];
  assign o[7523] = i[14];
  assign o[7524] = i[14];
  assign o[7525] = i[14];
  assign o[7526] = i[14];
  assign o[7527] = i[14];
  assign o[7528] = i[14];
  assign o[7529] = i[14];
  assign o[7530] = i[14];
  assign o[7531] = i[14];
  assign o[7532] = i[14];
  assign o[7533] = i[14];
  assign o[7534] = i[14];
  assign o[7535] = i[14];
  assign o[7536] = i[14];
  assign o[7537] = i[14];
  assign o[7538] = i[14];
  assign o[7539] = i[14];
  assign o[7540] = i[14];
  assign o[7541] = i[14];
  assign o[7542] = i[14];
  assign o[7543] = i[14];
  assign o[7544] = i[14];
  assign o[7545] = i[14];
  assign o[7546] = i[14];
  assign o[7547] = i[14];
  assign o[7548] = i[14];
  assign o[7549] = i[14];
  assign o[7550] = i[14];
  assign o[7551] = i[14];
  assign o[7552] = i[14];
  assign o[7553] = i[14];
  assign o[7554] = i[14];
  assign o[7555] = i[14];
  assign o[7556] = i[14];
  assign o[7557] = i[14];
  assign o[7558] = i[14];
  assign o[7559] = i[14];
  assign o[7560] = i[14];
  assign o[7561] = i[14];
  assign o[7562] = i[14];
  assign o[7563] = i[14];
  assign o[7564] = i[14];
  assign o[7565] = i[14];
  assign o[7566] = i[14];
  assign o[7567] = i[14];
  assign o[7568] = i[14];
  assign o[7569] = i[14];
  assign o[7570] = i[14];
  assign o[7571] = i[14];
  assign o[7572] = i[14];
  assign o[7573] = i[14];
  assign o[7574] = i[14];
  assign o[7575] = i[14];
  assign o[7576] = i[14];
  assign o[7577] = i[14];
  assign o[7578] = i[14];
  assign o[7579] = i[14];
  assign o[7580] = i[14];
  assign o[7581] = i[14];
  assign o[7582] = i[14];
  assign o[7583] = i[14];
  assign o[7584] = i[14];
  assign o[7585] = i[14];
  assign o[7586] = i[14];
  assign o[7587] = i[14];
  assign o[7588] = i[14];
  assign o[7589] = i[14];
  assign o[7590] = i[14];
  assign o[7591] = i[14];
  assign o[7592] = i[14];
  assign o[7593] = i[14];
  assign o[7594] = i[14];
  assign o[7595] = i[14];
  assign o[7596] = i[14];
  assign o[7597] = i[14];
  assign o[7598] = i[14];
  assign o[7599] = i[14];
  assign o[7600] = i[14];
  assign o[7601] = i[14];
  assign o[7602] = i[14];
  assign o[7603] = i[14];
  assign o[7604] = i[14];
  assign o[7605] = i[14];
  assign o[7606] = i[14];
  assign o[7607] = i[14];
  assign o[7608] = i[14];
  assign o[7609] = i[14];
  assign o[7610] = i[14];
  assign o[7611] = i[14];
  assign o[7612] = i[14];
  assign o[7613] = i[14];
  assign o[7614] = i[14];
  assign o[7615] = i[14];
  assign o[7616] = i[14];
  assign o[7617] = i[14];
  assign o[7618] = i[14];
  assign o[7619] = i[14];
  assign o[7620] = i[14];
  assign o[7621] = i[14];
  assign o[7622] = i[14];
  assign o[7623] = i[14];
  assign o[7624] = i[14];
  assign o[7625] = i[14];
  assign o[7626] = i[14];
  assign o[7627] = i[14];
  assign o[7628] = i[14];
  assign o[7629] = i[14];
  assign o[7630] = i[14];
  assign o[7631] = i[14];
  assign o[7632] = i[14];
  assign o[7633] = i[14];
  assign o[7634] = i[14];
  assign o[7635] = i[14];
  assign o[7636] = i[14];
  assign o[7637] = i[14];
  assign o[7638] = i[14];
  assign o[7639] = i[14];
  assign o[7640] = i[14];
  assign o[7641] = i[14];
  assign o[7642] = i[14];
  assign o[7643] = i[14];
  assign o[7644] = i[14];
  assign o[7645] = i[14];
  assign o[7646] = i[14];
  assign o[7647] = i[14];
  assign o[7648] = i[14];
  assign o[7649] = i[14];
  assign o[7650] = i[14];
  assign o[7651] = i[14];
  assign o[7652] = i[14];
  assign o[7653] = i[14];
  assign o[7654] = i[14];
  assign o[7655] = i[14];
  assign o[7656] = i[14];
  assign o[7657] = i[14];
  assign o[7658] = i[14];
  assign o[7659] = i[14];
  assign o[7660] = i[14];
  assign o[7661] = i[14];
  assign o[7662] = i[14];
  assign o[7663] = i[14];
  assign o[7664] = i[14];
  assign o[7665] = i[14];
  assign o[7666] = i[14];
  assign o[7667] = i[14];
  assign o[7668] = i[14];
  assign o[7669] = i[14];
  assign o[7670] = i[14];
  assign o[7671] = i[14];
  assign o[7672] = i[14];
  assign o[7673] = i[14];
  assign o[7674] = i[14];
  assign o[7675] = i[14];
  assign o[7676] = i[14];
  assign o[7677] = i[14];
  assign o[7678] = i[14];
  assign o[7679] = i[14];
  assign o[6656] = i[13];
  assign o[6657] = i[13];
  assign o[6658] = i[13];
  assign o[6659] = i[13];
  assign o[6660] = i[13];
  assign o[6661] = i[13];
  assign o[6662] = i[13];
  assign o[6663] = i[13];
  assign o[6664] = i[13];
  assign o[6665] = i[13];
  assign o[6666] = i[13];
  assign o[6667] = i[13];
  assign o[6668] = i[13];
  assign o[6669] = i[13];
  assign o[6670] = i[13];
  assign o[6671] = i[13];
  assign o[6672] = i[13];
  assign o[6673] = i[13];
  assign o[6674] = i[13];
  assign o[6675] = i[13];
  assign o[6676] = i[13];
  assign o[6677] = i[13];
  assign o[6678] = i[13];
  assign o[6679] = i[13];
  assign o[6680] = i[13];
  assign o[6681] = i[13];
  assign o[6682] = i[13];
  assign o[6683] = i[13];
  assign o[6684] = i[13];
  assign o[6685] = i[13];
  assign o[6686] = i[13];
  assign o[6687] = i[13];
  assign o[6688] = i[13];
  assign o[6689] = i[13];
  assign o[6690] = i[13];
  assign o[6691] = i[13];
  assign o[6692] = i[13];
  assign o[6693] = i[13];
  assign o[6694] = i[13];
  assign o[6695] = i[13];
  assign o[6696] = i[13];
  assign o[6697] = i[13];
  assign o[6698] = i[13];
  assign o[6699] = i[13];
  assign o[6700] = i[13];
  assign o[6701] = i[13];
  assign o[6702] = i[13];
  assign o[6703] = i[13];
  assign o[6704] = i[13];
  assign o[6705] = i[13];
  assign o[6706] = i[13];
  assign o[6707] = i[13];
  assign o[6708] = i[13];
  assign o[6709] = i[13];
  assign o[6710] = i[13];
  assign o[6711] = i[13];
  assign o[6712] = i[13];
  assign o[6713] = i[13];
  assign o[6714] = i[13];
  assign o[6715] = i[13];
  assign o[6716] = i[13];
  assign o[6717] = i[13];
  assign o[6718] = i[13];
  assign o[6719] = i[13];
  assign o[6720] = i[13];
  assign o[6721] = i[13];
  assign o[6722] = i[13];
  assign o[6723] = i[13];
  assign o[6724] = i[13];
  assign o[6725] = i[13];
  assign o[6726] = i[13];
  assign o[6727] = i[13];
  assign o[6728] = i[13];
  assign o[6729] = i[13];
  assign o[6730] = i[13];
  assign o[6731] = i[13];
  assign o[6732] = i[13];
  assign o[6733] = i[13];
  assign o[6734] = i[13];
  assign o[6735] = i[13];
  assign o[6736] = i[13];
  assign o[6737] = i[13];
  assign o[6738] = i[13];
  assign o[6739] = i[13];
  assign o[6740] = i[13];
  assign o[6741] = i[13];
  assign o[6742] = i[13];
  assign o[6743] = i[13];
  assign o[6744] = i[13];
  assign o[6745] = i[13];
  assign o[6746] = i[13];
  assign o[6747] = i[13];
  assign o[6748] = i[13];
  assign o[6749] = i[13];
  assign o[6750] = i[13];
  assign o[6751] = i[13];
  assign o[6752] = i[13];
  assign o[6753] = i[13];
  assign o[6754] = i[13];
  assign o[6755] = i[13];
  assign o[6756] = i[13];
  assign o[6757] = i[13];
  assign o[6758] = i[13];
  assign o[6759] = i[13];
  assign o[6760] = i[13];
  assign o[6761] = i[13];
  assign o[6762] = i[13];
  assign o[6763] = i[13];
  assign o[6764] = i[13];
  assign o[6765] = i[13];
  assign o[6766] = i[13];
  assign o[6767] = i[13];
  assign o[6768] = i[13];
  assign o[6769] = i[13];
  assign o[6770] = i[13];
  assign o[6771] = i[13];
  assign o[6772] = i[13];
  assign o[6773] = i[13];
  assign o[6774] = i[13];
  assign o[6775] = i[13];
  assign o[6776] = i[13];
  assign o[6777] = i[13];
  assign o[6778] = i[13];
  assign o[6779] = i[13];
  assign o[6780] = i[13];
  assign o[6781] = i[13];
  assign o[6782] = i[13];
  assign o[6783] = i[13];
  assign o[6784] = i[13];
  assign o[6785] = i[13];
  assign o[6786] = i[13];
  assign o[6787] = i[13];
  assign o[6788] = i[13];
  assign o[6789] = i[13];
  assign o[6790] = i[13];
  assign o[6791] = i[13];
  assign o[6792] = i[13];
  assign o[6793] = i[13];
  assign o[6794] = i[13];
  assign o[6795] = i[13];
  assign o[6796] = i[13];
  assign o[6797] = i[13];
  assign o[6798] = i[13];
  assign o[6799] = i[13];
  assign o[6800] = i[13];
  assign o[6801] = i[13];
  assign o[6802] = i[13];
  assign o[6803] = i[13];
  assign o[6804] = i[13];
  assign o[6805] = i[13];
  assign o[6806] = i[13];
  assign o[6807] = i[13];
  assign o[6808] = i[13];
  assign o[6809] = i[13];
  assign o[6810] = i[13];
  assign o[6811] = i[13];
  assign o[6812] = i[13];
  assign o[6813] = i[13];
  assign o[6814] = i[13];
  assign o[6815] = i[13];
  assign o[6816] = i[13];
  assign o[6817] = i[13];
  assign o[6818] = i[13];
  assign o[6819] = i[13];
  assign o[6820] = i[13];
  assign o[6821] = i[13];
  assign o[6822] = i[13];
  assign o[6823] = i[13];
  assign o[6824] = i[13];
  assign o[6825] = i[13];
  assign o[6826] = i[13];
  assign o[6827] = i[13];
  assign o[6828] = i[13];
  assign o[6829] = i[13];
  assign o[6830] = i[13];
  assign o[6831] = i[13];
  assign o[6832] = i[13];
  assign o[6833] = i[13];
  assign o[6834] = i[13];
  assign o[6835] = i[13];
  assign o[6836] = i[13];
  assign o[6837] = i[13];
  assign o[6838] = i[13];
  assign o[6839] = i[13];
  assign o[6840] = i[13];
  assign o[6841] = i[13];
  assign o[6842] = i[13];
  assign o[6843] = i[13];
  assign o[6844] = i[13];
  assign o[6845] = i[13];
  assign o[6846] = i[13];
  assign o[6847] = i[13];
  assign o[6848] = i[13];
  assign o[6849] = i[13];
  assign o[6850] = i[13];
  assign o[6851] = i[13];
  assign o[6852] = i[13];
  assign o[6853] = i[13];
  assign o[6854] = i[13];
  assign o[6855] = i[13];
  assign o[6856] = i[13];
  assign o[6857] = i[13];
  assign o[6858] = i[13];
  assign o[6859] = i[13];
  assign o[6860] = i[13];
  assign o[6861] = i[13];
  assign o[6862] = i[13];
  assign o[6863] = i[13];
  assign o[6864] = i[13];
  assign o[6865] = i[13];
  assign o[6866] = i[13];
  assign o[6867] = i[13];
  assign o[6868] = i[13];
  assign o[6869] = i[13];
  assign o[6870] = i[13];
  assign o[6871] = i[13];
  assign o[6872] = i[13];
  assign o[6873] = i[13];
  assign o[6874] = i[13];
  assign o[6875] = i[13];
  assign o[6876] = i[13];
  assign o[6877] = i[13];
  assign o[6878] = i[13];
  assign o[6879] = i[13];
  assign o[6880] = i[13];
  assign o[6881] = i[13];
  assign o[6882] = i[13];
  assign o[6883] = i[13];
  assign o[6884] = i[13];
  assign o[6885] = i[13];
  assign o[6886] = i[13];
  assign o[6887] = i[13];
  assign o[6888] = i[13];
  assign o[6889] = i[13];
  assign o[6890] = i[13];
  assign o[6891] = i[13];
  assign o[6892] = i[13];
  assign o[6893] = i[13];
  assign o[6894] = i[13];
  assign o[6895] = i[13];
  assign o[6896] = i[13];
  assign o[6897] = i[13];
  assign o[6898] = i[13];
  assign o[6899] = i[13];
  assign o[6900] = i[13];
  assign o[6901] = i[13];
  assign o[6902] = i[13];
  assign o[6903] = i[13];
  assign o[6904] = i[13];
  assign o[6905] = i[13];
  assign o[6906] = i[13];
  assign o[6907] = i[13];
  assign o[6908] = i[13];
  assign o[6909] = i[13];
  assign o[6910] = i[13];
  assign o[6911] = i[13];
  assign o[6912] = i[13];
  assign o[6913] = i[13];
  assign o[6914] = i[13];
  assign o[6915] = i[13];
  assign o[6916] = i[13];
  assign o[6917] = i[13];
  assign o[6918] = i[13];
  assign o[6919] = i[13];
  assign o[6920] = i[13];
  assign o[6921] = i[13];
  assign o[6922] = i[13];
  assign o[6923] = i[13];
  assign o[6924] = i[13];
  assign o[6925] = i[13];
  assign o[6926] = i[13];
  assign o[6927] = i[13];
  assign o[6928] = i[13];
  assign o[6929] = i[13];
  assign o[6930] = i[13];
  assign o[6931] = i[13];
  assign o[6932] = i[13];
  assign o[6933] = i[13];
  assign o[6934] = i[13];
  assign o[6935] = i[13];
  assign o[6936] = i[13];
  assign o[6937] = i[13];
  assign o[6938] = i[13];
  assign o[6939] = i[13];
  assign o[6940] = i[13];
  assign o[6941] = i[13];
  assign o[6942] = i[13];
  assign o[6943] = i[13];
  assign o[6944] = i[13];
  assign o[6945] = i[13];
  assign o[6946] = i[13];
  assign o[6947] = i[13];
  assign o[6948] = i[13];
  assign o[6949] = i[13];
  assign o[6950] = i[13];
  assign o[6951] = i[13];
  assign o[6952] = i[13];
  assign o[6953] = i[13];
  assign o[6954] = i[13];
  assign o[6955] = i[13];
  assign o[6956] = i[13];
  assign o[6957] = i[13];
  assign o[6958] = i[13];
  assign o[6959] = i[13];
  assign o[6960] = i[13];
  assign o[6961] = i[13];
  assign o[6962] = i[13];
  assign o[6963] = i[13];
  assign o[6964] = i[13];
  assign o[6965] = i[13];
  assign o[6966] = i[13];
  assign o[6967] = i[13];
  assign o[6968] = i[13];
  assign o[6969] = i[13];
  assign o[6970] = i[13];
  assign o[6971] = i[13];
  assign o[6972] = i[13];
  assign o[6973] = i[13];
  assign o[6974] = i[13];
  assign o[6975] = i[13];
  assign o[6976] = i[13];
  assign o[6977] = i[13];
  assign o[6978] = i[13];
  assign o[6979] = i[13];
  assign o[6980] = i[13];
  assign o[6981] = i[13];
  assign o[6982] = i[13];
  assign o[6983] = i[13];
  assign o[6984] = i[13];
  assign o[6985] = i[13];
  assign o[6986] = i[13];
  assign o[6987] = i[13];
  assign o[6988] = i[13];
  assign o[6989] = i[13];
  assign o[6990] = i[13];
  assign o[6991] = i[13];
  assign o[6992] = i[13];
  assign o[6993] = i[13];
  assign o[6994] = i[13];
  assign o[6995] = i[13];
  assign o[6996] = i[13];
  assign o[6997] = i[13];
  assign o[6998] = i[13];
  assign o[6999] = i[13];
  assign o[7000] = i[13];
  assign o[7001] = i[13];
  assign o[7002] = i[13];
  assign o[7003] = i[13];
  assign o[7004] = i[13];
  assign o[7005] = i[13];
  assign o[7006] = i[13];
  assign o[7007] = i[13];
  assign o[7008] = i[13];
  assign o[7009] = i[13];
  assign o[7010] = i[13];
  assign o[7011] = i[13];
  assign o[7012] = i[13];
  assign o[7013] = i[13];
  assign o[7014] = i[13];
  assign o[7015] = i[13];
  assign o[7016] = i[13];
  assign o[7017] = i[13];
  assign o[7018] = i[13];
  assign o[7019] = i[13];
  assign o[7020] = i[13];
  assign o[7021] = i[13];
  assign o[7022] = i[13];
  assign o[7023] = i[13];
  assign o[7024] = i[13];
  assign o[7025] = i[13];
  assign o[7026] = i[13];
  assign o[7027] = i[13];
  assign o[7028] = i[13];
  assign o[7029] = i[13];
  assign o[7030] = i[13];
  assign o[7031] = i[13];
  assign o[7032] = i[13];
  assign o[7033] = i[13];
  assign o[7034] = i[13];
  assign o[7035] = i[13];
  assign o[7036] = i[13];
  assign o[7037] = i[13];
  assign o[7038] = i[13];
  assign o[7039] = i[13];
  assign o[7040] = i[13];
  assign o[7041] = i[13];
  assign o[7042] = i[13];
  assign o[7043] = i[13];
  assign o[7044] = i[13];
  assign o[7045] = i[13];
  assign o[7046] = i[13];
  assign o[7047] = i[13];
  assign o[7048] = i[13];
  assign o[7049] = i[13];
  assign o[7050] = i[13];
  assign o[7051] = i[13];
  assign o[7052] = i[13];
  assign o[7053] = i[13];
  assign o[7054] = i[13];
  assign o[7055] = i[13];
  assign o[7056] = i[13];
  assign o[7057] = i[13];
  assign o[7058] = i[13];
  assign o[7059] = i[13];
  assign o[7060] = i[13];
  assign o[7061] = i[13];
  assign o[7062] = i[13];
  assign o[7063] = i[13];
  assign o[7064] = i[13];
  assign o[7065] = i[13];
  assign o[7066] = i[13];
  assign o[7067] = i[13];
  assign o[7068] = i[13];
  assign o[7069] = i[13];
  assign o[7070] = i[13];
  assign o[7071] = i[13];
  assign o[7072] = i[13];
  assign o[7073] = i[13];
  assign o[7074] = i[13];
  assign o[7075] = i[13];
  assign o[7076] = i[13];
  assign o[7077] = i[13];
  assign o[7078] = i[13];
  assign o[7079] = i[13];
  assign o[7080] = i[13];
  assign o[7081] = i[13];
  assign o[7082] = i[13];
  assign o[7083] = i[13];
  assign o[7084] = i[13];
  assign o[7085] = i[13];
  assign o[7086] = i[13];
  assign o[7087] = i[13];
  assign o[7088] = i[13];
  assign o[7089] = i[13];
  assign o[7090] = i[13];
  assign o[7091] = i[13];
  assign o[7092] = i[13];
  assign o[7093] = i[13];
  assign o[7094] = i[13];
  assign o[7095] = i[13];
  assign o[7096] = i[13];
  assign o[7097] = i[13];
  assign o[7098] = i[13];
  assign o[7099] = i[13];
  assign o[7100] = i[13];
  assign o[7101] = i[13];
  assign o[7102] = i[13];
  assign o[7103] = i[13];
  assign o[7104] = i[13];
  assign o[7105] = i[13];
  assign o[7106] = i[13];
  assign o[7107] = i[13];
  assign o[7108] = i[13];
  assign o[7109] = i[13];
  assign o[7110] = i[13];
  assign o[7111] = i[13];
  assign o[7112] = i[13];
  assign o[7113] = i[13];
  assign o[7114] = i[13];
  assign o[7115] = i[13];
  assign o[7116] = i[13];
  assign o[7117] = i[13];
  assign o[7118] = i[13];
  assign o[7119] = i[13];
  assign o[7120] = i[13];
  assign o[7121] = i[13];
  assign o[7122] = i[13];
  assign o[7123] = i[13];
  assign o[7124] = i[13];
  assign o[7125] = i[13];
  assign o[7126] = i[13];
  assign o[7127] = i[13];
  assign o[7128] = i[13];
  assign o[7129] = i[13];
  assign o[7130] = i[13];
  assign o[7131] = i[13];
  assign o[7132] = i[13];
  assign o[7133] = i[13];
  assign o[7134] = i[13];
  assign o[7135] = i[13];
  assign o[7136] = i[13];
  assign o[7137] = i[13];
  assign o[7138] = i[13];
  assign o[7139] = i[13];
  assign o[7140] = i[13];
  assign o[7141] = i[13];
  assign o[7142] = i[13];
  assign o[7143] = i[13];
  assign o[7144] = i[13];
  assign o[7145] = i[13];
  assign o[7146] = i[13];
  assign o[7147] = i[13];
  assign o[7148] = i[13];
  assign o[7149] = i[13];
  assign o[7150] = i[13];
  assign o[7151] = i[13];
  assign o[7152] = i[13];
  assign o[7153] = i[13];
  assign o[7154] = i[13];
  assign o[7155] = i[13];
  assign o[7156] = i[13];
  assign o[7157] = i[13];
  assign o[7158] = i[13];
  assign o[7159] = i[13];
  assign o[7160] = i[13];
  assign o[7161] = i[13];
  assign o[7162] = i[13];
  assign o[7163] = i[13];
  assign o[7164] = i[13];
  assign o[7165] = i[13];
  assign o[7166] = i[13];
  assign o[7167] = i[13];
  assign o[6144] = i[12];
  assign o[6145] = i[12];
  assign o[6146] = i[12];
  assign o[6147] = i[12];
  assign o[6148] = i[12];
  assign o[6149] = i[12];
  assign o[6150] = i[12];
  assign o[6151] = i[12];
  assign o[6152] = i[12];
  assign o[6153] = i[12];
  assign o[6154] = i[12];
  assign o[6155] = i[12];
  assign o[6156] = i[12];
  assign o[6157] = i[12];
  assign o[6158] = i[12];
  assign o[6159] = i[12];
  assign o[6160] = i[12];
  assign o[6161] = i[12];
  assign o[6162] = i[12];
  assign o[6163] = i[12];
  assign o[6164] = i[12];
  assign o[6165] = i[12];
  assign o[6166] = i[12];
  assign o[6167] = i[12];
  assign o[6168] = i[12];
  assign o[6169] = i[12];
  assign o[6170] = i[12];
  assign o[6171] = i[12];
  assign o[6172] = i[12];
  assign o[6173] = i[12];
  assign o[6174] = i[12];
  assign o[6175] = i[12];
  assign o[6176] = i[12];
  assign o[6177] = i[12];
  assign o[6178] = i[12];
  assign o[6179] = i[12];
  assign o[6180] = i[12];
  assign o[6181] = i[12];
  assign o[6182] = i[12];
  assign o[6183] = i[12];
  assign o[6184] = i[12];
  assign o[6185] = i[12];
  assign o[6186] = i[12];
  assign o[6187] = i[12];
  assign o[6188] = i[12];
  assign o[6189] = i[12];
  assign o[6190] = i[12];
  assign o[6191] = i[12];
  assign o[6192] = i[12];
  assign o[6193] = i[12];
  assign o[6194] = i[12];
  assign o[6195] = i[12];
  assign o[6196] = i[12];
  assign o[6197] = i[12];
  assign o[6198] = i[12];
  assign o[6199] = i[12];
  assign o[6200] = i[12];
  assign o[6201] = i[12];
  assign o[6202] = i[12];
  assign o[6203] = i[12];
  assign o[6204] = i[12];
  assign o[6205] = i[12];
  assign o[6206] = i[12];
  assign o[6207] = i[12];
  assign o[6208] = i[12];
  assign o[6209] = i[12];
  assign o[6210] = i[12];
  assign o[6211] = i[12];
  assign o[6212] = i[12];
  assign o[6213] = i[12];
  assign o[6214] = i[12];
  assign o[6215] = i[12];
  assign o[6216] = i[12];
  assign o[6217] = i[12];
  assign o[6218] = i[12];
  assign o[6219] = i[12];
  assign o[6220] = i[12];
  assign o[6221] = i[12];
  assign o[6222] = i[12];
  assign o[6223] = i[12];
  assign o[6224] = i[12];
  assign o[6225] = i[12];
  assign o[6226] = i[12];
  assign o[6227] = i[12];
  assign o[6228] = i[12];
  assign o[6229] = i[12];
  assign o[6230] = i[12];
  assign o[6231] = i[12];
  assign o[6232] = i[12];
  assign o[6233] = i[12];
  assign o[6234] = i[12];
  assign o[6235] = i[12];
  assign o[6236] = i[12];
  assign o[6237] = i[12];
  assign o[6238] = i[12];
  assign o[6239] = i[12];
  assign o[6240] = i[12];
  assign o[6241] = i[12];
  assign o[6242] = i[12];
  assign o[6243] = i[12];
  assign o[6244] = i[12];
  assign o[6245] = i[12];
  assign o[6246] = i[12];
  assign o[6247] = i[12];
  assign o[6248] = i[12];
  assign o[6249] = i[12];
  assign o[6250] = i[12];
  assign o[6251] = i[12];
  assign o[6252] = i[12];
  assign o[6253] = i[12];
  assign o[6254] = i[12];
  assign o[6255] = i[12];
  assign o[6256] = i[12];
  assign o[6257] = i[12];
  assign o[6258] = i[12];
  assign o[6259] = i[12];
  assign o[6260] = i[12];
  assign o[6261] = i[12];
  assign o[6262] = i[12];
  assign o[6263] = i[12];
  assign o[6264] = i[12];
  assign o[6265] = i[12];
  assign o[6266] = i[12];
  assign o[6267] = i[12];
  assign o[6268] = i[12];
  assign o[6269] = i[12];
  assign o[6270] = i[12];
  assign o[6271] = i[12];
  assign o[6272] = i[12];
  assign o[6273] = i[12];
  assign o[6274] = i[12];
  assign o[6275] = i[12];
  assign o[6276] = i[12];
  assign o[6277] = i[12];
  assign o[6278] = i[12];
  assign o[6279] = i[12];
  assign o[6280] = i[12];
  assign o[6281] = i[12];
  assign o[6282] = i[12];
  assign o[6283] = i[12];
  assign o[6284] = i[12];
  assign o[6285] = i[12];
  assign o[6286] = i[12];
  assign o[6287] = i[12];
  assign o[6288] = i[12];
  assign o[6289] = i[12];
  assign o[6290] = i[12];
  assign o[6291] = i[12];
  assign o[6292] = i[12];
  assign o[6293] = i[12];
  assign o[6294] = i[12];
  assign o[6295] = i[12];
  assign o[6296] = i[12];
  assign o[6297] = i[12];
  assign o[6298] = i[12];
  assign o[6299] = i[12];
  assign o[6300] = i[12];
  assign o[6301] = i[12];
  assign o[6302] = i[12];
  assign o[6303] = i[12];
  assign o[6304] = i[12];
  assign o[6305] = i[12];
  assign o[6306] = i[12];
  assign o[6307] = i[12];
  assign o[6308] = i[12];
  assign o[6309] = i[12];
  assign o[6310] = i[12];
  assign o[6311] = i[12];
  assign o[6312] = i[12];
  assign o[6313] = i[12];
  assign o[6314] = i[12];
  assign o[6315] = i[12];
  assign o[6316] = i[12];
  assign o[6317] = i[12];
  assign o[6318] = i[12];
  assign o[6319] = i[12];
  assign o[6320] = i[12];
  assign o[6321] = i[12];
  assign o[6322] = i[12];
  assign o[6323] = i[12];
  assign o[6324] = i[12];
  assign o[6325] = i[12];
  assign o[6326] = i[12];
  assign o[6327] = i[12];
  assign o[6328] = i[12];
  assign o[6329] = i[12];
  assign o[6330] = i[12];
  assign o[6331] = i[12];
  assign o[6332] = i[12];
  assign o[6333] = i[12];
  assign o[6334] = i[12];
  assign o[6335] = i[12];
  assign o[6336] = i[12];
  assign o[6337] = i[12];
  assign o[6338] = i[12];
  assign o[6339] = i[12];
  assign o[6340] = i[12];
  assign o[6341] = i[12];
  assign o[6342] = i[12];
  assign o[6343] = i[12];
  assign o[6344] = i[12];
  assign o[6345] = i[12];
  assign o[6346] = i[12];
  assign o[6347] = i[12];
  assign o[6348] = i[12];
  assign o[6349] = i[12];
  assign o[6350] = i[12];
  assign o[6351] = i[12];
  assign o[6352] = i[12];
  assign o[6353] = i[12];
  assign o[6354] = i[12];
  assign o[6355] = i[12];
  assign o[6356] = i[12];
  assign o[6357] = i[12];
  assign o[6358] = i[12];
  assign o[6359] = i[12];
  assign o[6360] = i[12];
  assign o[6361] = i[12];
  assign o[6362] = i[12];
  assign o[6363] = i[12];
  assign o[6364] = i[12];
  assign o[6365] = i[12];
  assign o[6366] = i[12];
  assign o[6367] = i[12];
  assign o[6368] = i[12];
  assign o[6369] = i[12];
  assign o[6370] = i[12];
  assign o[6371] = i[12];
  assign o[6372] = i[12];
  assign o[6373] = i[12];
  assign o[6374] = i[12];
  assign o[6375] = i[12];
  assign o[6376] = i[12];
  assign o[6377] = i[12];
  assign o[6378] = i[12];
  assign o[6379] = i[12];
  assign o[6380] = i[12];
  assign o[6381] = i[12];
  assign o[6382] = i[12];
  assign o[6383] = i[12];
  assign o[6384] = i[12];
  assign o[6385] = i[12];
  assign o[6386] = i[12];
  assign o[6387] = i[12];
  assign o[6388] = i[12];
  assign o[6389] = i[12];
  assign o[6390] = i[12];
  assign o[6391] = i[12];
  assign o[6392] = i[12];
  assign o[6393] = i[12];
  assign o[6394] = i[12];
  assign o[6395] = i[12];
  assign o[6396] = i[12];
  assign o[6397] = i[12];
  assign o[6398] = i[12];
  assign o[6399] = i[12];
  assign o[6400] = i[12];
  assign o[6401] = i[12];
  assign o[6402] = i[12];
  assign o[6403] = i[12];
  assign o[6404] = i[12];
  assign o[6405] = i[12];
  assign o[6406] = i[12];
  assign o[6407] = i[12];
  assign o[6408] = i[12];
  assign o[6409] = i[12];
  assign o[6410] = i[12];
  assign o[6411] = i[12];
  assign o[6412] = i[12];
  assign o[6413] = i[12];
  assign o[6414] = i[12];
  assign o[6415] = i[12];
  assign o[6416] = i[12];
  assign o[6417] = i[12];
  assign o[6418] = i[12];
  assign o[6419] = i[12];
  assign o[6420] = i[12];
  assign o[6421] = i[12];
  assign o[6422] = i[12];
  assign o[6423] = i[12];
  assign o[6424] = i[12];
  assign o[6425] = i[12];
  assign o[6426] = i[12];
  assign o[6427] = i[12];
  assign o[6428] = i[12];
  assign o[6429] = i[12];
  assign o[6430] = i[12];
  assign o[6431] = i[12];
  assign o[6432] = i[12];
  assign o[6433] = i[12];
  assign o[6434] = i[12];
  assign o[6435] = i[12];
  assign o[6436] = i[12];
  assign o[6437] = i[12];
  assign o[6438] = i[12];
  assign o[6439] = i[12];
  assign o[6440] = i[12];
  assign o[6441] = i[12];
  assign o[6442] = i[12];
  assign o[6443] = i[12];
  assign o[6444] = i[12];
  assign o[6445] = i[12];
  assign o[6446] = i[12];
  assign o[6447] = i[12];
  assign o[6448] = i[12];
  assign o[6449] = i[12];
  assign o[6450] = i[12];
  assign o[6451] = i[12];
  assign o[6452] = i[12];
  assign o[6453] = i[12];
  assign o[6454] = i[12];
  assign o[6455] = i[12];
  assign o[6456] = i[12];
  assign o[6457] = i[12];
  assign o[6458] = i[12];
  assign o[6459] = i[12];
  assign o[6460] = i[12];
  assign o[6461] = i[12];
  assign o[6462] = i[12];
  assign o[6463] = i[12];
  assign o[6464] = i[12];
  assign o[6465] = i[12];
  assign o[6466] = i[12];
  assign o[6467] = i[12];
  assign o[6468] = i[12];
  assign o[6469] = i[12];
  assign o[6470] = i[12];
  assign o[6471] = i[12];
  assign o[6472] = i[12];
  assign o[6473] = i[12];
  assign o[6474] = i[12];
  assign o[6475] = i[12];
  assign o[6476] = i[12];
  assign o[6477] = i[12];
  assign o[6478] = i[12];
  assign o[6479] = i[12];
  assign o[6480] = i[12];
  assign o[6481] = i[12];
  assign o[6482] = i[12];
  assign o[6483] = i[12];
  assign o[6484] = i[12];
  assign o[6485] = i[12];
  assign o[6486] = i[12];
  assign o[6487] = i[12];
  assign o[6488] = i[12];
  assign o[6489] = i[12];
  assign o[6490] = i[12];
  assign o[6491] = i[12];
  assign o[6492] = i[12];
  assign o[6493] = i[12];
  assign o[6494] = i[12];
  assign o[6495] = i[12];
  assign o[6496] = i[12];
  assign o[6497] = i[12];
  assign o[6498] = i[12];
  assign o[6499] = i[12];
  assign o[6500] = i[12];
  assign o[6501] = i[12];
  assign o[6502] = i[12];
  assign o[6503] = i[12];
  assign o[6504] = i[12];
  assign o[6505] = i[12];
  assign o[6506] = i[12];
  assign o[6507] = i[12];
  assign o[6508] = i[12];
  assign o[6509] = i[12];
  assign o[6510] = i[12];
  assign o[6511] = i[12];
  assign o[6512] = i[12];
  assign o[6513] = i[12];
  assign o[6514] = i[12];
  assign o[6515] = i[12];
  assign o[6516] = i[12];
  assign o[6517] = i[12];
  assign o[6518] = i[12];
  assign o[6519] = i[12];
  assign o[6520] = i[12];
  assign o[6521] = i[12];
  assign o[6522] = i[12];
  assign o[6523] = i[12];
  assign o[6524] = i[12];
  assign o[6525] = i[12];
  assign o[6526] = i[12];
  assign o[6527] = i[12];
  assign o[6528] = i[12];
  assign o[6529] = i[12];
  assign o[6530] = i[12];
  assign o[6531] = i[12];
  assign o[6532] = i[12];
  assign o[6533] = i[12];
  assign o[6534] = i[12];
  assign o[6535] = i[12];
  assign o[6536] = i[12];
  assign o[6537] = i[12];
  assign o[6538] = i[12];
  assign o[6539] = i[12];
  assign o[6540] = i[12];
  assign o[6541] = i[12];
  assign o[6542] = i[12];
  assign o[6543] = i[12];
  assign o[6544] = i[12];
  assign o[6545] = i[12];
  assign o[6546] = i[12];
  assign o[6547] = i[12];
  assign o[6548] = i[12];
  assign o[6549] = i[12];
  assign o[6550] = i[12];
  assign o[6551] = i[12];
  assign o[6552] = i[12];
  assign o[6553] = i[12];
  assign o[6554] = i[12];
  assign o[6555] = i[12];
  assign o[6556] = i[12];
  assign o[6557] = i[12];
  assign o[6558] = i[12];
  assign o[6559] = i[12];
  assign o[6560] = i[12];
  assign o[6561] = i[12];
  assign o[6562] = i[12];
  assign o[6563] = i[12];
  assign o[6564] = i[12];
  assign o[6565] = i[12];
  assign o[6566] = i[12];
  assign o[6567] = i[12];
  assign o[6568] = i[12];
  assign o[6569] = i[12];
  assign o[6570] = i[12];
  assign o[6571] = i[12];
  assign o[6572] = i[12];
  assign o[6573] = i[12];
  assign o[6574] = i[12];
  assign o[6575] = i[12];
  assign o[6576] = i[12];
  assign o[6577] = i[12];
  assign o[6578] = i[12];
  assign o[6579] = i[12];
  assign o[6580] = i[12];
  assign o[6581] = i[12];
  assign o[6582] = i[12];
  assign o[6583] = i[12];
  assign o[6584] = i[12];
  assign o[6585] = i[12];
  assign o[6586] = i[12];
  assign o[6587] = i[12];
  assign o[6588] = i[12];
  assign o[6589] = i[12];
  assign o[6590] = i[12];
  assign o[6591] = i[12];
  assign o[6592] = i[12];
  assign o[6593] = i[12];
  assign o[6594] = i[12];
  assign o[6595] = i[12];
  assign o[6596] = i[12];
  assign o[6597] = i[12];
  assign o[6598] = i[12];
  assign o[6599] = i[12];
  assign o[6600] = i[12];
  assign o[6601] = i[12];
  assign o[6602] = i[12];
  assign o[6603] = i[12];
  assign o[6604] = i[12];
  assign o[6605] = i[12];
  assign o[6606] = i[12];
  assign o[6607] = i[12];
  assign o[6608] = i[12];
  assign o[6609] = i[12];
  assign o[6610] = i[12];
  assign o[6611] = i[12];
  assign o[6612] = i[12];
  assign o[6613] = i[12];
  assign o[6614] = i[12];
  assign o[6615] = i[12];
  assign o[6616] = i[12];
  assign o[6617] = i[12];
  assign o[6618] = i[12];
  assign o[6619] = i[12];
  assign o[6620] = i[12];
  assign o[6621] = i[12];
  assign o[6622] = i[12];
  assign o[6623] = i[12];
  assign o[6624] = i[12];
  assign o[6625] = i[12];
  assign o[6626] = i[12];
  assign o[6627] = i[12];
  assign o[6628] = i[12];
  assign o[6629] = i[12];
  assign o[6630] = i[12];
  assign o[6631] = i[12];
  assign o[6632] = i[12];
  assign o[6633] = i[12];
  assign o[6634] = i[12];
  assign o[6635] = i[12];
  assign o[6636] = i[12];
  assign o[6637] = i[12];
  assign o[6638] = i[12];
  assign o[6639] = i[12];
  assign o[6640] = i[12];
  assign o[6641] = i[12];
  assign o[6642] = i[12];
  assign o[6643] = i[12];
  assign o[6644] = i[12];
  assign o[6645] = i[12];
  assign o[6646] = i[12];
  assign o[6647] = i[12];
  assign o[6648] = i[12];
  assign o[6649] = i[12];
  assign o[6650] = i[12];
  assign o[6651] = i[12];
  assign o[6652] = i[12];
  assign o[6653] = i[12];
  assign o[6654] = i[12];
  assign o[6655] = i[12];
  assign o[5632] = i[11];
  assign o[5633] = i[11];
  assign o[5634] = i[11];
  assign o[5635] = i[11];
  assign o[5636] = i[11];
  assign o[5637] = i[11];
  assign o[5638] = i[11];
  assign o[5639] = i[11];
  assign o[5640] = i[11];
  assign o[5641] = i[11];
  assign o[5642] = i[11];
  assign o[5643] = i[11];
  assign o[5644] = i[11];
  assign o[5645] = i[11];
  assign o[5646] = i[11];
  assign o[5647] = i[11];
  assign o[5648] = i[11];
  assign o[5649] = i[11];
  assign o[5650] = i[11];
  assign o[5651] = i[11];
  assign o[5652] = i[11];
  assign o[5653] = i[11];
  assign o[5654] = i[11];
  assign o[5655] = i[11];
  assign o[5656] = i[11];
  assign o[5657] = i[11];
  assign o[5658] = i[11];
  assign o[5659] = i[11];
  assign o[5660] = i[11];
  assign o[5661] = i[11];
  assign o[5662] = i[11];
  assign o[5663] = i[11];
  assign o[5664] = i[11];
  assign o[5665] = i[11];
  assign o[5666] = i[11];
  assign o[5667] = i[11];
  assign o[5668] = i[11];
  assign o[5669] = i[11];
  assign o[5670] = i[11];
  assign o[5671] = i[11];
  assign o[5672] = i[11];
  assign o[5673] = i[11];
  assign o[5674] = i[11];
  assign o[5675] = i[11];
  assign o[5676] = i[11];
  assign o[5677] = i[11];
  assign o[5678] = i[11];
  assign o[5679] = i[11];
  assign o[5680] = i[11];
  assign o[5681] = i[11];
  assign o[5682] = i[11];
  assign o[5683] = i[11];
  assign o[5684] = i[11];
  assign o[5685] = i[11];
  assign o[5686] = i[11];
  assign o[5687] = i[11];
  assign o[5688] = i[11];
  assign o[5689] = i[11];
  assign o[5690] = i[11];
  assign o[5691] = i[11];
  assign o[5692] = i[11];
  assign o[5693] = i[11];
  assign o[5694] = i[11];
  assign o[5695] = i[11];
  assign o[5696] = i[11];
  assign o[5697] = i[11];
  assign o[5698] = i[11];
  assign o[5699] = i[11];
  assign o[5700] = i[11];
  assign o[5701] = i[11];
  assign o[5702] = i[11];
  assign o[5703] = i[11];
  assign o[5704] = i[11];
  assign o[5705] = i[11];
  assign o[5706] = i[11];
  assign o[5707] = i[11];
  assign o[5708] = i[11];
  assign o[5709] = i[11];
  assign o[5710] = i[11];
  assign o[5711] = i[11];
  assign o[5712] = i[11];
  assign o[5713] = i[11];
  assign o[5714] = i[11];
  assign o[5715] = i[11];
  assign o[5716] = i[11];
  assign o[5717] = i[11];
  assign o[5718] = i[11];
  assign o[5719] = i[11];
  assign o[5720] = i[11];
  assign o[5721] = i[11];
  assign o[5722] = i[11];
  assign o[5723] = i[11];
  assign o[5724] = i[11];
  assign o[5725] = i[11];
  assign o[5726] = i[11];
  assign o[5727] = i[11];
  assign o[5728] = i[11];
  assign o[5729] = i[11];
  assign o[5730] = i[11];
  assign o[5731] = i[11];
  assign o[5732] = i[11];
  assign o[5733] = i[11];
  assign o[5734] = i[11];
  assign o[5735] = i[11];
  assign o[5736] = i[11];
  assign o[5737] = i[11];
  assign o[5738] = i[11];
  assign o[5739] = i[11];
  assign o[5740] = i[11];
  assign o[5741] = i[11];
  assign o[5742] = i[11];
  assign o[5743] = i[11];
  assign o[5744] = i[11];
  assign o[5745] = i[11];
  assign o[5746] = i[11];
  assign o[5747] = i[11];
  assign o[5748] = i[11];
  assign o[5749] = i[11];
  assign o[5750] = i[11];
  assign o[5751] = i[11];
  assign o[5752] = i[11];
  assign o[5753] = i[11];
  assign o[5754] = i[11];
  assign o[5755] = i[11];
  assign o[5756] = i[11];
  assign o[5757] = i[11];
  assign o[5758] = i[11];
  assign o[5759] = i[11];
  assign o[5760] = i[11];
  assign o[5761] = i[11];
  assign o[5762] = i[11];
  assign o[5763] = i[11];
  assign o[5764] = i[11];
  assign o[5765] = i[11];
  assign o[5766] = i[11];
  assign o[5767] = i[11];
  assign o[5768] = i[11];
  assign o[5769] = i[11];
  assign o[5770] = i[11];
  assign o[5771] = i[11];
  assign o[5772] = i[11];
  assign o[5773] = i[11];
  assign o[5774] = i[11];
  assign o[5775] = i[11];
  assign o[5776] = i[11];
  assign o[5777] = i[11];
  assign o[5778] = i[11];
  assign o[5779] = i[11];
  assign o[5780] = i[11];
  assign o[5781] = i[11];
  assign o[5782] = i[11];
  assign o[5783] = i[11];
  assign o[5784] = i[11];
  assign o[5785] = i[11];
  assign o[5786] = i[11];
  assign o[5787] = i[11];
  assign o[5788] = i[11];
  assign o[5789] = i[11];
  assign o[5790] = i[11];
  assign o[5791] = i[11];
  assign o[5792] = i[11];
  assign o[5793] = i[11];
  assign o[5794] = i[11];
  assign o[5795] = i[11];
  assign o[5796] = i[11];
  assign o[5797] = i[11];
  assign o[5798] = i[11];
  assign o[5799] = i[11];
  assign o[5800] = i[11];
  assign o[5801] = i[11];
  assign o[5802] = i[11];
  assign o[5803] = i[11];
  assign o[5804] = i[11];
  assign o[5805] = i[11];
  assign o[5806] = i[11];
  assign o[5807] = i[11];
  assign o[5808] = i[11];
  assign o[5809] = i[11];
  assign o[5810] = i[11];
  assign o[5811] = i[11];
  assign o[5812] = i[11];
  assign o[5813] = i[11];
  assign o[5814] = i[11];
  assign o[5815] = i[11];
  assign o[5816] = i[11];
  assign o[5817] = i[11];
  assign o[5818] = i[11];
  assign o[5819] = i[11];
  assign o[5820] = i[11];
  assign o[5821] = i[11];
  assign o[5822] = i[11];
  assign o[5823] = i[11];
  assign o[5824] = i[11];
  assign o[5825] = i[11];
  assign o[5826] = i[11];
  assign o[5827] = i[11];
  assign o[5828] = i[11];
  assign o[5829] = i[11];
  assign o[5830] = i[11];
  assign o[5831] = i[11];
  assign o[5832] = i[11];
  assign o[5833] = i[11];
  assign o[5834] = i[11];
  assign o[5835] = i[11];
  assign o[5836] = i[11];
  assign o[5837] = i[11];
  assign o[5838] = i[11];
  assign o[5839] = i[11];
  assign o[5840] = i[11];
  assign o[5841] = i[11];
  assign o[5842] = i[11];
  assign o[5843] = i[11];
  assign o[5844] = i[11];
  assign o[5845] = i[11];
  assign o[5846] = i[11];
  assign o[5847] = i[11];
  assign o[5848] = i[11];
  assign o[5849] = i[11];
  assign o[5850] = i[11];
  assign o[5851] = i[11];
  assign o[5852] = i[11];
  assign o[5853] = i[11];
  assign o[5854] = i[11];
  assign o[5855] = i[11];
  assign o[5856] = i[11];
  assign o[5857] = i[11];
  assign o[5858] = i[11];
  assign o[5859] = i[11];
  assign o[5860] = i[11];
  assign o[5861] = i[11];
  assign o[5862] = i[11];
  assign o[5863] = i[11];
  assign o[5864] = i[11];
  assign o[5865] = i[11];
  assign o[5866] = i[11];
  assign o[5867] = i[11];
  assign o[5868] = i[11];
  assign o[5869] = i[11];
  assign o[5870] = i[11];
  assign o[5871] = i[11];
  assign o[5872] = i[11];
  assign o[5873] = i[11];
  assign o[5874] = i[11];
  assign o[5875] = i[11];
  assign o[5876] = i[11];
  assign o[5877] = i[11];
  assign o[5878] = i[11];
  assign o[5879] = i[11];
  assign o[5880] = i[11];
  assign o[5881] = i[11];
  assign o[5882] = i[11];
  assign o[5883] = i[11];
  assign o[5884] = i[11];
  assign o[5885] = i[11];
  assign o[5886] = i[11];
  assign o[5887] = i[11];
  assign o[5888] = i[11];
  assign o[5889] = i[11];
  assign o[5890] = i[11];
  assign o[5891] = i[11];
  assign o[5892] = i[11];
  assign o[5893] = i[11];
  assign o[5894] = i[11];
  assign o[5895] = i[11];
  assign o[5896] = i[11];
  assign o[5897] = i[11];
  assign o[5898] = i[11];
  assign o[5899] = i[11];
  assign o[5900] = i[11];
  assign o[5901] = i[11];
  assign o[5902] = i[11];
  assign o[5903] = i[11];
  assign o[5904] = i[11];
  assign o[5905] = i[11];
  assign o[5906] = i[11];
  assign o[5907] = i[11];
  assign o[5908] = i[11];
  assign o[5909] = i[11];
  assign o[5910] = i[11];
  assign o[5911] = i[11];
  assign o[5912] = i[11];
  assign o[5913] = i[11];
  assign o[5914] = i[11];
  assign o[5915] = i[11];
  assign o[5916] = i[11];
  assign o[5917] = i[11];
  assign o[5918] = i[11];
  assign o[5919] = i[11];
  assign o[5920] = i[11];
  assign o[5921] = i[11];
  assign o[5922] = i[11];
  assign o[5923] = i[11];
  assign o[5924] = i[11];
  assign o[5925] = i[11];
  assign o[5926] = i[11];
  assign o[5927] = i[11];
  assign o[5928] = i[11];
  assign o[5929] = i[11];
  assign o[5930] = i[11];
  assign o[5931] = i[11];
  assign o[5932] = i[11];
  assign o[5933] = i[11];
  assign o[5934] = i[11];
  assign o[5935] = i[11];
  assign o[5936] = i[11];
  assign o[5937] = i[11];
  assign o[5938] = i[11];
  assign o[5939] = i[11];
  assign o[5940] = i[11];
  assign o[5941] = i[11];
  assign o[5942] = i[11];
  assign o[5943] = i[11];
  assign o[5944] = i[11];
  assign o[5945] = i[11];
  assign o[5946] = i[11];
  assign o[5947] = i[11];
  assign o[5948] = i[11];
  assign o[5949] = i[11];
  assign o[5950] = i[11];
  assign o[5951] = i[11];
  assign o[5952] = i[11];
  assign o[5953] = i[11];
  assign o[5954] = i[11];
  assign o[5955] = i[11];
  assign o[5956] = i[11];
  assign o[5957] = i[11];
  assign o[5958] = i[11];
  assign o[5959] = i[11];
  assign o[5960] = i[11];
  assign o[5961] = i[11];
  assign o[5962] = i[11];
  assign o[5963] = i[11];
  assign o[5964] = i[11];
  assign o[5965] = i[11];
  assign o[5966] = i[11];
  assign o[5967] = i[11];
  assign o[5968] = i[11];
  assign o[5969] = i[11];
  assign o[5970] = i[11];
  assign o[5971] = i[11];
  assign o[5972] = i[11];
  assign o[5973] = i[11];
  assign o[5974] = i[11];
  assign o[5975] = i[11];
  assign o[5976] = i[11];
  assign o[5977] = i[11];
  assign o[5978] = i[11];
  assign o[5979] = i[11];
  assign o[5980] = i[11];
  assign o[5981] = i[11];
  assign o[5982] = i[11];
  assign o[5983] = i[11];
  assign o[5984] = i[11];
  assign o[5985] = i[11];
  assign o[5986] = i[11];
  assign o[5987] = i[11];
  assign o[5988] = i[11];
  assign o[5989] = i[11];
  assign o[5990] = i[11];
  assign o[5991] = i[11];
  assign o[5992] = i[11];
  assign o[5993] = i[11];
  assign o[5994] = i[11];
  assign o[5995] = i[11];
  assign o[5996] = i[11];
  assign o[5997] = i[11];
  assign o[5998] = i[11];
  assign o[5999] = i[11];
  assign o[6000] = i[11];
  assign o[6001] = i[11];
  assign o[6002] = i[11];
  assign o[6003] = i[11];
  assign o[6004] = i[11];
  assign o[6005] = i[11];
  assign o[6006] = i[11];
  assign o[6007] = i[11];
  assign o[6008] = i[11];
  assign o[6009] = i[11];
  assign o[6010] = i[11];
  assign o[6011] = i[11];
  assign o[6012] = i[11];
  assign o[6013] = i[11];
  assign o[6014] = i[11];
  assign o[6015] = i[11];
  assign o[6016] = i[11];
  assign o[6017] = i[11];
  assign o[6018] = i[11];
  assign o[6019] = i[11];
  assign o[6020] = i[11];
  assign o[6021] = i[11];
  assign o[6022] = i[11];
  assign o[6023] = i[11];
  assign o[6024] = i[11];
  assign o[6025] = i[11];
  assign o[6026] = i[11];
  assign o[6027] = i[11];
  assign o[6028] = i[11];
  assign o[6029] = i[11];
  assign o[6030] = i[11];
  assign o[6031] = i[11];
  assign o[6032] = i[11];
  assign o[6033] = i[11];
  assign o[6034] = i[11];
  assign o[6035] = i[11];
  assign o[6036] = i[11];
  assign o[6037] = i[11];
  assign o[6038] = i[11];
  assign o[6039] = i[11];
  assign o[6040] = i[11];
  assign o[6041] = i[11];
  assign o[6042] = i[11];
  assign o[6043] = i[11];
  assign o[6044] = i[11];
  assign o[6045] = i[11];
  assign o[6046] = i[11];
  assign o[6047] = i[11];
  assign o[6048] = i[11];
  assign o[6049] = i[11];
  assign o[6050] = i[11];
  assign o[6051] = i[11];
  assign o[6052] = i[11];
  assign o[6053] = i[11];
  assign o[6054] = i[11];
  assign o[6055] = i[11];
  assign o[6056] = i[11];
  assign o[6057] = i[11];
  assign o[6058] = i[11];
  assign o[6059] = i[11];
  assign o[6060] = i[11];
  assign o[6061] = i[11];
  assign o[6062] = i[11];
  assign o[6063] = i[11];
  assign o[6064] = i[11];
  assign o[6065] = i[11];
  assign o[6066] = i[11];
  assign o[6067] = i[11];
  assign o[6068] = i[11];
  assign o[6069] = i[11];
  assign o[6070] = i[11];
  assign o[6071] = i[11];
  assign o[6072] = i[11];
  assign o[6073] = i[11];
  assign o[6074] = i[11];
  assign o[6075] = i[11];
  assign o[6076] = i[11];
  assign o[6077] = i[11];
  assign o[6078] = i[11];
  assign o[6079] = i[11];
  assign o[6080] = i[11];
  assign o[6081] = i[11];
  assign o[6082] = i[11];
  assign o[6083] = i[11];
  assign o[6084] = i[11];
  assign o[6085] = i[11];
  assign o[6086] = i[11];
  assign o[6087] = i[11];
  assign o[6088] = i[11];
  assign o[6089] = i[11];
  assign o[6090] = i[11];
  assign o[6091] = i[11];
  assign o[6092] = i[11];
  assign o[6093] = i[11];
  assign o[6094] = i[11];
  assign o[6095] = i[11];
  assign o[6096] = i[11];
  assign o[6097] = i[11];
  assign o[6098] = i[11];
  assign o[6099] = i[11];
  assign o[6100] = i[11];
  assign o[6101] = i[11];
  assign o[6102] = i[11];
  assign o[6103] = i[11];
  assign o[6104] = i[11];
  assign o[6105] = i[11];
  assign o[6106] = i[11];
  assign o[6107] = i[11];
  assign o[6108] = i[11];
  assign o[6109] = i[11];
  assign o[6110] = i[11];
  assign o[6111] = i[11];
  assign o[6112] = i[11];
  assign o[6113] = i[11];
  assign o[6114] = i[11];
  assign o[6115] = i[11];
  assign o[6116] = i[11];
  assign o[6117] = i[11];
  assign o[6118] = i[11];
  assign o[6119] = i[11];
  assign o[6120] = i[11];
  assign o[6121] = i[11];
  assign o[6122] = i[11];
  assign o[6123] = i[11];
  assign o[6124] = i[11];
  assign o[6125] = i[11];
  assign o[6126] = i[11];
  assign o[6127] = i[11];
  assign o[6128] = i[11];
  assign o[6129] = i[11];
  assign o[6130] = i[11];
  assign o[6131] = i[11];
  assign o[6132] = i[11];
  assign o[6133] = i[11];
  assign o[6134] = i[11];
  assign o[6135] = i[11];
  assign o[6136] = i[11];
  assign o[6137] = i[11];
  assign o[6138] = i[11];
  assign o[6139] = i[11];
  assign o[6140] = i[11];
  assign o[6141] = i[11];
  assign o[6142] = i[11];
  assign o[6143] = i[11];
  assign o[5120] = i[10];
  assign o[5121] = i[10];
  assign o[5122] = i[10];
  assign o[5123] = i[10];
  assign o[5124] = i[10];
  assign o[5125] = i[10];
  assign o[5126] = i[10];
  assign o[5127] = i[10];
  assign o[5128] = i[10];
  assign o[5129] = i[10];
  assign o[5130] = i[10];
  assign o[5131] = i[10];
  assign o[5132] = i[10];
  assign o[5133] = i[10];
  assign o[5134] = i[10];
  assign o[5135] = i[10];
  assign o[5136] = i[10];
  assign o[5137] = i[10];
  assign o[5138] = i[10];
  assign o[5139] = i[10];
  assign o[5140] = i[10];
  assign o[5141] = i[10];
  assign o[5142] = i[10];
  assign o[5143] = i[10];
  assign o[5144] = i[10];
  assign o[5145] = i[10];
  assign o[5146] = i[10];
  assign o[5147] = i[10];
  assign o[5148] = i[10];
  assign o[5149] = i[10];
  assign o[5150] = i[10];
  assign o[5151] = i[10];
  assign o[5152] = i[10];
  assign o[5153] = i[10];
  assign o[5154] = i[10];
  assign o[5155] = i[10];
  assign o[5156] = i[10];
  assign o[5157] = i[10];
  assign o[5158] = i[10];
  assign o[5159] = i[10];
  assign o[5160] = i[10];
  assign o[5161] = i[10];
  assign o[5162] = i[10];
  assign o[5163] = i[10];
  assign o[5164] = i[10];
  assign o[5165] = i[10];
  assign o[5166] = i[10];
  assign o[5167] = i[10];
  assign o[5168] = i[10];
  assign o[5169] = i[10];
  assign o[5170] = i[10];
  assign o[5171] = i[10];
  assign o[5172] = i[10];
  assign o[5173] = i[10];
  assign o[5174] = i[10];
  assign o[5175] = i[10];
  assign o[5176] = i[10];
  assign o[5177] = i[10];
  assign o[5178] = i[10];
  assign o[5179] = i[10];
  assign o[5180] = i[10];
  assign o[5181] = i[10];
  assign o[5182] = i[10];
  assign o[5183] = i[10];
  assign o[5184] = i[10];
  assign o[5185] = i[10];
  assign o[5186] = i[10];
  assign o[5187] = i[10];
  assign o[5188] = i[10];
  assign o[5189] = i[10];
  assign o[5190] = i[10];
  assign o[5191] = i[10];
  assign o[5192] = i[10];
  assign o[5193] = i[10];
  assign o[5194] = i[10];
  assign o[5195] = i[10];
  assign o[5196] = i[10];
  assign o[5197] = i[10];
  assign o[5198] = i[10];
  assign o[5199] = i[10];
  assign o[5200] = i[10];
  assign o[5201] = i[10];
  assign o[5202] = i[10];
  assign o[5203] = i[10];
  assign o[5204] = i[10];
  assign o[5205] = i[10];
  assign o[5206] = i[10];
  assign o[5207] = i[10];
  assign o[5208] = i[10];
  assign o[5209] = i[10];
  assign o[5210] = i[10];
  assign o[5211] = i[10];
  assign o[5212] = i[10];
  assign o[5213] = i[10];
  assign o[5214] = i[10];
  assign o[5215] = i[10];
  assign o[5216] = i[10];
  assign o[5217] = i[10];
  assign o[5218] = i[10];
  assign o[5219] = i[10];
  assign o[5220] = i[10];
  assign o[5221] = i[10];
  assign o[5222] = i[10];
  assign o[5223] = i[10];
  assign o[5224] = i[10];
  assign o[5225] = i[10];
  assign o[5226] = i[10];
  assign o[5227] = i[10];
  assign o[5228] = i[10];
  assign o[5229] = i[10];
  assign o[5230] = i[10];
  assign o[5231] = i[10];
  assign o[5232] = i[10];
  assign o[5233] = i[10];
  assign o[5234] = i[10];
  assign o[5235] = i[10];
  assign o[5236] = i[10];
  assign o[5237] = i[10];
  assign o[5238] = i[10];
  assign o[5239] = i[10];
  assign o[5240] = i[10];
  assign o[5241] = i[10];
  assign o[5242] = i[10];
  assign o[5243] = i[10];
  assign o[5244] = i[10];
  assign o[5245] = i[10];
  assign o[5246] = i[10];
  assign o[5247] = i[10];
  assign o[5248] = i[10];
  assign o[5249] = i[10];
  assign o[5250] = i[10];
  assign o[5251] = i[10];
  assign o[5252] = i[10];
  assign o[5253] = i[10];
  assign o[5254] = i[10];
  assign o[5255] = i[10];
  assign o[5256] = i[10];
  assign o[5257] = i[10];
  assign o[5258] = i[10];
  assign o[5259] = i[10];
  assign o[5260] = i[10];
  assign o[5261] = i[10];
  assign o[5262] = i[10];
  assign o[5263] = i[10];
  assign o[5264] = i[10];
  assign o[5265] = i[10];
  assign o[5266] = i[10];
  assign o[5267] = i[10];
  assign o[5268] = i[10];
  assign o[5269] = i[10];
  assign o[5270] = i[10];
  assign o[5271] = i[10];
  assign o[5272] = i[10];
  assign o[5273] = i[10];
  assign o[5274] = i[10];
  assign o[5275] = i[10];
  assign o[5276] = i[10];
  assign o[5277] = i[10];
  assign o[5278] = i[10];
  assign o[5279] = i[10];
  assign o[5280] = i[10];
  assign o[5281] = i[10];
  assign o[5282] = i[10];
  assign o[5283] = i[10];
  assign o[5284] = i[10];
  assign o[5285] = i[10];
  assign o[5286] = i[10];
  assign o[5287] = i[10];
  assign o[5288] = i[10];
  assign o[5289] = i[10];
  assign o[5290] = i[10];
  assign o[5291] = i[10];
  assign o[5292] = i[10];
  assign o[5293] = i[10];
  assign o[5294] = i[10];
  assign o[5295] = i[10];
  assign o[5296] = i[10];
  assign o[5297] = i[10];
  assign o[5298] = i[10];
  assign o[5299] = i[10];
  assign o[5300] = i[10];
  assign o[5301] = i[10];
  assign o[5302] = i[10];
  assign o[5303] = i[10];
  assign o[5304] = i[10];
  assign o[5305] = i[10];
  assign o[5306] = i[10];
  assign o[5307] = i[10];
  assign o[5308] = i[10];
  assign o[5309] = i[10];
  assign o[5310] = i[10];
  assign o[5311] = i[10];
  assign o[5312] = i[10];
  assign o[5313] = i[10];
  assign o[5314] = i[10];
  assign o[5315] = i[10];
  assign o[5316] = i[10];
  assign o[5317] = i[10];
  assign o[5318] = i[10];
  assign o[5319] = i[10];
  assign o[5320] = i[10];
  assign o[5321] = i[10];
  assign o[5322] = i[10];
  assign o[5323] = i[10];
  assign o[5324] = i[10];
  assign o[5325] = i[10];
  assign o[5326] = i[10];
  assign o[5327] = i[10];
  assign o[5328] = i[10];
  assign o[5329] = i[10];
  assign o[5330] = i[10];
  assign o[5331] = i[10];
  assign o[5332] = i[10];
  assign o[5333] = i[10];
  assign o[5334] = i[10];
  assign o[5335] = i[10];
  assign o[5336] = i[10];
  assign o[5337] = i[10];
  assign o[5338] = i[10];
  assign o[5339] = i[10];
  assign o[5340] = i[10];
  assign o[5341] = i[10];
  assign o[5342] = i[10];
  assign o[5343] = i[10];
  assign o[5344] = i[10];
  assign o[5345] = i[10];
  assign o[5346] = i[10];
  assign o[5347] = i[10];
  assign o[5348] = i[10];
  assign o[5349] = i[10];
  assign o[5350] = i[10];
  assign o[5351] = i[10];
  assign o[5352] = i[10];
  assign o[5353] = i[10];
  assign o[5354] = i[10];
  assign o[5355] = i[10];
  assign o[5356] = i[10];
  assign o[5357] = i[10];
  assign o[5358] = i[10];
  assign o[5359] = i[10];
  assign o[5360] = i[10];
  assign o[5361] = i[10];
  assign o[5362] = i[10];
  assign o[5363] = i[10];
  assign o[5364] = i[10];
  assign o[5365] = i[10];
  assign o[5366] = i[10];
  assign o[5367] = i[10];
  assign o[5368] = i[10];
  assign o[5369] = i[10];
  assign o[5370] = i[10];
  assign o[5371] = i[10];
  assign o[5372] = i[10];
  assign o[5373] = i[10];
  assign o[5374] = i[10];
  assign o[5375] = i[10];
  assign o[5376] = i[10];
  assign o[5377] = i[10];
  assign o[5378] = i[10];
  assign o[5379] = i[10];
  assign o[5380] = i[10];
  assign o[5381] = i[10];
  assign o[5382] = i[10];
  assign o[5383] = i[10];
  assign o[5384] = i[10];
  assign o[5385] = i[10];
  assign o[5386] = i[10];
  assign o[5387] = i[10];
  assign o[5388] = i[10];
  assign o[5389] = i[10];
  assign o[5390] = i[10];
  assign o[5391] = i[10];
  assign o[5392] = i[10];
  assign o[5393] = i[10];
  assign o[5394] = i[10];
  assign o[5395] = i[10];
  assign o[5396] = i[10];
  assign o[5397] = i[10];
  assign o[5398] = i[10];
  assign o[5399] = i[10];
  assign o[5400] = i[10];
  assign o[5401] = i[10];
  assign o[5402] = i[10];
  assign o[5403] = i[10];
  assign o[5404] = i[10];
  assign o[5405] = i[10];
  assign o[5406] = i[10];
  assign o[5407] = i[10];
  assign o[5408] = i[10];
  assign o[5409] = i[10];
  assign o[5410] = i[10];
  assign o[5411] = i[10];
  assign o[5412] = i[10];
  assign o[5413] = i[10];
  assign o[5414] = i[10];
  assign o[5415] = i[10];
  assign o[5416] = i[10];
  assign o[5417] = i[10];
  assign o[5418] = i[10];
  assign o[5419] = i[10];
  assign o[5420] = i[10];
  assign o[5421] = i[10];
  assign o[5422] = i[10];
  assign o[5423] = i[10];
  assign o[5424] = i[10];
  assign o[5425] = i[10];
  assign o[5426] = i[10];
  assign o[5427] = i[10];
  assign o[5428] = i[10];
  assign o[5429] = i[10];
  assign o[5430] = i[10];
  assign o[5431] = i[10];
  assign o[5432] = i[10];
  assign o[5433] = i[10];
  assign o[5434] = i[10];
  assign o[5435] = i[10];
  assign o[5436] = i[10];
  assign o[5437] = i[10];
  assign o[5438] = i[10];
  assign o[5439] = i[10];
  assign o[5440] = i[10];
  assign o[5441] = i[10];
  assign o[5442] = i[10];
  assign o[5443] = i[10];
  assign o[5444] = i[10];
  assign o[5445] = i[10];
  assign o[5446] = i[10];
  assign o[5447] = i[10];
  assign o[5448] = i[10];
  assign o[5449] = i[10];
  assign o[5450] = i[10];
  assign o[5451] = i[10];
  assign o[5452] = i[10];
  assign o[5453] = i[10];
  assign o[5454] = i[10];
  assign o[5455] = i[10];
  assign o[5456] = i[10];
  assign o[5457] = i[10];
  assign o[5458] = i[10];
  assign o[5459] = i[10];
  assign o[5460] = i[10];
  assign o[5461] = i[10];
  assign o[5462] = i[10];
  assign o[5463] = i[10];
  assign o[5464] = i[10];
  assign o[5465] = i[10];
  assign o[5466] = i[10];
  assign o[5467] = i[10];
  assign o[5468] = i[10];
  assign o[5469] = i[10];
  assign o[5470] = i[10];
  assign o[5471] = i[10];
  assign o[5472] = i[10];
  assign o[5473] = i[10];
  assign o[5474] = i[10];
  assign o[5475] = i[10];
  assign o[5476] = i[10];
  assign o[5477] = i[10];
  assign o[5478] = i[10];
  assign o[5479] = i[10];
  assign o[5480] = i[10];
  assign o[5481] = i[10];
  assign o[5482] = i[10];
  assign o[5483] = i[10];
  assign o[5484] = i[10];
  assign o[5485] = i[10];
  assign o[5486] = i[10];
  assign o[5487] = i[10];
  assign o[5488] = i[10];
  assign o[5489] = i[10];
  assign o[5490] = i[10];
  assign o[5491] = i[10];
  assign o[5492] = i[10];
  assign o[5493] = i[10];
  assign o[5494] = i[10];
  assign o[5495] = i[10];
  assign o[5496] = i[10];
  assign o[5497] = i[10];
  assign o[5498] = i[10];
  assign o[5499] = i[10];
  assign o[5500] = i[10];
  assign o[5501] = i[10];
  assign o[5502] = i[10];
  assign o[5503] = i[10];
  assign o[5504] = i[10];
  assign o[5505] = i[10];
  assign o[5506] = i[10];
  assign o[5507] = i[10];
  assign o[5508] = i[10];
  assign o[5509] = i[10];
  assign o[5510] = i[10];
  assign o[5511] = i[10];
  assign o[5512] = i[10];
  assign o[5513] = i[10];
  assign o[5514] = i[10];
  assign o[5515] = i[10];
  assign o[5516] = i[10];
  assign o[5517] = i[10];
  assign o[5518] = i[10];
  assign o[5519] = i[10];
  assign o[5520] = i[10];
  assign o[5521] = i[10];
  assign o[5522] = i[10];
  assign o[5523] = i[10];
  assign o[5524] = i[10];
  assign o[5525] = i[10];
  assign o[5526] = i[10];
  assign o[5527] = i[10];
  assign o[5528] = i[10];
  assign o[5529] = i[10];
  assign o[5530] = i[10];
  assign o[5531] = i[10];
  assign o[5532] = i[10];
  assign o[5533] = i[10];
  assign o[5534] = i[10];
  assign o[5535] = i[10];
  assign o[5536] = i[10];
  assign o[5537] = i[10];
  assign o[5538] = i[10];
  assign o[5539] = i[10];
  assign o[5540] = i[10];
  assign o[5541] = i[10];
  assign o[5542] = i[10];
  assign o[5543] = i[10];
  assign o[5544] = i[10];
  assign o[5545] = i[10];
  assign o[5546] = i[10];
  assign o[5547] = i[10];
  assign o[5548] = i[10];
  assign o[5549] = i[10];
  assign o[5550] = i[10];
  assign o[5551] = i[10];
  assign o[5552] = i[10];
  assign o[5553] = i[10];
  assign o[5554] = i[10];
  assign o[5555] = i[10];
  assign o[5556] = i[10];
  assign o[5557] = i[10];
  assign o[5558] = i[10];
  assign o[5559] = i[10];
  assign o[5560] = i[10];
  assign o[5561] = i[10];
  assign o[5562] = i[10];
  assign o[5563] = i[10];
  assign o[5564] = i[10];
  assign o[5565] = i[10];
  assign o[5566] = i[10];
  assign o[5567] = i[10];
  assign o[5568] = i[10];
  assign o[5569] = i[10];
  assign o[5570] = i[10];
  assign o[5571] = i[10];
  assign o[5572] = i[10];
  assign o[5573] = i[10];
  assign o[5574] = i[10];
  assign o[5575] = i[10];
  assign o[5576] = i[10];
  assign o[5577] = i[10];
  assign o[5578] = i[10];
  assign o[5579] = i[10];
  assign o[5580] = i[10];
  assign o[5581] = i[10];
  assign o[5582] = i[10];
  assign o[5583] = i[10];
  assign o[5584] = i[10];
  assign o[5585] = i[10];
  assign o[5586] = i[10];
  assign o[5587] = i[10];
  assign o[5588] = i[10];
  assign o[5589] = i[10];
  assign o[5590] = i[10];
  assign o[5591] = i[10];
  assign o[5592] = i[10];
  assign o[5593] = i[10];
  assign o[5594] = i[10];
  assign o[5595] = i[10];
  assign o[5596] = i[10];
  assign o[5597] = i[10];
  assign o[5598] = i[10];
  assign o[5599] = i[10];
  assign o[5600] = i[10];
  assign o[5601] = i[10];
  assign o[5602] = i[10];
  assign o[5603] = i[10];
  assign o[5604] = i[10];
  assign o[5605] = i[10];
  assign o[5606] = i[10];
  assign o[5607] = i[10];
  assign o[5608] = i[10];
  assign o[5609] = i[10];
  assign o[5610] = i[10];
  assign o[5611] = i[10];
  assign o[5612] = i[10];
  assign o[5613] = i[10];
  assign o[5614] = i[10];
  assign o[5615] = i[10];
  assign o[5616] = i[10];
  assign o[5617] = i[10];
  assign o[5618] = i[10];
  assign o[5619] = i[10];
  assign o[5620] = i[10];
  assign o[5621] = i[10];
  assign o[5622] = i[10];
  assign o[5623] = i[10];
  assign o[5624] = i[10];
  assign o[5625] = i[10];
  assign o[5626] = i[10];
  assign o[5627] = i[10];
  assign o[5628] = i[10];
  assign o[5629] = i[10];
  assign o[5630] = i[10];
  assign o[5631] = i[10];
  assign o[4608] = i[9];
  assign o[4609] = i[9];
  assign o[4610] = i[9];
  assign o[4611] = i[9];
  assign o[4612] = i[9];
  assign o[4613] = i[9];
  assign o[4614] = i[9];
  assign o[4615] = i[9];
  assign o[4616] = i[9];
  assign o[4617] = i[9];
  assign o[4618] = i[9];
  assign o[4619] = i[9];
  assign o[4620] = i[9];
  assign o[4621] = i[9];
  assign o[4622] = i[9];
  assign o[4623] = i[9];
  assign o[4624] = i[9];
  assign o[4625] = i[9];
  assign o[4626] = i[9];
  assign o[4627] = i[9];
  assign o[4628] = i[9];
  assign o[4629] = i[9];
  assign o[4630] = i[9];
  assign o[4631] = i[9];
  assign o[4632] = i[9];
  assign o[4633] = i[9];
  assign o[4634] = i[9];
  assign o[4635] = i[9];
  assign o[4636] = i[9];
  assign o[4637] = i[9];
  assign o[4638] = i[9];
  assign o[4639] = i[9];
  assign o[4640] = i[9];
  assign o[4641] = i[9];
  assign o[4642] = i[9];
  assign o[4643] = i[9];
  assign o[4644] = i[9];
  assign o[4645] = i[9];
  assign o[4646] = i[9];
  assign o[4647] = i[9];
  assign o[4648] = i[9];
  assign o[4649] = i[9];
  assign o[4650] = i[9];
  assign o[4651] = i[9];
  assign o[4652] = i[9];
  assign o[4653] = i[9];
  assign o[4654] = i[9];
  assign o[4655] = i[9];
  assign o[4656] = i[9];
  assign o[4657] = i[9];
  assign o[4658] = i[9];
  assign o[4659] = i[9];
  assign o[4660] = i[9];
  assign o[4661] = i[9];
  assign o[4662] = i[9];
  assign o[4663] = i[9];
  assign o[4664] = i[9];
  assign o[4665] = i[9];
  assign o[4666] = i[9];
  assign o[4667] = i[9];
  assign o[4668] = i[9];
  assign o[4669] = i[9];
  assign o[4670] = i[9];
  assign o[4671] = i[9];
  assign o[4672] = i[9];
  assign o[4673] = i[9];
  assign o[4674] = i[9];
  assign o[4675] = i[9];
  assign o[4676] = i[9];
  assign o[4677] = i[9];
  assign o[4678] = i[9];
  assign o[4679] = i[9];
  assign o[4680] = i[9];
  assign o[4681] = i[9];
  assign o[4682] = i[9];
  assign o[4683] = i[9];
  assign o[4684] = i[9];
  assign o[4685] = i[9];
  assign o[4686] = i[9];
  assign o[4687] = i[9];
  assign o[4688] = i[9];
  assign o[4689] = i[9];
  assign o[4690] = i[9];
  assign o[4691] = i[9];
  assign o[4692] = i[9];
  assign o[4693] = i[9];
  assign o[4694] = i[9];
  assign o[4695] = i[9];
  assign o[4696] = i[9];
  assign o[4697] = i[9];
  assign o[4698] = i[9];
  assign o[4699] = i[9];
  assign o[4700] = i[9];
  assign o[4701] = i[9];
  assign o[4702] = i[9];
  assign o[4703] = i[9];
  assign o[4704] = i[9];
  assign o[4705] = i[9];
  assign o[4706] = i[9];
  assign o[4707] = i[9];
  assign o[4708] = i[9];
  assign o[4709] = i[9];
  assign o[4710] = i[9];
  assign o[4711] = i[9];
  assign o[4712] = i[9];
  assign o[4713] = i[9];
  assign o[4714] = i[9];
  assign o[4715] = i[9];
  assign o[4716] = i[9];
  assign o[4717] = i[9];
  assign o[4718] = i[9];
  assign o[4719] = i[9];
  assign o[4720] = i[9];
  assign o[4721] = i[9];
  assign o[4722] = i[9];
  assign o[4723] = i[9];
  assign o[4724] = i[9];
  assign o[4725] = i[9];
  assign o[4726] = i[9];
  assign o[4727] = i[9];
  assign o[4728] = i[9];
  assign o[4729] = i[9];
  assign o[4730] = i[9];
  assign o[4731] = i[9];
  assign o[4732] = i[9];
  assign o[4733] = i[9];
  assign o[4734] = i[9];
  assign o[4735] = i[9];
  assign o[4736] = i[9];
  assign o[4737] = i[9];
  assign o[4738] = i[9];
  assign o[4739] = i[9];
  assign o[4740] = i[9];
  assign o[4741] = i[9];
  assign o[4742] = i[9];
  assign o[4743] = i[9];
  assign o[4744] = i[9];
  assign o[4745] = i[9];
  assign o[4746] = i[9];
  assign o[4747] = i[9];
  assign o[4748] = i[9];
  assign o[4749] = i[9];
  assign o[4750] = i[9];
  assign o[4751] = i[9];
  assign o[4752] = i[9];
  assign o[4753] = i[9];
  assign o[4754] = i[9];
  assign o[4755] = i[9];
  assign o[4756] = i[9];
  assign o[4757] = i[9];
  assign o[4758] = i[9];
  assign o[4759] = i[9];
  assign o[4760] = i[9];
  assign o[4761] = i[9];
  assign o[4762] = i[9];
  assign o[4763] = i[9];
  assign o[4764] = i[9];
  assign o[4765] = i[9];
  assign o[4766] = i[9];
  assign o[4767] = i[9];
  assign o[4768] = i[9];
  assign o[4769] = i[9];
  assign o[4770] = i[9];
  assign o[4771] = i[9];
  assign o[4772] = i[9];
  assign o[4773] = i[9];
  assign o[4774] = i[9];
  assign o[4775] = i[9];
  assign o[4776] = i[9];
  assign o[4777] = i[9];
  assign o[4778] = i[9];
  assign o[4779] = i[9];
  assign o[4780] = i[9];
  assign o[4781] = i[9];
  assign o[4782] = i[9];
  assign o[4783] = i[9];
  assign o[4784] = i[9];
  assign o[4785] = i[9];
  assign o[4786] = i[9];
  assign o[4787] = i[9];
  assign o[4788] = i[9];
  assign o[4789] = i[9];
  assign o[4790] = i[9];
  assign o[4791] = i[9];
  assign o[4792] = i[9];
  assign o[4793] = i[9];
  assign o[4794] = i[9];
  assign o[4795] = i[9];
  assign o[4796] = i[9];
  assign o[4797] = i[9];
  assign o[4798] = i[9];
  assign o[4799] = i[9];
  assign o[4800] = i[9];
  assign o[4801] = i[9];
  assign o[4802] = i[9];
  assign o[4803] = i[9];
  assign o[4804] = i[9];
  assign o[4805] = i[9];
  assign o[4806] = i[9];
  assign o[4807] = i[9];
  assign o[4808] = i[9];
  assign o[4809] = i[9];
  assign o[4810] = i[9];
  assign o[4811] = i[9];
  assign o[4812] = i[9];
  assign o[4813] = i[9];
  assign o[4814] = i[9];
  assign o[4815] = i[9];
  assign o[4816] = i[9];
  assign o[4817] = i[9];
  assign o[4818] = i[9];
  assign o[4819] = i[9];
  assign o[4820] = i[9];
  assign o[4821] = i[9];
  assign o[4822] = i[9];
  assign o[4823] = i[9];
  assign o[4824] = i[9];
  assign o[4825] = i[9];
  assign o[4826] = i[9];
  assign o[4827] = i[9];
  assign o[4828] = i[9];
  assign o[4829] = i[9];
  assign o[4830] = i[9];
  assign o[4831] = i[9];
  assign o[4832] = i[9];
  assign o[4833] = i[9];
  assign o[4834] = i[9];
  assign o[4835] = i[9];
  assign o[4836] = i[9];
  assign o[4837] = i[9];
  assign o[4838] = i[9];
  assign o[4839] = i[9];
  assign o[4840] = i[9];
  assign o[4841] = i[9];
  assign o[4842] = i[9];
  assign o[4843] = i[9];
  assign o[4844] = i[9];
  assign o[4845] = i[9];
  assign o[4846] = i[9];
  assign o[4847] = i[9];
  assign o[4848] = i[9];
  assign o[4849] = i[9];
  assign o[4850] = i[9];
  assign o[4851] = i[9];
  assign o[4852] = i[9];
  assign o[4853] = i[9];
  assign o[4854] = i[9];
  assign o[4855] = i[9];
  assign o[4856] = i[9];
  assign o[4857] = i[9];
  assign o[4858] = i[9];
  assign o[4859] = i[9];
  assign o[4860] = i[9];
  assign o[4861] = i[9];
  assign o[4862] = i[9];
  assign o[4863] = i[9];
  assign o[4864] = i[9];
  assign o[4865] = i[9];
  assign o[4866] = i[9];
  assign o[4867] = i[9];
  assign o[4868] = i[9];
  assign o[4869] = i[9];
  assign o[4870] = i[9];
  assign o[4871] = i[9];
  assign o[4872] = i[9];
  assign o[4873] = i[9];
  assign o[4874] = i[9];
  assign o[4875] = i[9];
  assign o[4876] = i[9];
  assign o[4877] = i[9];
  assign o[4878] = i[9];
  assign o[4879] = i[9];
  assign o[4880] = i[9];
  assign o[4881] = i[9];
  assign o[4882] = i[9];
  assign o[4883] = i[9];
  assign o[4884] = i[9];
  assign o[4885] = i[9];
  assign o[4886] = i[9];
  assign o[4887] = i[9];
  assign o[4888] = i[9];
  assign o[4889] = i[9];
  assign o[4890] = i[9];
  assign o[4891] = i[9];
  assign o[4892] = i[9];
  assign o[4893] = i[9];
  assign o[4894] = i[9];
  assign o[4895] = i[9];
  assign o[4896] = i[9];
  assign o[4897] = i[9];
  assign o[4898] = i[9];
  assign o[4899] = i[9];
  assign o[4900] = i[9];
  assign o[4901] = i[9];
  assign o[4902] = i[9];
  assign o[4903] = i[9];
  assign o[4904] = i[9];
  assign o[4905] = i[9];
  assign o[4906] = i[9];
  assign o[4907] = i[9];
  assign o[4908] = i[9];
  assign o[4909] = i[9];
  assign o[4910] = i[9];
  assign o[4911] = i[9];
  assign o[4912] = i[9];
  assign o[4913] = i[9];
  assign o[4914] = i[9];
  assign o[4915] = i[9];
  assign o[4916] = i[9];
  assign o[4917] = i[9];
  assign o[4918] = i[9];
  assign o[4919] = i[9];
  assign o[4920] = i[9];
  assign o[4921] = i[9];
  assign o[4922] = i[9];
  assign o[4923] = i[9];
  assign o[4924] = i[9];
  assign o[4925] = i[9];
  assign o[4926] = i[9];
  assign o[4927] = i[9];
  assign o[4928] = i[9];
  assign o[4929] = i[9];
  assign o[4930] = i[9];
  assign o[4931] = i[9];
  assign o[4932] = i[9];
  assign o[4933] = i[9];
  assign o[4934] = i[9];
  assign o[4935] = i[9];
  assign o[4936] = i[9];
  assign o[4937] = i[9];
  assign o[4938] = i[9];
  assign o[4939] = i[9];
  assign o[4940] = i[9];
  assign o[4941] = i[9];
  assign o[4942] = i[9];
  assign o[4943] = i[9];
  assign o[4944] = i[9];
  assign o[4945] = i[9];
  assign o[4946] = i[9];
  assign o[4947] = i[9];
  assign o[4948] = i[9];
  assign o[4949] = i[9];
  assign o[4950] = i[9];
  assign o[4951] = i[9];
  assign o[4952] = i[9];
  assign o[4953] = i[9];
  assign o[4954] = i[9];
  assign o[4955] = i[9];
  assign o[4956] = i[9];
  assign o[4957] = i[9];
  assign o[4958] = i[9];
  assign o[4959] = i[9];
  assign o[4960] = i[9];
  assign o[4961] = i[9];
  assign o[4962] = i[9];
  assign o[4963] = i[9];
  assign o[4964] = i[9];
  assign o[4965] = i[9];
  assign o[4966] = i[9];
  assign o[4967] = i[9];
  assign o[4968] = i[9];
  assign o[4969] = i[9];
  assign o[4970] = i[9];
  assign o[4971] = i[9];
  assign o[4972] = i[9];
  assign o[4973] = i[9];
  assign o[4974] = i[9];
  assign o[4975] = i[9];
  assign o[4976] = i[9];
  assign o[4977] = i[9];
  assign o[4978] = i[9];
  assign o[4979] = i[9];
  assign o[4980] = i[9];
  assign o[4981] = i[9];
  assign o[4982] = i[9];
  assign o[4983] = i[9];
  assign o[4984] = i[9];
  assign o[4985] = i[9];
  assign o[4986] = i[9];
  assign o[4987] = i[9];
  assign o[4988] = i[9];
  assign o[4989] = i[9];
  assign o[4990] = i[9];
  assign o[4991] = i[9];
  assign o[4992] = i[9];
  assign o[4993] = i[9];
  assign o[4994] = i[9];
  assign o[4995] = i[9];
  assign o[4996] = i[9];
  assign o[4997] = i[9];
  assign o[4998] = i[9];
  assign o[4999] = i[9];
  assign o[5000] = i[9];
  assign o[5001] = i[9];
  assign o[5002] = i[9];
  assign o[5003] = i[9];
  assign o[5004] = i[9];
  assign o[5005] = i[9];
  assign o[5006] = i[9];
  assign o[5007] = i[9];
  assign o[5008] = i[9];
  assign o[5009] = i[9];
  assign o[5010] = i[9];
  assign o[5011] = i[9];
  assign o[5012] = i[9];
  assign o[5013] = i[9];
  assign o[5014] = i[9];
  assign o[5015] = i[9];
  assign o[5016] = i[9];
  assign o[5017] = i[9];
  assign o[5018] = i[9];
  assign o[5019] = i[9];
  assign o[5020] = i[9];
  assign o[5021] = i[9];
  assign o[5022] = i[9];
  assign o[5023] = i[9];
  assign o[5024] = i[9];
  assign o[5025] = i[9];
  assign o[5026] = i[9];
  assign o[5027] = i[9];
  assign o[5028] = i[9];
  assign o[5029] = i[9];
  assign o[5030] = i[9];
  assign o[5031] = i[9];
  assign o[5032] = i[9];
  assign o[5033] = i[9];
  assign o[5034] = i[9];
  assign o[5035] = i[9];
  assign o[5036] = i[9];
  assign o[5037] = i[9];
  assign o[5038] = i[9];
  assign o[5039] = i[9];
  assign o[5040] = i[9];
  assign o[5041] = i[9];
  assign o[5042] = i[9];
  assign o[5043] = i[9];
  assign o[5044] = i[9];
  assign o[5045] = i[9];
  assign o[5046] = i[9];
  assign o[5047] = i[9];
  assign o[5048] = i[9];
  assign o[5049] = i[9];
  assign o[5050] = i[9];
  assign o[5051] = i[9];
  assign o[5052] = i[9];
  assign o[5053] = i[9];
  assign o[5054] = i[9];
  assign o[5055] = i[9];
  assign o[5056] = i[9];
  assign o[5057] = i[9];
  assign o[5058] = i[9];
  assign o[5059] = i[9];
  assign o[5060] = i[9];
  assign o[5061] = i[9];
  assign o[5062] = i[9];
  assign o[5063] = i[9];
  assign o[5064] = i[9];
  assign o[5065] = i[9];
  assign o[5066] = i[9];
  assign o[5067] = i[9];
  assign o[5068] = i[9];
  assign o[5069] = i[9];
  assign o[5070] = i[9];
  assign o[5071] = i[9];
  assign o[5072] = i[9];
  assign o[5073] = i[9];
  assign o[5074] = i[9];
  assign o[5075] = i[9];
  assign o[5076] = i[9];
  assign o[5077] = i[9];
  assign o[5078] = i[9];
  assign o[5079] = i[9];
  assign o[5080] = i[9];
  assign o[5081] = i[9];
  assign o[5082] = i[9];
  assign o[5083] = i[9];
  assign o[5084] = i[9];
  assign o[5085] = i[9];
  assign o[5086] = i[9];
  assign o[5087] = i[9];
  assign o[5088] = i[9];
  assign o[5089] = i[9];
  assign o[5090] = i[9];
  assign o[5091] = i[9];
  assign o[5092] = i[9];
  assign o[5093] = i[9];
  assign o[5094] = i[9];
  assign o[5095] = i[9];
  assign o[5096] = i[9];
  assign o[5097] = i[9];
  assign o[5098] = i[9];
  assign o[5099] = i[9];
  assign o[5100] = i[9];
  assign o[5101] = i[9];
  assign o[5102] = i[9];
  assign o[5103] = i[9];
  assign o[5104] = i[9];
  assign o[5105] = i[9];
  assign o[5106] = i[9];
  assign o[5107] = i[9];
  assign o[5108] = i[9];
  assign o[5109] = i[9];
  assign o[5110] = i[9];
  assign o[5111] = i[9];
  assign o[5112] = i[9];
  assign o[5113] = i[9];
  assign o[5114] = i[9];
  assign o[5115] = i[9];
  assign o[5116] = i[9];
  assign o[5117] = i[9];
  assign o[5118] = i[9];
  assign o[5119] = i[9];
  assign o[4096] = i[8];
  assign o[4097] = i[8];
  assign o[4098] = i[8];
  assign o[4099] = i[8];
  assign o[4100] = i[8];
  assign o[4101] = i[8];
  assign o[4102] = i[8];
  assign o[4103] = i[8];
  assign o[4104] = i[8];
  assign o[4105] = i[8];
  assign o[4106] = i[8];
  assign o[4107] = i[8];
  assign o[4108] = i[8];
  assign o[4109] = i[8];
  assign o[4110] = i[8];
  assign o[4111] = i[8];
  assign o[4112] = i[8];
  assign o[4113] = i[8];
  assign o[4114] = i[8];
  assign o[4115] = i[8];
  assign o[4116] = i[8];
  assign o[4117] = i[8];
  assign o[4118] = i[8];
  assign o[4119] = i[8];
  assign o[4120] = i[8];
  assign o[4121] = i[8];
  assign o[4122] = i[8];
  assign o[4123] = i[8];
  assign o[4124] = i[8];
  assign o[4125] = i[8];
  assign o[4126] = i[8];
  assign o[4127] = i[8];
  assign o[4128] = i[8];
  assign o[4129] = i[8];
  assign o[4130] = i[8];
  assign o[4131] = i[8];
  assign o[4132] = i[8];
  assign o[4133] = i[8];
  assign o[4134] = i[8];
  assign o[4135] = i[8];
  assign o[4136] = i[8];
  assign o[4137] = i[8];
  assign o[4138] = i[8];
  assign o[4139] = i[8];
  assign o[4140] = i[8];
  assign o[4141] = i[8];
  assign o[4142] = i[8];
  assign o[4143] = i[8];
  assign o[4144] = i[8];
  assign o[4145] = i[8];
  assign o[4146] = i[8];
  assign o[4147] = i[8];
  assign o[4148] = i[8];
  assign o[4149] = i[8];
  assign o[4150] = i[8];
  assign o[4151] = i[8];
  assign o[4152] = i[8];
  assign o[4153] = i[8];
  assign o[4154] = i[8];
  assign o[4155] = i[8];
  assign o[4156] = i[8];
  assign o[4157] = i[8];
  assign o[4158] = i[8];
  assign o[4159] = i[8];
  assign o[4160] = i[8];
  assign o[4161] = i[8];
  assign o[4162] = i[8];
  assign o[4163] = i[8];
  assign o[4164] = i[8];
  assign o[4165] = i[8];
  assign o[4166] = i[8];
  assign o[4167] = i[8];
  assign o[4168] = i[8];
  assign o[4169] = i[8];
  assign o[4170] = i[8];
  assign o[4171] = i[8];
  assign o[4172] = i[8];
  assign o[4173] = i[8];
  assign o[4174] = i[8];
  assign o[4175] = i[8];
  assign o[4176] = i[8];
  assign o[4177] = i[8];
  assign o[4178] = i[8];
  assign o[4179] = i[8];
  assign o[4180] = i[8];
  assign o[4181] = i[8];
  assign o[4182] = i[8];
  assign o[4183] = i[8];
  assign o[4184] = i[8];
  assign o[4185] = i[8];
  assign o[4186] = i[8];
  assign o[4187] = i[8];
  assign o[4188] = i[8];
  assign o[4189] = i[8];
  assign o[4190] = i[8];
  assign o[4191] = i[8];
  assign o[4192] = i[8];
  assign o[4193] = i[8];
  assign o[4194] = i[8];
  assign o[4195] = i[8];
  assign o[4196] = i[8];
  assign o[4197] = i[8];
  assign o[4198] = i[8];
  assign o[4199] = i[8];
  assign o[4200] = i[8];
  assign o[4201] = i[8];
  assign o[4202] = i[8];
  assign o[4203] = i[8];
  assign o[4204] = i[8];
  assign o[4205] = i[8];
  assign o[4206] = i[8];
  assign o[4207] = i[8];
  assign o[4208] = i[8];
  assign o[4209] = i[8];
  assign o[4210] = i[8];
  assign o[4211] = i[8];
  assign o[4212] = i[8];
  assign o[4213] = i[8];
  assign o[4214] = i[8];
  assign o[4215] = i[8];
  assign o[4216] = i[8];
  assign o[4217] = i[8];
  assign o[4218] = i[8];
  assign o[4219] = i[8];
  assign o[4220] = i[8];
  assign o[4221] = i[8];
  assign o[4222] = i[8];
  assign o[4223] = i[8];
  assign o[4224] = i[8];
  assign o[4225] = i[8];
  assign o[4226] = i[8];
  assign o[4227] = i[8];
  assign o[4228] = i[8];
  assign o[4229] = i[8];
  assign o[4230] = i[8];
  assign o[4231] = i[8];
  assign o[4232] = i[8];
  assign o[4233] = i[8];
  assign o[4234] = i[8];
  assign o[4235] = i[8];
  assign o[4236] = i[8];
  assign o[4237] = i[8];
  assign o[4238] = i[8];
  assign o[4239] = i[8];
  assign o[4240] = i[8];
  assign o[4241] = i[8];
  assign o[4242] = i[8];
  assign o[4243] = i[8];
  assign o[4244] = i[8];
  assign o[4245] = i[8];
  assign o[4246] = i[8];
  assign o[4247] = i[8];
  assign o[4248] = i[8];
  assign o[4249] = i[8];
  assign o[4250] = i[8];
  assign o[4251] = i[8];
  assign o[4252] = i[8];
  assign o[4253] = i[8];
  assign o[4254] = i[8];
  assign o[4255] = i[8];
  assign o[4256] = i[8];
  assign o[4257] = i[8];
  assign o[4258] = i[8];
  assign o[4259] = i[8];
  assign o[4260] = i[8];
  assign o[4261] = i[8];
  assign o[4262] = i[8];
  assign o[4263] = i[8];
  assign o[4264] = i[8];
  assign o[4265] = i[8];
  assign o[4266] = i[8];
  assign o[4267] = i[8];
  assign o[4268] = i[8];
  assign o[4269] = i[8];
  assign o[4270] = i[8];
  assign o[4271] = i[8];
  assign o[4272] = i[8];
  assign o[4273] = i[8];
  assign o[4274] = i[8];
  assign o[4275] = i[8];
  assign o[4276] = i[8];
  assign o[4277] = i[8];
  assign o[4278] = i[8];
  assign o[4279] = i[8];
  assign o[4280] = i[8];
  assign o[4281] = i[8];
  assign o[4282] = i[8];
  assign o[4283] = i[8];
  assign o[4284] = i[8];
  assign o[4285] = i[8];
  assign o[4286] = i[8];
  assign o[4287] = i[8];
  assign o[4288] = i[8];
  assign o[4289] = i[8];
  assign o[4290] = i[8];
  assign o[4291] = i[8];
  assign o[4292] = i[8];
  assign o[4293] = i[8];
  assign o[4294] = i[8];
  assign o[4295] = i[8];
  assign o[4296] = i[8];
  assign o[4297] = i[8];
  assign o[4298] = i[8];
  assign o[4299] = i[8];
  assign o[4300] = i[8];
  assign o[4301] = i[8];
  assign o[4302] = i[8];
  assign o[4303] = i[8];
  assign o[4304] = i[8];
  assign o[4305] = i[8];
  assign o[4306] = i[8];
  assign o[4307] = i[8];
  assign o[4308] = i[8];
  assign o[4309] = i[8];
  assign o[4310] = i[8];
  assign o[4311] = i[8];
  assign o[4312] = i[8];
  assign o[4313] = i[8];
  assign o[4314] = i[8];
  assign o[4315] = i[8];
  assign o[4316] = i[8];
  assign o[4317] = i[8];
  assign o[4318] = i[8];
  assign o[4319] = i[8];
  assign o[4320] = i[8];
  assign o[4321] = i[8];
  assign o[4322] = i[8];
  assign o[4323] = i[8];
  assign o[4324] = i[8];
  assign o[4325] = i[8];
  assign o[4326] = i[8];
  assign o[4327] = i[8];
  assign o[4328] = i[8];
  assign o[4329] = i[8];
  assign o[4330] = i[8];
  assign o[4331] = i[8];
  assign o[4332] = i[8];
  assign o[4333] = i[8];
  assign o[4334] = i[8];
  assign o[4335] = i[8];
  assign o[4336] = i[8];
  assign o[4337] = i[8];
  assign o[4338] = i[8];
  assign o[4339] = i[8];
  assign o[4340] = i[8];
  assign o[4341] = i[8];
  assign o[4342] = i[8];
  assign o[4343] = i[8];
  assign o[4344] = i[8];
  assign o[4345] = i[8];
  assign o[4346] = i[8];
  assign o[4347] = i[8];
  assign o[4348] = i[8];
  assign o[4349] = i[8];
  assign o[4350] = i[8];
  assign o[4351] = i[8];
  assign o[4352] = i[8];
  assign o[4353] = i[8];
  assign o[4354] = i[8];
  assign o[4355] = i[8];
  assign o[4356] = i[8];
  assign o[4357] = i[8];
  assign o[4358] = i[8];
  assign o[4359] = i[8];
  assign o[4360] = i[8];
  assign o[4361] = i[8];
  assign o[4362] = i[8];
  assign o[4363] = i[8];
  assign o[4364] = i[8];
  assign o[4365] = i[8];
  assign o[4366] = i[8];
  assign o[4367] = i[8];
  assign o[4368] = i[8];
  assign o[4369] = i[8];
  assign o[4370] = i[8];
  assign o[4371] = i[8];
  assign o[4372] = i[8];
  assign o[4373] = i[8];
  assign o[4374] = i[8];
  assign o[4375] = i[8];
  assign o[4376] = i[8];
  assign o[4377] = i[8];
  assign o[4378] = i[8];
  assign o[4379] = i[8];
  assign o[4380] = i[8];
  assign o[4381] = i[8];
  assign o[4382] = i[8];
  assign o[4383] = i[8];
  assign o[4384] = i[8];
  assign o[4385] = i[8];
  assign o[4386] = i[8];
  assign o[4387] = i[8];
  assign o[4388] = i[8];
  assign o[4389] = i[8];
  assign o[4390] = i[8];
  assign o[4391] = i[8];
  assign o[4392] = i[8];
  assign o[4393] = i[8];
  assign o[4394] = i[8];
  assign o[4395] = i[8];
  assign o[4396] = i[8];
  assign o[4397] = i[8];
  assign o[4398] = i[8];
  assign o[4399] = i[8];
  assign o[4400] = i[8];
  assign o[4401] = i[8];
  assign o[4402] = i[8];
  assign o[4403] = i[8];
  assign o[4404] = i[8];
  assign o[4405] = i[8];
  assign o[4406] = i[8];
  assign o[4407] = i[8];
  assign o[4408] = i[8];
  assign o[4409] = i[8];
  assign o[4410] = i[8];
  assign o[4411] = i[8];
  assign o[4412] = i[8];
  assign o[4413] = i[8];
  assign o[4414] = i[8];
  assign o[4415] = i[8];
  assign o[4416] = i[8];
  assign o[4417] = i[8];
  assign o[4418] = i[8];
  assign o[4419] = i[8];
  assign o[4420] = i[8];
  assign o[4421] = i[8];
  assign o[4422] = i[8];
  assign o[4423] = i[8];
  assign o[4424] = i[8];
  assign o[4425] = i[8];
  assign o[4426] = i[8];
  assign o[4427] = i[8];
  assign o[4428] = i[8];
  assign o[4429] = i[8];
  assign o[4430] = i[8];
  assign o[4431] = i[8];
  assign o[4432] = i[8];
  assign o[4433] = i[8];
  assign o[4434] = i[8];
  assign o[4435] = i[8];
  assign o[4436] = i[8];
  assign o[4437] = i[8];
  assign o[4438] = i[8];
  assign o[4439] = i[8];
  assign o[4440] = i[8];
  assign o[4441] = i[8];
  assign o[4442] = i[8];
  assign o[4443] = i[8];
  assign o[4444] = i[8];
  assign o[4445] = i[8];
  assign o[4446] = i[8];
  assign o[4447] = i[8];
  assign o[4448] = i[8];
  assign o[4449] = i[8];
  assign o[4450] = i[8];
  assign o[4451] = i[8];
  assign o[4452] = i[8];
  assign o[4453] = i[8];
  assign o[4454] = i[8];
  assign o[4455] = i[8];
  assign o[4456] = i[8];
  assign o[4457] = i[8];
  assign o[4458] = i[8];
  assign o[4459] = i[8];
  assign o[4460] = i[8];
  assign o[4461] = i[8];
  assign o[4462] = i[8];
  assign o[4463] = i[8];
  assign o[4464] = i[8];
  assign o[4465] = i[8];
  assign o[4466] = i[8];
  assign o[4467] = i[8];
  assign o[4468] = i[8];
  assign o[4469] = i[8];
  assign o[4470] = i[8];
  assign o[4471] = i[8];
  assign o[4472] = i[8];
  assign o[4473] = i[8];
  assign o[4474] = i[8];
  assign o[4475] = i[8];
  assign o[4476] = i[8];
  assign o[4477] = i[8];
  assign o[4478] = i[8];
  assign o[4479] = i[8];
  assign o[4480] = i[8];
  assign o[4481] = i[8];
  assign o[4482] = i[8];
  assign o[4483] = i[8];
  assign o[4484] = i[8];
  assign o[4485] = i[8];
  assign o[4486] = i[8];
  assign o[4487] = i[8];
  assign o[4488] = i[8];
  assign o[4489] = i[8];
  assign o[4490] = i[8];
  assign o[4491] = i[8];
  assign o[4492] = i[8];
  assign o[4493] = i[8];
  assign o[4494] = i[8];
  assign o[4495] = i[8];
  assign o[4496] = i[8];
  assign o[4497] = i[8];
  assign o[4498] = i[8];
  assign o[4499] = i[8];
  assign o[4500] = i[8];
  assign o[4501] = i[8];
  assign o[4502] = i[8];
  assign o[4503] = i[8];
  assign o[4504] = i[8];
  assign o[4505] = i[8];
  assign o[4506] = i[8];
  assign o[4507] = i[8];
  assign o[4508] = i[8];
  assign o[4509] = i[8];
  assign o[4510] = i[8];
  assign o[4511] = i[8];
  assign o[4512] = i[8];
  assign o[4513] = i[8];
  assign o[4514] = i[8];
  assign o[4515] = i[8];
  assign o[4516] = i[8];
  assign o[4517] = i[8];
  assign o[4518] = i[8];
  assign o[4519] = i[8];
  assign o[4520] = i[8];
  assign o[4521] = i[8];
  assign o[4522] = i[8];
  assign o[4523] = i[8];
  assign o[4524] = i[8];
  assign o[4525] = i[8];
  assign o[4526] = i[8];
  assign o[4527] = i[8];
  assign o[4528] = i[8];
  assign o[4529] = i[8];
  assign o[4530] = i[8];
  assign o[4531] = i[8];
  assign o[4532] = i[8];
  assign o[4533] = i[8];
  assign o[4534] = i[8];
  assign o[4535] = i[8];
  assign o[4536] = i[8];
  assign o[4537] = i[8];
  assign o[4538] = i[8];
  assign o[4539] = i[8];
  assign o[4540] = i[8];
  assign o[4541] = i[8];
  assign o[4542] = i[8];
  assign o[4543] = i[8];
  assign o[4544] = i[8];
  assign o[4545] = i[8];
  assign o[4546] = i[8];
  assign o[4547] = i[8];
  assign o[4548] = i[8];
  assign o[4549] = i[8];
  assign o[4550] = i[8];
  assign o[4551] = i[8];
  assign o[4552] = i[8];
  assign o[4553] = i[8];
  assign o[4554] = i[8];
  assign o[4555] = i[8];
  assign o[4556] = i[8];
  assign o[4557] = i[8];
  assign o[4558] = i[8];
  assign o[4559] = i[8];
  assign o[4560] = i[8];
  assign o[4561] = i[8];
  assign o[4562] = i[8];
  assign o[4563] = i[8];
  assign o[4564] = i[8];
  assign o[4565] = i[8];
  assign o[4566] = i[8];
  assign o[4567] = i[8];
  assign o[4568] = i[8];
  assign o[4569] = i[8];
  assign o[4570] = i[8];
  assign o[4571] = i[8];
  assign o[4572] = i[8];
  assign o[4573] = i[8];
  assign o[4574] = i[8];
  assign o[4575] = i[8];
  assign o[4576] = i[8];
  assign o[4577] = i[8];
  assign o[4578] = i[8];
  assign o[4579] = i[8];
  assign o[4580] = i[8];
  assign o[4581] = i[8];
  assign o[4582] = i[8];
  assign o[4583] = i[8];
  assign o[4584] = i[8];
  assign o[4585] = i[8];
  assign o[4586] = i[8];
  assign o[4587] = i[8];
  assign o[4588] = i[8];
  assign o[4589] = i[8];
  assign o[4590] = i[8];
  assign o[4591] = i[8];
  assign o[4592] = i[8];
  assign o[4593] = i[8];
  assign o[4594] = i[8];
  assign o[4595] = i[8];
  assign o[4596] = i[8];
  assign o[4597] = i[8];
  assign o[4598] = i[8];
  assign o[4599] = i[8];
  assign o[4600] = i[8];
  assign o[4601] = i[8];
  assign o[4602] = i[8];
  assign o[4603] = i[8];
  assign o[4604] = i[8];
  assign o[4605] = i[8];
  assign o[4606] = i[8];
  assign o[4607] = i[8];
  assign o[3584] = i[7];
  assign o[3585] = i[7];
  assign o[3586] = i[7];
  assign o[3587] = i[7];
  assign o[3588] = i[7];
  assign o[3589] = i[7];
  assign o[3590] = i[7];
  assign o[3591] = i[7];
  assign o[3592] = i[7];
  assign o[3593] = i[7];
  assign o[3594] = i[7];
  assign o[3595] = i[7];
  assign o[3596] = i[7];
  assign o[3597] = i[7];
  assign o[3598] = i[7];
  assign o[3599] = i[7];
  assign o[3600] = i[7];
  assign o[3601] = i[7];
  assign o[3602] = i[7];
  assign o[3603] = i[7];
  assign o[3604] = i[7];
  assign o[3605] = i[7];
  assign o[3606] = i[7];
  assign o[3607] = i[7];
  assign o[3608] = i[7];
  assign o[3609] = i[7];
  assign o[3610] = i[7];
  assign o[3611] = i[7];
  assign o[3612] = i[7];
  assign o[3613] = i[7];
  assign o[3614] = i[7];
  assign o[3615] = i[7];
  assign o[3616] = i[7];
  assign o[3617] = i[7];
  assign o[3618] = i[7];
  assign o[3619] = i[7];
  assign o[3620] = i[7];
  assign o[3621] = i[7];
  assign o[3622] = i[7];
  assign o[3623] = i[7];
  assign o[3624] = i[7];
  assign o[3625] = i[7];
  assign o[3626] = i[7];
  assign o[3627] = i[7];
  assign o[3628] = i[7];
  assign o[3629] = i[7];
  assign o[3630] = i[7];
  assign o[3631] = i[7];
  assign o[3632] = i[7];
  assign o[3633] = i[7];
  assign o[3634] = i[7];
  assign o[3635] = i[7];
  assign o[3636] = i[7];
  assign o[3637] = i[7];
  assign o[3638] = i[7];
  assign o[3639] = i[7];
  assign o[3640] = i[7];
  assign o[3641] = i[7];
  assign o[3642] = i[7];
  assign o[3643] = i[7];
  assign o[3644] = i[7];
  assign o[3645] = i[7];
  assign o[3646] = i[7];
  assign o[3647] = i[7];
  assign o[3648] = i[7];
  assign o[3649] = i[7];
  assign o[3650] = i[7];
  assign o[3651] = i[7];
  assign o[3652] = i[7];
  assign o[3653] = i[7];
  assign o[3654] = i[7];
  assign o[3655] = i[7];
  assign o[3656] = i[7];
  assign o[3657] = i[7];
  assign o[3658] = i[7];
  assign o[3659] = i[7];
  assign o[3660] = i[7];
  assign o[3661] = i[7];
  assign o[3662] = i[7];
  assign o[3663] = i[7];
  assign o[3664] = i[7];
  assign o[3665] = i[7];
  assign o[3666] = i[7];
  assign o[3667] = i[7];
  assign o[3668] = i[7];
  assign o[3669] = i[7];
  assign o[3670] = i[7];
  assign o[3671] = i[7];
  assign o[3672] = i[7];
  assign o[3673] = i[7];
  assign o[3674] = i[7];
  assign o[3675] = i[7];
  assign o[3676] = i[7];
  assign o[3677] = i[7];
  assign o[3678] = i[7];
  assign o[3679] = i[7];
  assign o[3680] = i[7];
  assign o[3681] = i[7];
  assign o[3682] = i[7];
  assign o[3683] = i[7];
  assign o[3684] = i[7];
  assign o[3685] = i[7];
  assign o[3686] = i[7];
  assign o[3687] = i[7];
  assign o[3688] = i[7];
  assign o[3689] = i[7];
  assign o[3690] = i[7];
  assign o[3691] = i[7];
  assign o[3692] = i[7];
  assign o[3693] = i[7];
  assign o[3694] = i[7];
  assign o[3695] = i[7];
  assign o[3696] = i[7];
  assign o[3697] = i[7];
  assign o[3698] = i[7];
  assign o[3699] = i[7];
  assign o[3700] = i[7];
  assign o[3701] = i[7];
  assign o[3702] = i[7];
  assign o[3703] = i[7];
  assign o[3704] = i[7];
  assign o[3705] = i[7];
  assign o[3706] = i[7];
  assign o[3707] = i[7];
  assign o[3708] = i[7];
  assign o[3709] = i[7];
  assign o[3710] = i[7];
  assign o[3711] = i[7];
  assign o[3712] = i[7];
  assign o[3713] = i[7];
  assign o[3714] = i[7];
  assign o[3715] = i[7];
  assign o[3716] = i[7];
  assign o[3717] = i[7];
  assign o[3718] = i[7];
  assign o[3719] = i[7];
  assign o[3720] = i[7];
  assign o[3721] = i[7];
  assign o[3722] = i[7];
  assign o[3723] = i[7];
  assign o[3724] = i[7];
  assign o[3725] = i[7];
  assign o[3726] = i[7];
  assign o[3727] = i[7];
  assign o[3728] = i[7];
  assign o[3729] = i[7];
  assign o[3730] = i[7];
  assign o[3731] = i[7];
  assign o[3732] = i[7];
  assign o[3733] = i[7];
  assign o[3734] = i[7];
  assign o[3735] = i[7];
  assign o[3736] = i[7];
  assign o[3737] = i[7];
  assign o[3738] = i[7];
  assign o[3739] = i[7];
  assign o[3740] = i[7];
  assign o[3741] = i[7];
  assign o[3742] = i[7];
  assign o[3743] = i[7];
  assign o[3744] = i[7];
  assign o[3745] = i[7];
  assign o[3746] = i[7];
  assign o[3747] = i[7];
  assign o[3748] = i[7];
  assign o[3749] = i[7];
  assign o[3750] = i[7];
  assign o[3751] = i[7];
  assign o[3752] = i[7];
  assign o[3753] = i[7];
  assign o[3754] = i[7];
  assign o[3755] = i[7];
  assign o[3756] = i[7];
  assign o[3757] = i[7];
  assign o[3758] = i[7];
  assign o[3759] = i[7];
  assign o[3760] = i[7];
  assign o[3761] = i[7];
  assign o[3762] = i[7];
  assign o[3763] = i[7];
  assign o[3764] = i[7];
  assign o[3765] = i[7];
  assign o[3766] = i[7];
  assign o[3767] = i[7];
  assign o[3768] = i[7];
  assign o[3769] = i[7];
  assign o[3770] = i[7];
  assign o[3771] = i[7];
  assign o[3772] = i[7];
  assign o[3773] = i[7];
  assign o[3774] = i[7];
  assign o[3775] = i[7];
  assign o[3776] = i[7];
  assign o[3777] = i[7];
  assign o[3778] = i[7];
  assign o[3779] = i[7];
  assign o[3780] = i[7];
  assign o[3781] = i[7];
  assign o[3782] = i[7];
  assign o[3783] = i[7];
  assign o[3784] = i[7];
  assign o[3785] = i[7];
  assign o[3786] = i[7];
  assign o[3787] = i[7];
  assign o[3788] = i[7];
  assign o[3789] = i[7];
  assign o[3790] = i[7];
  assign o[3791] = i[7];
  assign o[3792] = i[7];
  assign o[3793] = i[7];
  assign o[3794] = i[7];
  assign o[3795] = i[7];
  assign o[3796] = i[7];
  assign o[3797] = i[7];
  assign o[3798] = i[7];
  assign o[3799] = i[7];
  assign o[3800] = i[7];
  assign o[3801] = i[7];
  assign o[3802] = i[7];
  assign o[3803] = i[7];
  assign o[3804] = i[7];
  assign o[3805] = i[7];
  assign o[3806] = i[7];
  assign o[3807] = i[7];
  assign o[3808] = i[7];
  assign o[3809] = i[7];
  assign o[3810] = i[7];
  assign o[3811] = i[7];
  assign o[3812] = i[7];
  assign o[3813] = i[7];
  assign o[3814] = i[7];
  assign o[3815] = i[7];
  assign o[3816] = i[7];
  assign o[3817] = i[7];
  assign o[3818] = i[7];
  assign o[3819] = i[7];
  assign o[3820] = i[7];
  assign o[3821] = i[7];
  assign o[3822] = i[7];
  assign o[3823] = i[7];
  assign o[3824] = i[7];
  assign o[3825] = i[7];
  assign o[3826] = i[7];
  assign o[3827] = i[7];
  assign o[3828] = i[7];
  assign o[3829] = i[7];
  assign o[3830] = i[7];
  assign o[3831] = i[7];
  assign o[3832] = i[7];
  assign o[3833] = i[7];
  assign o[3834] = i[7];
  assign o[3835] = i[7];
  assign o[3836] = i[7];
  assign o[3837] = i[7];
  assign o[3838] = i[7];
  assign o[3839] = i[7];
  assign o[3840] = i[7];
  assign o[3841] = i[7];
  assign o[3842] = i[7];
  assign o[3843] = i[7];
  assign o[3844] = i[7];
  assign o[3845] = i[7];
  assign o[3846] = i[7];
  assign o[3847] = i[7];
  assign o[3848] = i[7];
  assign o[3849] = i[7];
  assign o[3850] = i[7];
  assign o[3851] = i[7];
  assign o[3852] = i[7];
  assign o[3853] = i[7];
  assign o[3854] = i[7];
  assign o[3855] = i[7];
  assign o[3856] = i[7];
  assign o[3857] = i[7];
  assign o[3858] = i[7];
  assign o[3859] = i[7];
  assign o[3860] = i[7];
  assign o[3861] = i[7];
  assign o[3862] = i[7];
  assign o[3863] = i[7];
  assign o[3864] = i[7];
  assign o[3865] = i[7];
  assign o[3866] = i[7];
  assign o[3867] = i[7];
  assign o[3868] = i[7];
  assign o[3869] = i[7];
  assign o[3870] = i[7];
  assign o[3871] = i[7];
  assign o[3872] = i[7];
  assign o[3873] = i[7];
  assign o[3874] = i[7];
  assign o[3875] = i[7];
  assign o[3876] = i[7];
  assign o[3877] = i[7];
  assign o[3878] = i[7];
  assign o[3879] = i[7];
  assign o[3880] = i[7];
  assign o[3881] = i[7];
  assign o[3882] = i[7];
  assign o[3883] = i[7];
  assign o[3884] = i[7];
  assign o[3885] = i[7];
  assign o[3886] = i[7];
  assign o[3887] = i[7];
  assign o[3888] = i[7];
  assign o[3889] = i[7];
  assign o[3890] = i[7];
  assign o[3891] = i[7];
  assign o[3892] = i[7];
  assign o[3893] = i[7];
  assign o[3894] = i[7];
  assign o[3895] = i[7];
  assign o[3896] = i[7];
  assign o[3897] = i[7];
  assign o[3898] = i[7];
  assign o[3899] = i[7];
  assign o[3900] = i[7];
  assign o[3901] = i[7];
  assign o[3902] = i[7];
  assign o[3903] = i[7];
  assign o[3904] = i[7];
  assign o[3905] = i[7];
  assign o[3906] = i[7];
  assign o[3907] = i[7];
  assign o[3908] = i[7];
  assign o[3909] = i[7];
  assign o[3910] = i[7];
  assign o[3911] = i[7];
  assign o[3912] = i[7];
  assign o[3913] = i[7];
  assign o[3914] = i[7];
  assign o[3915] = i[7];
  assign o[3916] = i[7];
  assign o[3917] = i[7];
  assign o[3918] = i[7];
  assign o[3919] = i[7];
  assign o[3920] = i[7];
  assign o[3921] = i[7];
  assign o[3922] = i[7];
  assign o[3923] = i[7];
  assign o[3924] = i[7];
  assign o[3925] = i[7];
  assign o[3926] = i[7];
  assign o[3927] = i[7];
  assign o[3928] = i[7];
  assign o[3929] = i[7];
  assign o[3930] = i[7];
  assign o[3931] = i[7];
  assign o[3932] = i[7];
  assign o[3933] = i[7];
  assign o[3934] = i[7];
  assign o[3935] = i[7];
  assign o[3936] = i[7];
  assign o[3937] = i[7];
  assign o[3938] = i[7];
  assign o[3939] = i[7];
  assign o[3940] = i[7];
  assign o[3941] = i[7];
  assign o[3942] = i[7];
  assign o[3943] = i[7];
  assign o[3944] = i[7];
  assign o[3945] = i[7];
  assign o[3946] = i[7];
  assign o[3947] = i[7];
  assign o[3948] = i[7];
  assign o[3949] = i[7];
  assign o[3950] = i[7];
  assign o[3951] = i[7];
  assign o[3952] = i[7];
  assign o[3953] = i[7];
  assign o[3954] = i[7];
  assign o[3955] = i[7];
  assign o[3956] = i[7];
  assign o[3957] = i[7];
  assign o[3958] = i[7];
  assign o[3959] = i[7];
  assign o[3960] = i[7];
  assign o[3961] = i[7];
  assign o[3962] = i[7];
  assign o[3963] = i[7];
  assign o[3964] = i[7];
  assign o[3965] = i[7];
  assign o[3966] = i[7];
  assign o[3967] = i[7];
  assign o[3968] = i[7];
  assign o[3969] = i[7];
  assign o[3970] = i[7];
  assign o[3971] = i[7];
  assign o[3972] = i[7];
  assign o[3973] = i[7];
  assign o[3974] = i[7];
  assign o[3975] = i[7];
  assign o[3976] = i[7];
  assign o[3977] = i[7];
  assign o[3978] = i[7];
  assign o[3979] = i[7];
  assign o[3980] = i[7];
  assign o[3981] = i[7];
  assign o[3982] = i[7];
  assign o[3983] = i[7];
  assign o[3984] = i[7];
  assign o[3985] = i[7];
  assign o[3986] = i[7];
  assign o[3987] = i[7];
  assign o[3988] = i[7];
  assign o[3989] = i[7];
  assign o[3990] = i[7];
  assign o[3991] = i[7];
  assign o[3992] = i[7];
  assign o[3993] = i[7];
  assign o[3994] = i[7];
  assign o[3995] = i[7];
  assign o[3996] = i[7];
  assign o[3997] = i[7];
  assign o[3998] = i[7];
  assign o[3999] = i[7];
  assign o[4000] = i[7];
  assign o[4001] = i[7];
  assign o[4002] = i[7];
  assign o[4003] = i[7];
  assign o[4004] = i[7];
  assign o[4005] = i[7];
  assign o[4006] = i[7];
  assign o[4007] = i[7];
  assign o[4008] = i[7];
  assign o[4009] = i[7];
  assign o[4010] = i[7];
  assign o[4011] = i[7];
  assign o[4012] = i[7];
  assign o[4013] = i[7];
  assign o[4014] = i[7];
  assign o[4015] = i[7];
  assign o[4016] = i[7];
  assign o[4017] = i[7];
  assign o[4018] = i[7];
  assign o[4019] = i[7];
  assign o[4020] = i[7];
  assign o[4021] = i[7];
  assign o[4022] = i[7];
  assign o[4023] = i[7];
  assign o[4024] = i[7];
  assign o[4025] = i[7];
  assign o[4026] = i[7];
  assign o[4027] = i[7];
  assign o[4028] = i[7];
  assign o[4029] = i[7];
  assign o[4030] = i[7];
  assign o[4031] = i[7];
  assign o[4032] = i[7];
  assign o[4033] = i[7];
  assign o[4034] = i[7];
  assign o[4035] = i[7];
  assign o[4036] = i[7];
  assign o[4037] = i[7];
  assign o[4038] = i[7];
  assign o[4039] = i[7];
  assign o[4040] = i[7];
  assign o[4041] = i[7];
  assign o[4042] = i[7];
  assign o[4043] = i[7];
  assign o[4044] = i[7];
  assign o[4045] = i[7];
  assign o[4046] = i[7];
  assign o[4047] = i[7];
  assign o[4048] = i[7];
  assign o[4049] = i[7];
  assign o[4050] = i[7];
  assign o[4051] = i[7];
  assign o[4052] = i[7];
  assign o[4053] = i[7];
  assign o[4054] = i[7];
  assign o[4055] = i[7];
  assign o[4056] = i[7];
  assign o[4057] = i[7];
  assign o[4058] = i[7];
  assign o[4059] = i[7];
  assign o[4060] = i[7];
  assign o[4061] = i[7];
  assign o[4062] = i[7];
  assign o[4063] = i[7];
  assign o[4064] = i[7];
  assign o[4065] = i[7];
  assign o[4066] = i[7];
  assign o[4067] = i[7];
  assign o[4068] = i[7];
  assign o[4069] = i[7];
  assign o[4070] = i[7];
  assign o[4071] = i[7];
  assign o[4072] = i[7];
  assign o[4073] = i[7];
  assign o[4074] = i[7];
  assign o[4075] = i[7];
  assign o[4076] = i[7];
  assign o[4077] = i[7];
  assign o[4078] = i[7];
  assign o[4079] = i[7];
  assign o[4080] = i[7];
  assign o[4081] = i[7];
  assign o[4082] = i[7];
  assign o[4083] = i[7];
  assign o[4084] = i[7];
  assign o[4085] = i[7];
  assign o[4086] = i[7];
  assign o[4087] = i[7];
  assign o[4088] = i[7];
  assign o[4089] = i[7];
  assign o[4090] = i[7];
  assign o[4091] = i[7];
  assign o[4092] = i[7];
  assign o[4093] = i[7];
  assign o[4094] = i[7];
  assign o[4095] = i[7];
  assign o[3072] = i[6];
  assign o[3073] = i[6];
  assign o[3074] = i[6];
  assign o[3075] = i[6];
  assign o[3076] = i[6];
  assign o[3077] = i[6];
  assign o[3078] = i[6];
  assign o[3079] = i[6];
  assign o[3080] = i[6];
  assign o[3081] = i[6];
  assign o[3082] = i[6];
  assign o[3083] = i[6];
  assign o[3084] = i[6];
  assign o[3085] = i[6];
  assign o[3086] = i[6];
  assign o[3087] = i[6];
  assign o[3088] = i[6];
  assign o[3089] = i[6];
  assign o[3090] = i[6];
  assign o[3091] = i[6];
  assign o[3092] = i[6];
  assign o[3093] = i[6];
  assign o[3094] = i[6];
  assign o[3095] = i[6];
  assign o[3096] = i[6];
  assign o[3097] = i[6];
  assign o[3098] = i[6];
  assign o[3099] = i[6];
  assign o[3100] = i[6];
  assign o[3101] = i[6];
  assign o[3102] = i[6];
  assign o[3103] = i[6];
  assign o[3104] = i[6];
  assign o[3105] = i[6];
  assign o[3106] = i[6];
  assign o[3107] = i[6];
  assign o[3108] = i[6];
  assign o[3109] = i[6];
  assign o[3110] = i[6];
  assign o[3111] = i[6];
  assign o[3112] = i[6];
  assign o[3113] = i[6];
  assign o[3114] = i[6];
  assign o[3115] = i[6];
  assign o[3116] = i[6];
  assign o[3117] = i[6];
  assign o[3118] = i[6];
  assign o[3119] = i[6];
  assign o[3120] = i[6];
  assign o[3121] = i[6];
  assign o[3122] = i[6];
  assign o[3123] = i[6];
  assign o[3124] = i[6];
  assign o[3125] = i[6];
  assign o[3126] = i[6];
  assign o[3127] = i[6];
  assign o[3128] = i[6];
  assign o[3129] = i[6];
  assign o[3130] = i[6];
  assign o[3131] = i[6];
  assign o[3132] = i[6];
  assign o[3133] = i[6];
  assign o[3134] = i[6];
  assign o[3135] = i[6];
  assign o[3136] = i[6];
  assign o[3137] = i[6];
  assign o[3138] = i[6];
  assign o[3139] = i[6];
  assign o[3140] = i[6];
  assign o[3141] = i[6];
  assign o[3142] = i[6];
  assign o[3143] = i[6];
  assign o[3144] = i[6];
  assign o[3145] = i[6];
  assign o[3146] = i[6];
  assign o[3147] = i[6];
  assign o[3148] = i[6];
  assign o[3149] = i[6];
  assign o[3150] = i[6];
  assign o[3151] = i[6];
  assign o[3152] = i[6];
  assign o[3153] = i[6];
  assign o[3154] = i[6];
  assign o[3155] = i[6];
  assign o[3156] = i[6];
  assign o[3157] = i[6];
  assign o[3158] = i[6];
  assign o[3159] = i[6];
  assign o[3160] = i[6];
  assign o[3161] = i[6];
  assign o[3162] = i[6];
  assign o[3163] = i[6];
  assign o[3164] = i[6];
  assign o[3165] = i[6];
  assign o[3166] = i[6];
  assign o[3167] = i[6];
  assign o[3168] = i[6];
  assign o[3169] = i[6];
  assign o[3170] = i[6];
  assign o[3171] = i[6];
  assign o[3172] = i[6];
  assign o[3173] = i[6];
  assign o[3174] = i[6];
  assign o[3175] = i[6];
  assign o[3176] = i[6];
  assign o[3177] = i[6];
  assign o[3178] = i[6];
  assign o[3179] = i[6];
  assign o[3180] = i[6];
  assign o[3181] = i[6];
  assign o[3182] = i[6];
  assign o[3183] = i[6];
  assign o[3184] = i[6];
  assign o[3185] = i[6];
  assign o[3186] = i[6];
  assign o[3187] = i[6];
  assign o[3188] = i[6];
  assign o[3189] = i[6];
  assign o[3190] = i[6];
  assign o[3191] = i[6];
  assign o[3192] = i[6];
  assign o[3193] = i[6];
  assign o[3194] = i[6];
  assign o[3195] = i[6];
  assign o[3196] = i[6];
  assign o[3197] = i[6];
  assign o[3198] = i[6];
  assign o[3199] = i[6];
  assign o[3200] = i[6];
  assign o[3201] = i[6];
  assign o[3202] = i[6];
  assign o[3203] = i[6];
  assign o[3204] = i[6];
  assign o[3205] = i[6];
  assign o[3206] = i[6];
  assign o[3207] = i[6];
  assign o[3208] = i[6];
  assign o[3209] = i[6];
  assign o[3210] = i[6];
  assign o[3211] = i[6];
  assign o[3212] = i[6];
  assign o[3213] = i[6];
  assign o[3214] = i[6];
  assign o[3215] = i[6];
  assign o[3216] = i[6];
  assign o[3217] = i[6];
  assign o[3218] = i[6];
  assign o[3219] = i[6];
  assign o[3220] = i[6];
  assign o[3221] = i[6];
  assign o[3222] = i[6];
  assign o[3223] = i[6];
  assign o[3224] = i[6];
  assign o[3225] = i[6];
  assign o[3226] = i[6];
  assign o[3227] = i[6];
  assign o[3228] = i[6];
  assign o[3229] = i[6];
  assign o[3230] = i[6];
  assign o[3231] = i[6];
  assign o[3232] = i[6];
  assign o[3233] = i[6];
  assign o[3234] = i[6];
  assign o[3235] = i[6];
  assign o[3236] = i[6];
  assign o[3237] = i[6];
  assign o[3238] = i[6];
  assign o[3239] = i[6];
  assign o[3240] = i[6];
  assign o[3241] = i[6];
  assign o[3242] = i[6];
  assign o[3243] = i[6];
  assign o[3244] = i[6];
  assign o[3245] = i[6];
  assign o[3246] = i[6];
  assign o[3247] = i[6];
  assign o[3248] = i[6];
  assign o[3249] = i[6];
  assign o[3250] = i[6];
  assign o[3251] = i[6];
  assign o[3252] = i[6];
  assign o[3253] = i[6];
  assign o[3254] = i[6];
  assign o[3255] = i[6];
  assign o[3256] = i[6];
  assign o[3257] = i[6];
  assign o[3258] = i[6];
  assign o[3259] = i[6];
  assign o[3260] = i[6];
  assign o[3261] = i[6];
  assign o[3262] = i[6];
  assign o[3263] = i[6];
  assign o[3264] = i[6];
  assign o[3265] = i[6];
  assign o[3266] = i[6];
  assign o[3267] = i[6];
  assign o[3268] = i[6];
  assign o[3269] = i[6];
  assign o[3270] = i[6];
  assign o[3271] = i[6];
  assign o[3272] = i[6];
  assign o[3273] = i[6];
  assign o[3274] = i[6];
  assign o[3275] = i[6];
  assign o[3276] = i[6];
  assign o[3277] = i[6];
  assign o[3278] = i[6];
  assign o[3279] = i[6];
  assign o[3280] = i[6];
  assign o[3281] = i[6];
  assign o[3282] = i[6];
  assign o[3283] = i[6];
  assign o[3284] = i[6];
  assign o[3285] = i[6];
  assign o[3286] = i[6];
  assign o[3287] = i[6];
  assign o[3288] = i[6];
  assign o[3289] = i[6];
  assign o[3290] = i[6];
  assign o[3291] = i[6];
  assign o[3292] = i[6];
  assign o[3293] = i[6];
  assign o[3294] = i[6];
  assign o[3295] = i[6];
  assign o[3296] = i[6];
  assign o[3297] = i[6];
  assign o[3298] = i[6];
  assign o[3299] = i[6];
  assign o[3300] = i[6];
  assign o[3301] = i[6];
  assign o[3302] = i[6];
  assign o[3303] = i[6];
  assign o[3304] = i[6];
  assign o[3305] = i[6];
  assign o[3306] = i[6];
  assign o[3307] = i[6];
  assign o[3308] = i[6];
  assign o[3309] = i[6];
  assign o[3310] = i[6];
  assign o[3311] = i[6];
  assign o[3312] = i[6];
  assign o[3313] = i[6];
  assign o[3314] = i[6];
  assign o[3315] = i[6];
  assign o[3316] = i[6];
  assign o[3317] = i[6];
  assign o[3318] = i[6];
  assign o[3319] = i[6];
  assign o[3320] = i[6];
  assign o[3321] = i[6];
  assign o[3322] = i[6];
  assign o[3323] = i[6];
  assign o[3324] = i[6];
  assign o[3325] = i[6];
  assign o[3326] = i[6];
  assign o[3327] = i[6];
  assign o[3328] = i[6];
  assign o[3329] = i[6];
  assign o[3330] = i[6];
  assign o[3331] = i[6];
  assign o[3332] = i[6];
  assign o[3333] = i[6];
  assign o[3334] = i[6];
  assign o[3335] = i[6];
  assign o[3336] = i[6];
  assign o[3337] = i[6];
  assign o[3338] = i[6];
  assign o[3339] = i[6];
  assign o[3340] = i[6];
  assign o[3341] = i[6];
  assign o[3342] = i[6];
  assign o[3343] = i[6];
  assign o[3344] = i[6];
  assign o[3345] = i[6];
  assign o[3346] = i[6];
  assign o[3347] = i[6];
  assign o[3348] = i[6];
  assign o[3349] = i[6];
  assign o[3350] = i[6];
  assign o[3351] = i[6];
  assign o[3352] = i[6];
  assign o[3353] = i[6];
  assign o[3354] = i[6];
  assign o[3355] = i[6];
  assign o[3356] = i[6];
  assign o[3357] = i[6];
  assign o[3358] = i[6];
  assign o[3359] = i[6];
  assign o[3360] = i[6];
  assign o[3361] = i[6];
  assign o[3362] = i[6];
  assign o[3363] = i[6];
  assign o[3364] = i[6];
  assign o[3365] = i[6];
  assign o[3366] = i[6];
  assign o[3367] = i[6];
  assign o[3368] = i[6];
  assign o[3369] = i[6];
  assign o[3370] = i[6];
  assign o[3371] = i[6];
  assign o[3372] = i[6];
  assign o[3373] = i[6];
  assign o[3374] = i[6];
  assign o[3375] = i[6];
  assign o[3376] = i[6];
  assign o[3377] = i[6];
  assign o[3378] = i[6];
  assign o[3379] = i[6];
  assign o[3380] = i[6];
  assign o[3381] = i[6];
  assign o[3382] = i[6];
  assign o[3383] = i[6];
  assign o[3384] = i[6];
  assign o[3385] = i[6];
  assign o[3386] = i[6];
  assign o[3387] = i[6];
  assign o[3388] = i[6];
  assign o[3389] = i[6];
  assign o[3390] = i[6];
  assign o[3391] = i[6];
  assign o[3392] = i[6];
  assign o[3393] = i[6];
  assign o[3394] = i[6];
  assign o[3395] = i[6];
  assign o[3396] = i[6];
  assign o[3397] = i[6];
  assign o[3398] = i[6];
  assign o[3399] = i[6];
  assign o[3400] = i[6];
  assign o[3401] = i[6];
  assign o[3402] = i[6];
  assign o[3403] = i[6];
  assign o[3404] = i[6];
  assign o[3405] = i[6];
  assign o[3406] = i[6];
  assign o[3407] = i[6];
  assign o[3408] = i[6];
  assign o[3409] = i[6];
  assign o[3410] = i[6];
  assign o[3411] = i[6];
  assign o[3412] = i[6];
  assign o[3413] = i[6];
  assign o[3414] = i[6];
  assign o[3415] = i[6];
  assign o[3416] = i[6];
  assign o[3417] = i[6];
  assign o[3418] = i[6];
  assign o[3419] = i[6];
  assign o[3420] = i[6];
  assign o[3421] = i[6];
  assign o[3422] = i[6];
  assign o[3423] = i[6];
  assign o[3424] = i[6];
  assign o[3425] = i[6];
  assign o[3426] = i[6];
  assign o[3427] = i[6];
  assign o[3428] = i[6];
  assign o[3429] = i[6];
  assign o[3430] = i[6];
  assign o[3431] = i[6];
  assign o[3432] = i[6];
  assign o[3433] = i[6];
  assign o[3434] = i[6];
  assign o[3435] = i[6];
  assign o[3436] = i[6];
  assign o[3437] = i[6];
  assign o[3438] = i[6];
  assign o[3439] = i[6];
  assign o[3440] = i[6];
  assign o[3441] = i[6];
  assign o[3442] = i[6];
  assign o[3443] = i[6];
  assign o[3444] = i[6];
  assign o[3445] = i[6];
  assign o[3446] = i[6];
  assign o[3447] = i[6];
  assign o[3448] = i[6];
  assign o[3449] = i[6];
  assign o[3450] = i[6];
  assign o[3451] = i[6];
  assign o[3452] = i[6];
  assign o[3453] = i[6];
  assign o[3454] = i[6];
  assign o[3455] = i[6];
  assign o[3456] = i[6];
  assign o[3457] = i[6];
  assign o[3458] = i[6];
  assign o[3459] = i[6];
  assign o[3460] = i[6];
  assign o[3461] = i[6];
  assign o[3462] = i[6];
  assign o[3463] = i[6];
  assign o[3464] = i[6];
  assign o[3465] = i[6];
  assign o[3466] = i[6];
  assign o[3467] = i[6];
  assign o[3468] = i[6];
  assign o[3469] = i[6];
  assign o[3470] = i[6];
  assign o[3471] = i[6];
  assign o[3472] = i[6];
  assign o[3473] = i[6];
  assign o[3474] = i[6];
  assign o[3475] = i[6];
  assign o[3476] = i[6];
  assign o[3477] = i[6];
  assign o[3478] = i[6];
  assign o[3479] = i[6];
  assign o[3480] = i[6];
  assign o[3481] = i[6];
  assign o[3482] = i[6];
  assign o[3483] = i[6];
  assign o[3484] = i[6];
  assign o[3485] = i[6];
  assign o[3486] = i[6];
  assign o[3487] = i[6];
  assign o[3488] = i[6];
  assign o[3489] = i[6];
  assign o[3490] = i[6];
  assign o[3491] = i[6];
  assign o[3492] = i[6];
  assign o[3493] = i[6];
  assign o[3494] = i[6];
  assign o[3495] = i[6];
  assign o[3496] = i[6];
  assign o[3497] = i[6];
  assign o[3498] = i[6];
  assign o[3499] = i[6];
  assign o[3500] = i[6];
  assign o[3501] = i[6];
  assign o[3502] = i[6];
  assign o[3503] = i[6];
  assign o[3504] = i[6];
  assign o[3505] = i[6];
  assign o[3506] = i[6];
  assign o[3507] = i[6];
  assign o[3508] = i[6];
  assign o[3509] = i[6];
  assign o[3510] = i[6];
  assign o[3511] = i[6];
  assign o[3512] = i[6];
  assign o[3513] = i[6];
  assign o[3514] = i[6];
  assign o[3515] = i[6];
  assign o[3516] = i[6];
  assign o[3517] = i[6];
  assign o[3518] = i[6];
  assign o[3519] = i[6];
  assign o[3520] = i[6];
  assign o[3521] = i[6];
  assign o[3522] = i[6];
  assign o[3523] = i[6];
  assign o[3524] = i[6];
  assign o[3525] = i[6];
  assign o[3526] = i[6];
  assign o[3527] = i[6];
  assign o[3528] = i[6];
  assign o[3529] = i[6];
  assign o[3530] = i[6];
  assign o[3531] = i[6];
  assign o[3532] = i[6];
  assign o[3533] = i[6];
  assign o[3534] = i[6];
  assign o[3535] = i[6];
  assign o[3536] = i[6];
  assign o[3537] = i[6];
  assign o[3538] = i[6];
  assign o[3539] = i[6];
  assign o[3540] = i[6];
  assign o[3541] = i[6];
  assign o[3542] = i[6];
  assign o[3543] = i[6];
  assign o[3544] = i[6];
  assign o[3545] = i[6];
  assign o[3546] = i[6];
  assign o[3547] = i[6];
  assign o[3548] = i[6];
  assign o[3549] = i[6];
  assign o[3550] = i[6];
  assign o[3551] = i[6];
  assign o[3552] = i[6];
  assign o[3553] = i[6];
  assign o[3554] = i[6];
  assign o[3555] = i[6];
  assign o[3556] = i[6];
  assign o[3557] = i[6];
  assign o[3558] = i[6];
  assign o[3559] = i[6];
  assign o[3560] = i[6];
  assign o[3561] = i[6];
  assign o[3562] = i[6];
  assign o[3563] = i[6];
  assign o[3564] = i[6];
  assign o[3565] = i[6];
  assign o[3566] = i[6];
  assign o[3567] = i[6];
  assign o[3568] = i[6];
  assign o[3569] = i[6];
  assign o[3570] = i[6];
  assign o[3571] = i[6];
  assign o[3572] = i[6];
  assign o[3573] = i[6];
  assign o[3574] = i[6];
  assign o[3575] = i[6];
  assign o[3576] = i[6];
  assign o[3577] = i[6];
  assign o[3578] = i[6];
  assign o[3579] = i[6];
  assign o[3580] = i[6];
  assign o[3581] = i[6];
  assign o[3582] = i[6];
  assign o[3583] = i[6];
  assign o[2560] = i[5];
  assign o[2561] = i[5];
  assign o[2562] = i[5];
  assign o[2563] = i[5];
  assign o[2564] = i[5];
  assign o[2565] = i[5];
  assign o[2566] = i[5];
  assign o[2567] = i[5];
  assign o[2568] = i[5];
  assign o[2569] = i[5];
  assign o[2570] = i[5];
  assign o[2571] = i[5];
  assign o[2572] = i[5];
  assign o[2573] = i[5];
  assign o[2574] = i[5];
  assign o[2575] = i[5];
  assign o[2576] = i[5];
  assign o[2577] = i[5];
  assign o[2578] = i[5];
  assign o[2579] = i[5];
  assign o[2580] = i[5];
  assign o[2581] = i[5];
  assign o[2582] = i[5];
  assign o[2583] = i[5];
  assign o[2584] = i[5];
  assign o[2585] = i[5];
  assign o[2586] = i[5];
  assign o[2587] = i[5];
  assign o[2588] = i[5];
  assign o[2589] = i[5];
  assign o[2590] = i[5];
  assign o[2591] = i[5];
  assign o[2592] = i[5];
  assign o[2593] = i[5];
  assign o[2594] = i[5];
  assign o[2595] = i[5];
  assign o[2596] = i[5];
  assign o[2597] = i[5];
  assign o[2598] = i[5];
  assign o[2599] = i[5];
  assign o[2600] = i[5];
  assign o[2601] = i[5];
  assign o[2602] = i[5];
  assign o[2603] = i[5];
  assign o[2604] = i[5];
  assign o[2605] = i[5];
  assign o[2606] = i[5];
  assign o[2607] = i[5];
  assign o[2608] = i[5];
  assign o[2609] = i[5];
  assign o[2610] = i[5];
  assign o[2611] = i[5];
  assign o[2612] = i[5];
  assign o[2613] = i[5];
  assign o[2614] = i[5];
  assign o[2615] = i[5];
  assign o[2616] = i[5];
  assign o[2617] = i[5];
  assign o[2618] = i[5];
  assign o[2619] = i[5];
  assign o[2620] = i[5];
  assign o[2621] = i[5];
  assign o[2622] = i[5];
  assign o[2623] = i[5];
  assign o[2624] = i[5];
  assign o[2625] = i[5];
  assign o[2626] = i[5];
  assign o[2627] = i[5];
  assign o[2628] = i[5];
  assign o[2629] = i[5];
  assign o[2630] = i[5];
  assign o[2631] = i[5];
  assign o[2632] = i[5];
  assign o[2633] = i[5];
  assign o[2634] = i[5];
  assign o[2635] = i[5];
  assign o[2636] = i[5];
  assign o[2637] = i[5];
  assign o[2638] = i[5];
  assign o[2639] = i[5];
  assign o[2640] = i[5];
  assign o[2641] = i[5];
  assign o[2642] = i[5];
  assign o[2643] = i[5];
  assign o[2644] = i[5];
  assign o[2645] = i[5];
  assign o[2646] = i[5];
  assign o[2647] = i[5];
  assign o[2648] = i[5];
  assign o[2649] = i[5];
  assign o[2650] = i[5];
  assign o[2651] = i[5];
  assign o[2652] = i[5];
  assign o[2653] = i[5];
  assign o[2654] = i[5];
  assign o[2655] = i[5];
  assign o[2656] = i[5];
  assign o[2657] = i[5];
  assign o[2658] = i[5];
  assign o[2659] = i[5];
  assign o[2660] = i[5];
  assign o[2661] = i[5];
  assign o[2662] = i[5];
  assign o[2663] = i[5];
  assign o[2664] = i[5];
  assign o[2665] = i[5];
  assign o[2666] = i[5];
  assign o[2667] = i[5];
  assign o[2668] = i[5];
  assign o[2669] = i[5];
  assign o[2670] = i[5];
  assign o[2671] = i[5];
  assign o[2672] = i[5];
  assign o[2673] = i[5];
  assign o[2674] = i[5];
  assign o[2675] = i[5];
  assign o[2676] = i[5];
  assign o[2677] = i[5];
  assign o[2678] = i[5];
  assign o[2679] = i[5];
  assign o[2680] = i[5];
  assign o[2681] = i[5];
  assign o[2682] = i[5];
  assign o[2683] = i[5];
  assign o[2684] = i[5];
  assign o[2685] = i[5];
  assign o[2686] = i[5];
  assign o[2687] = i[5];
  assign o[2688] = i[5];
  assign o[2689] = i[5];
  assign o[2690] = i[5];
  assign o[2691] = i[5];
  assign o[2692] = i[5];
  assign o[2693] = i[5];
  assign o[2694] = i[5];
  assign o[2695] = i[5];
  assign o[2696] = i[5];
  assign o[2697] = i[5];
  assign o[2698] = i[5];
  assign o[2699] = i[5];
  assign o[2700] = i[5];
  assign o[2701] = i[5];
  assign o[2702] = i[5];
  assign o[2703] = i[5];
  assign o[2704] = i[5];
  assign o[2705] = i[5];
  assign o[2706] = i[5];
  assign o[2707] = i[5];
  assign o[2708] = i[5];
  assign o[2709] = i[5];
  assign o[2710] = i[5];
  assign o[2711] = i[5];
  assign o[2712] = i[5];
  assign o[2713] = i[5];
  assign o[2714] = i[5];
  assign o[2715] = i[5];
  assign o[2716] = i[5];
  assign o[2717] = i[5];
  assign o[2718] = i[5];
  assign o[2719] = i[5];
  assign o[2720] = i[5];
  assign o[2721] = i[5];
  assign o[2722] = i[5];
  assign o[2723] = i[5];
  assign o[2724] = i[5];
  assign o[2725] = i[5];
  assign o[2726] = i[5];
  assign o[2727] = i[5];
  assign o[2728] = i[5];
  assign o[2729] = i[5];
  assign o[2730] = i[5];
  assign o[2731] = i[5];
  assign o[2732] = i[5];
  assign o[2733] = i[5];
  assign o[2734] = i[5];
  assign o[2735] = i[5];
  assign o[2736] = i[5];
  assign o[2737] = i[5];
  assign o[2738] = i[5];
  assign o[2739] = i[5];
  assign o[2740] = i[5];
  assign o[2741] = i[5];
  assign o[2742] = i[5];
  assign o[2743] = i[5];
  assign o[2744] = i[5];
  assign o[2745] = i[5];
  assign o[2746] = i[5];
  assign o[2747] = i[5];
  assign o[2748] = i[5];
  assign o[2749] = i[5];
  assign o[2750] = i[5];
  assign o[2751] = i[5];
  assign o[2752] = i[5];
  assign o[2753] = i[5];
  assign o[2754] = i[5];
  assign o[2755] = i[5];
  assign o[2756] = i[5];
  assign o[2757] = i[5];
  assign o[2758] = i[5];
  assign o[2759] = i[5];
  assign o[2760] = i[5];
  assign o[2761] = i[5];
  assign o[2762] = i[5];
  assign o[2763] = i[5];
  assign o[2764] = i[5];
  assign o[2765] = i[5];
  assign o[2766] = i[5];
  assign o[2767] = i[5];
  assign o[2768] = i[5];
  assign o[2769] = i[5];
  assign o[2770] = i[5];
  assign o[2771] = i[5];
  assign o[2772] = i[5];
  assign o[2773] = i[5];
  assign o[2774] = i[5];
  assign o[2775] = i[5];
  assign o[2776] = i[5];
  assign o[2777] = i[5];
  assign o[2778] = i[5];
  assign o[2779] = i[5];
  assign o[2780] = i[5];
  assign o[2781] = i[5];
  assign o[2782] = i[5];
  assign o[2783] = i[5];
  assign o[2784] = i[5];
  assign o[2785] = i[5];
  assign o[2786] = i[5];
  assign o[2787] = i[5];
  assign o[2788] = i[5];
  assign o[2789] = i[5];
  assign o[2790] = i[5];
  assign o[2791] = i[5];
  assign o[2792] = i[5];
  assign o[2793] = i[5];
  assign o[2794] = i[5];
  assign o[2795] = i[5];
  assign o[2796] = i[5];
  assign o[2797] = i[5];
  assign o[2798] = i[5];
  assign o[2799] = i[5];
  assign o[2800] = i[5];
  assign o[2801] = i[5];
  assign o[2802] = i[5];
  assign o[2803] = i[5];
  assign o[2804] = i[5];
  assign o[2805] = i[5];
  assign o[2806] = i[5];
  assign o[2807] = i[5];
  assign o[2808] = i[5];
  assign o[2809] = i[5];
  assign o[2810] = i[5];
  assign o[2811] = i[5];
  assign o[2812] = i[5];
  assign o[2813] = i[5];
  assign o[2814] = i[5];
  assign o[2815] = i[5];
  assign o[2816] = i[5];
  assign o[2817] = i[5];
  assign o[2818] = i[5];
  assign o[2819] = i[5];
  assign o[2820] = i[5];
  assign o[2821] = i[5];
  assign o[2822] = i[5];
  assign o[2823] = i[5];
  assign o[2824] = i[5];
  assign o[2825] = i[5];
  assign o[2826] = i[5];
  assign o[2827] = i[5];
  assign o[2828] = i[5];
  assign o[2829] = i[5];
  assign o[2830] = i[5];
  assign o[2831] = i[5];
  assign o[2832] = i[5];
  assign o[2833] = i[5];
  assign o[2834] = i[5];
  assign o[2835] = i[5];
  assign o[2836] = i[5];
  assign o[2837] = i[5];
  assign o[2838] = i[5];
  assign o[2839] = i[5];
  assign o[2840] = i[5];
  assign o[2841] = i[5];
  assign o[2842] = i[5];
  assign o[2843] = i[5];
  assign o[2844] = i[5];
  assign o[2845] = i[5];
  assign o[2846] = i[5];
  assign o[2847] = i[5];
  assign o[2848] = i[5];
  assign o[2849] = i[5];
  assign o[2850] = i[5];
  assign o[2851] = i[5];
  assign o[2852] = i[5];
  assign o[2853] = i[5];
  assign o[2854] = i[5];
  assign o[2855] = i[5];
  assign o[2856] = i[5];
  assign o[2857] = i[5];
  assign o[2858] = i[5];
  assign o[2859] = i[5];
  assign o[2860] = i[5];
  assign o[2861] = i[5];
  assign o[2862] = i[5];
  assign o[2863] = i[5];
  assign o[2864] = i[5];
  assign o[2865] = i[5];
  assign o[2866] = i[5];
  assign o[2867] = i[5];
  assign o[2868] = i[5];
  assign o[2869] = i[5];
  assign o[2870] = i[5];
  assign o[2871] = i[5];
  assign o[2872] = i[5];
  assign o[2873] = i[5];
  assign o[2874] = i[5];
  assign o[2875] = i[5];
  assign o[2876] = i[5];
  assign o[2877] = i[5];
  assign o[2878] = i[5];
  assign o[2879] = i[5];
  assign o[2880] = i[5];
  assign o[2881] = i[5];
  assign o[2882] = i[5];
  assign o[2883] = i[5];
  assign o[2884] = i[5];
  assign o[2885] = i[5];
  assign o[2886] = i[5];
  assign o[2887] = i[5];
  assign o[2888] = i[5];
  assign o[2889] = i[5];
  assign o[2890] = i[5];
  assign o[2891] = i[5];
  assign o[2892] = i[5];
  assign o[2893] = i[5];
  assign o[2894] = i[5];
  assign o[2895] = i[5];
  assign o[2896] = i[5];
  assign o[2897] = i[5];
  assign o[2898] = i[5];
  assign o[2899] = i[5];
  assign o[2900] = i[5];
  assign o[2901] = i[5];
  assign o[2902] = i[5];
  assign o[2903] = i[5];
  assign o[2904] = i[5];
  assign o[2905] = i[5];
  assign o[2906] = i[5];
  assign o[2907] = i[5];
  assign o[2908] = i[5];
  assign o[2909] = i[5];
  assign o[2910] = i[5];
  assign o[2911] = i[5];
  assign o[2912] = i[5];
  assign o[2913] = i[5];
  assign o[2914] = i[5];
  assign o[2915] = i[5];
  assign o[2916] = i[5];
  assign o[2917] = i[5];
  assign o[2918] = i[5];
  assign o[2919] = i[5];
  assign o[2920] = i[5];
  assign o[2921] = i[5];
  assign o[2922] = i[5];
  assign o[2923] = i[5];
  assign o[2924] = i[5];
  assign o[2925] = i[5];
  assign o[2926] = i[5];
  assign o[2927] = i[5];
  assign o[2928] = i[5];
  assign o[2929] = i[5];
  assign o[2930] = i[5];
  assign o[2931] = i[5];
  assign o[2932] = i[5];
  assign o[2933] = i[5];
  assign o[2934] = i[5];
  assign o[2935] = i[5];
  assign o[2936] = i[5];
  assign o[2937] = i[5];
  assign o[2938] = i[5];
  assign o[2939] = i[5];
  assign o[2940] = i[5];
  assign o[2941] = i[5];
  assign o[2942] = i[5];
  assign o[2943] = i[5];
  assign o[2944] = i[5];
  assign o[2945] = i[5];
  assign o[2946] = i[5];
  assign o[2947] = i[5];
  assign o[2948] = i[5];
  assign o[2949] = i[5];
  assign o[2950] = i[5];
  assign o[2951] = i[5];
  assign o[2952] = i[5];
  assign o[2953] = i[5];
  assign o[2954] = i[5];
  assign o[2955] = i[5];
  assign o[2956] = i[5];
  assign o[2957] = i[5];
  assign o[2958] = i[5];
  assign o[2959] = i[5];
  assign o[2960] = i[5];
  assign o[2961] = i[5];
  assign o[2962] = i[5];
  assign o[2963] = i[5];
  assign o[2964] = i[5];
  assign o[2965] = i[5];
  assign o[2966] = i[5];
  assign o[2967] = i[5];
  assign o[2968] = i[5];
  assign o[2969] = i[5];
  assign o[2970] = i[5];
  assign o[2971] = i[5];
  assign o[2972] = i[5];
  assign o[2973] = i[5];
  assign o[2974] = i[5];
  assign o[2975] = i[5];
  assign o[2976] = i[5];
  assign o[2977] = i[5];
  assign o[2978] = i[5];
  assign o[2979] = i[5];
  assign o[2980] = i[5];
  assign o[2981] = i[5];
  assign o[2982] = i[5];
  assign o[2983] = i[5];
  assign o[2984] = i[5];
  assign o[2985] = i[5];
  assign o[2986] = i[5];
  assign o[2987] = i[5];
  assign o[2988] = i[5];
  assign o[2989] = i[5];
  assign o[2990] = i[5];
  assign o[2991] = i[5];
  assign o[2992] = i[5];
  assign o[2993] = i[5];
  assign o[2994] = i[5];
  assign o[2995] = i[5];
  assign o[2996] = i[5];
  assign o[2997] = i[5];
  assign o[2998] = i[5];
  assign o[2999] = i[5];
  assign o[3000] = i[5];
  assign o[3001] = i[5];
  assign o[3002] = i[5];
  assign o[3003] = i[5];
  assign o[3004] = i[5];
  assign o[3005] = i[5];
  assign o[3006] = i[5];
  assign o[3007] = i[5];
  assign o[3008] = i[5];
  assign o[3009] = i[5];
  assign o[3010] = i[5];
  assign o[3011] = i[5];
  assign o[3012] = i[5];
  assign o[3013] = i[5];
  assign o[3014] = i[5];
  assign o[3015] = i[5];
  assign o[3016] = i[5];
  assign o[3017] = i[5];
  assign o[3018] = i[5];
  assign o[3019] = i[5];
  assign o[3020] = i[5];
  assign o[3021] = i[5];
  assign o[3022] = i[5];
  assign o[3023] = i[5];
  assign o[3024] = i[5];
  assign o[3025] = i[5];
  assign o[3026] = i[5];
  assign o[3027] = i[5];
  assign o[3028] = i[5];
  assign o[3029] = i[5];
  assign o[3030] = i[5];
  assign o[3031] = i[5];
  assign o[3032] = i[5];
  assign o[3033] = i[5];
  assign o[3034] = i[5];
  assign o[3035] = i[5];
  assign o[3036] = i[5];
  assign o[3037] = i[5];
  assign o[3038] = i[5];
  assign o[3039] = i[5];
  assign o[3040] = i[5];
  assign o[3041] = i[5];
  assign o[3042] = i[5];
  assign o[3043] = i[5];
  assign o[3044] = i[5];
  assign o[3045] = i[5];
  assign o[3046] = i[5];
  assign o[3047] = i[5];
  assign o[3048] = i[5];
  assign o[3049] = i[5];
  assign o[3050] = i[5];
  assign o[3051] = i[5];
  assign o[3052] = i[5];
  assign o[3053] = i[5];
  assign o[3054] = i[5];
  assign o[3055] = i[5];
  assign o[3056] = i[5];
  assign o[3057] = i[5];
  assign o[3058] = i[5];
  assign o[3059] = i[5];
  assign o[3060] = i[5];
  assign o[3061] = i[5];
  assign o[3062] = i[5];
  assign o[3063] = i[5];
  assign o[3064] = i[5];
  assign o[3065] = i[5];
  assign o[3066] = i[5];
  assign o[3067] = i[5];
  assign o[3068] = i[5];
  assign o[3069] = i[5];
  assign o[3070] = i[5];
  assign o[3071] = i[5];
  assign o[2048] = i[4];
  assign o[2049] = i[4];
  assign o[2050] = i[4];
  assign o[2051] = i[4];
  assign o[2052] = i[4];
  assign o[2053] = i[4];
  assign o[2054] = i[4];
  assign o[2055] = i[4];
  assign o[2056] = i[4];
  assign o[2057] = i[4];
  assign o[2058] = i[4];
  assign o[2059] = i[4];
  assign o[2060] = i[4];
  assign o[2061] = i[4];
  assign o[2062] = i[4];
  assign o[2063] = i[4];
  assign o[2064] = i[4];
  assign o[2065] = i[4];
  assign o[2066] = i[4];
  assign o[2067] = i[4];
  assign o[2068] = i[4];
  assign o[2069] = i[4];
  assign o[2070] = i[4];
  assign o[2071] = i[4];
  assign o[2072] = i[4];
  assign o[2073] = i[4];
  assign o[2074] = i[4];
  assign o[2075] = i[4];
  assign o[2076] = i[4];
  assign o[2077] = i[4];
  assign o[2078] = i[4];
  assign o[2079] = i[4];
  assign o[2080] = i[4];
  assign o[2081] = i[4];
  assign o[2082] = i[4];
  assign o[2083] = i[4];
  assign o[2084] = i[4];
  assign o[2085] = i[4];
  assign o[2086] = i[4];
  assign o[2087] = i[4];
  assign o[2088] = i[4];
  assign o[2089] = i[4];
  assign o[2090] = i[4];
  assign o[2091] = i[4];
  assign o[2092] = i[4];
  assign o[2093] = i[4];
  assign o[2094] = i[4];
  assign o[2095] = i[4];
  assign o[2096] = i[4];
  assign o[2097] = i[4];
  assign o[2098] = i[4];
  assign o[2099] = i[4];
  assign o[2100] = i[4];
  assign o[2101] = i[4];
  assign o[2102] = i[4];
  assign o[2103] = i[4];
  assign o[2104] = i[4];
  assign o[2105] = i[4];
  assign o[2106] = i[4];
  assign o[2107] = i[4];
  assign o[2108] = i[4];
  assign o[2109] = i[4];
  assign o[2110] = i[4];
  assign o[2111] = i[4];
  assign o[2112] = i[4];
  assign o[2113] = i[4];
  assign o[2114] = i[4];
  assign o[2115] = i[4];
  assign o[2116] = i[4];
  assign o[2117] = i[4];
  assign o[2118] = i[4];
  assign o[2119] = i[4];
  assign o[2120] = i[4];
  assign o[2121] = i[4];
  assign o[2122] = i[4];
  assign o[2123] = i[4];
  assign o[2124] = i[4];
  assign o[2125] = i[4];
  assign o[2126] = i[4];
  assign o[2127] = i[4];
  assign o[2128] = i[4];
  assign o[2129] = i[4];
  assign o[2130] = i[4];
  assign o[2131] = i[4];
  assign o[2132] = i[4];
  assign o[2133] = i[4];
  assign o[2134] = i[4];
  assign o[2135] = i[4];
  assign o[2136] = i[4];
  assign o[2137] = i[4];
  assign o[2138] = i[4];
  assign o[2139] = i[4];
  assign o[2140] = i[4];
  assign o[2141] = i[4];
  assign o[2142] = i[4];
  assign o[2143] = i[4];
  assign o[2144] = i[4];
  assign o[2145] = i[4];
  assign o[2146] = i[4];
  assign o[2147] = i[4];
  assign o[2148] = i[4];
  assign o[2149] = i[4];
  assign o[2150] = i[4];
  assign o[2151] = i[4];
  assign o[2152] = i[4];
  assign o[2153] = i[4];
  assign o[2154] = i[4];
  assign o[2155] = i[4];
  assign o[2156] = i[4];
  assign o[2157] = i[4];
  assign o[2158] = i[4];
  assign o[2159] = i[4];
  assign o[2160] = i[4];
  assign o[2161] = i[4];
  assign o[2162] = i[4];
  assign o[2163] = i[4];
  assign o[2164] = i[4];
  assign o[2165] = i[4];
  assign o[2166] = i[4];
  assign o[2167] = i[4];
  assign o[2168] = i[4];
  assign o[2169] = i[4];
  assign o[2170] = i[4];
  assign o[2171] = i[4];
  assign o[2172] = i[4];
  assign o[2173] = i[4];
  assign o[2174] = i[4];
  assign o[2175] = i[4];
  assign o[2176] = i[4];
  assign o[2177] = i[4];
  assign o[2178] = i[4];
  assign o[2179] = i[4];
  assign o[2180] = i[4];
  assign o[2181] = i[4];
  assign o[2182] = i[4];
  assign o[2183] = i[4];
  assign o[2184] = i[4];
  assign o[2185] = i[4];
  assign o[2186] = i[4];
  assign o[2187] = i[4];
  assign o[2188] = i[4];
  assign o[2189] = i[4];
  assign o[2190] = i[4];
  assign o[2191] = i[4];
  assign o[2192] = i[4];
  assign o[2193] = i[4];
  assign o[2194] = i[4];
  assign o[2195] = i[4];
  assign o[2196] = i[4];
  assign o[2197] = i[4];
  assign o[2198] = i[4];
  assign o[2199] = i[4];
  assign o[2200] = i[4];
  assign o[2201] = i[4];
  assign o[2202] = i[4];
  assign o[2203] = i[4];
  assign o[2204] = i[4];
  assign o[2205] = i[4];
  assign o[2206] = i[4];
  assign o[2207] = i[4];
  assign o[2208] = i[4];
  assign o[2209] = i[4];
  assign o[2210] = i[4];
  assign o[2211] = i[4];
  assign o[2212] = i[4];
  assign o[2213] = i[4];
  assign o[2214] = i[4];
  assign o[2215] = i[4];
  assign o[2216] = i[4];
  assign o[2217] = i[4];
  assign o[2218] = i[4];
  assign o[2219] = i[4];
  assign o[2220] = i[4];
  assign o[2221] = i[4];
  assign o[2222] = i[4];
  assign o[2223] = i[4];
  assign o[2224] = i[4];
  assign o[2225] = i[4];
  assign o[2226] = i[4];
  assign o[2227] = i[4];
  assign o[2228] = i[4];
  assign o[2229] = i[4];
  assign o[2230] = i[4];
  assign o[2231] = i[4];
  assign o[2232] = i[4];
  assign o[2233] = i[4];
  assign o[2234] = i[4];
  assign o[2235] = i[4];
  assign o[2236] = i[4];
  assign o[2237] = i[4];
  assign o[2238] = i[4];
  assign o[2239] = i[4];
  assign o[2240] = i[4];
  assign o[2241] = i[4];
  assign o[2242] = i[4];
  assign o[2243] = i[4];
  assign o[2244] = i[4];
  assign o[2245] = i[4];
  assign o[2246] = i[4];
  assign o[2247] = i[4];
  assign o[2248] = i[4];
  assign o[2249] = i[4];
  assign o[2250] = i[4];
  assign o[2251] = i[4];
  assign o[2252] = i[4];
  assign o[2253] = i[4];
  assign o[2254] = i[4];
  assign o[2255] = i[4];
  assign o[2256] = i[4];
  assign o[2257] = i[4];
  assign o[2258] = i[4];
  assign o[2259] = i[4];
  assign o[2260] = i[4];
  assign o[2261] = i[4];
  assign o[2262] = i[4];
  assign o[2263] = i[4];
  assign o[2264] = i[4];
  assign o[2265] = i[4];
  assign o[2266] = i[4];
  assign o[2267] = i[4];
  assign o[2268] = i[4];
  assign o[2269] = i[4];
  assign o[2270] = i[4];
  assign o[2271] = i[4];
  assign o[2272] = i[4];
  assign o[2273] = i[4];
  assign o[2274] = i[4];
  assign o[2275] = i[4];
  assign o[2276] = i[4];
  assign o[2277] = i[4];
  assign o[2278] = i[4];
  assign o[2279] = i[4];
  assign o[2280] = i[4];
  assign o[2281] = i[4];
  assign o[2282] = i[4];
  assign o[2283] = i[4];
  assign o[2284] = i[4];
  assign o[2285] = i[4];
  assign o[2286] = i[4];
  assign o[2287] = i[4];
  assign o[2288] = i[4];
  assign o[2289] = i[4];
  assign o[2290] = i[4];
  assign o[2291] = i[4];
  assign o[2292] = i[4];
  assign o[2293] = i[4];
  assign o[2294] = i[4];
  assign o[2295] = i[4];
  assign o[2296] = i[4];
  assign o[2297] = i[4];
  assign o[2298] = i[4];
  assign o[2299] = i[4];
  assign o[2300] = i[4];
  assign o[2301] = i[4];
  assign o[2302] = i[4];
  assign o[2303] = i[4];
  assign o[2304] = i[4];
  assign o[2305] = i[4];
  assign o[2306] = i[4];
  assign o[2307] = i[4];
  assign o[2308] = i[4];
  assign o[2309] = i[4];
  assign o[2310] = i[4];
  assign o[2311] = i[4];
  assign o[2312] = i[4];
  assign o[2313] = i[4];
  assign o[2314] = i[4];
  assign o[2315] = i[4];
  assign o[2316] = i[4];
  assign o[2317] = i[4];
  assign o[2318] = i[4];
  assign o[2319] = i[4];
  assign o[2320] = i[4];
  assign o[2321] = i[4];
  assign o[2322] = i[4];
  assign o[2323] = i[4];
  assign o[2324] = i[4];
  assign o[2325] = i[4];
  assign o[2326] = i[4];
  assign o[2327] = i[4];
  assign o[2328] = i[4];
  assign o[2329] = i[4];
  assign o[2330] = i[4];
  assign o[2331] = i[4];
  assign o[2332] = i[4];
  assign o[2333] = i[4];
  assign o[2334] = i[4];
  assign o[2335] = i[4];
  assign o[2336] = i[4];
  assign o[2337] = i[4];
  assign o[2338] = i[4];
  assign o[2339] = i[4];
  assign o[2340] = i[4];
  assign o[2341] = i[4];
  assign o[2342] = i[4];
  assign o[2343] = i[4];
  assign o[2344] = i[4];
  assign o[2345] = i[4];
  assign o[2346] = i[4];
  assign o[2347] = i[4];
  assign o[2348] = i[4];
  assign o[2349] = i[4];
  assign o[2350] = i[4];
  assign o[2351] = i[4];
  assign o[2352] = i[4];
  assign o[2353] = i[4];
  assign o[2354] = i[4];
  assign o[2355] = i[4];
  assign o[2356] = i[4];
  assign o[2357] = i[4];
  assign o[2358] = i[4];
  assign o[2359] = i[4];
  assign o[2360] = i[4];
  assign o[2361] = i[4];
  assign o[2362] = i[4];
  assign o[2363] = i[4];
  assign o[2364] = i[4];
  assign o[2365] = i[4];
  assign o[2366] = i[4];
  assign o[2367] = i[4];
  assign o[2368] = i[4];
  assign o[2369] = i[4];
  assign o[2370] = i[4];
  assign o[2371] = i[4];
  assign o[2372] = i[4];
  assign o[2373] = i[4];
  assign o[2374] = i[4];
  assign o[2375] = i[4];
  assign o[2376] = i[4];
  assign o[2377] = i[4];
  assign o[2378] = i[4];
  assign o[2379] = i[4];
  assign o[2380] = i[4];
  assign o[2381] = i[4];
  assign o[2382] = i[4];
  assign o[2383] = i[4];
  assign o[2384] = i[4];
  assign o[2385] = i[4];
  assign o[2386] = i[4];
  assign o[2387] = i[4];
  assign o[2388] = i[4];
  assign o[2389] = i[4];
  assign o[2390] = i[4];
  assign o[2391] = i[4];
  assign o[2392] = i[4];
  assign o[2393] = i[4];
  assign o[2394] = i[4];
  assign o[2395] = i[4];
  assign o[2396] = i[4];
  assign o[2397] = i[4];
  assign o[2398] = i[4];
  assign o[2399] = i[4];
  assign o[2400] = i[4];
  assign o[2401] = i[4];
  assign o[2402] = i[4];
  assign o[2403] = i[4];
  assign o[2404] = i[4];
  assign o[2405] = i[4];
  assign o[2406] = i[4];
  assign o[2407] = i[4];
  assign o[2408] = i[4];
  assign o[2409] = i[4];
  assign o[2410] = i[4];
  assign o[2411] = i[4];
  assign o[2412] = i[4];
  assign o[2413] = i[4];
  assign o[2414] = i[4];
  assign o[2415] = i[4];
  assign o[2416] = i[4];
  assign o[2417] = i[4];
  assign o[2418] = i[4];
  assign o[2419] = i[4];
  assign o[2420] = i[4];
  assign o[2421] = i[4];
  assign o[2422] = i[4];
  assign o[2423] = i[4];
  assign o[2424] = i[4];
  assign o[2425] = i[4];
  assign o[2426] = i[4];
  assign o[2427] = i[4];
  assign o[2428] = i[4];
  assign o[2429] = i[4];
  assign o[2430] = i[4];
  assign o[2431] = i[4];
  assign o[2432] = i[4];
  assign o[2433] = i[4];
  assign o[2434] = i[4];
  assign o[2435] = i[4];
  assign o[2436] = i[4];
  assign o[2437] = i[4];
  assign o[2438] = i[4];
  assign o[2439] = i[4];
  assign o[2440] = i[4];
  assign o[2441] = i[4];
  assign o[2442] = i[4];
  assign o[2443] = i[4];
  assign o[2444] = i[4];
  assign o[2445] = i[4];
  assign o[2446] = i[4];
  assign o[2447] = i[4];
  assign o[2448] = i[4];
  assign o[2449] = i[4];
  assign o[2450] = i[4];
  assign o[2451] = i[4];
  assign o[2452] = i[4];
  assign o[2453] = i[4];
  assign o[2454] = i[4];
  assign o[2455] = i[4];
  assign o[2456] = i[4];
  assign o[2457] = i[4];
  assign o[2458] = i[4];
  assign o[2459] = i[4];
  assign o[2460] = i[4];
  assign o[2461] = i[4];
  assign o[2462] = i[4];
  assign o[2463] = i[4];
  assign o[2464] = i[4];
  assign o[2465] = i[4];
  assign o[2466] = i[4];
  assign o[2467] = i[4];
  assign o[2468] = i[4];
  assign o[2469] = i[4];
  assign o[2470] = i[4];
  assign o[2471] = i[4];
  assign o[2472] = i[4];
  assign o[2473] = i[4];
  assign o[2474] = i[4];
  assign o[2475] = i[4];
  assign o[2476] = i[4];
  assign o[2477] = i[4];
  assign o[2478] = i[4];
  assign o[2479] = i[4];
  assign o[2480] = i[4];
  assign o[2481] = i[4];
  assign o[2482] = i[4];
  assign o[2483] = i[4];
  assign o[2484] = i[4];
  assign o[2485] = i[4];
  assign o[2486] = i[4];
  assign o[2487] = i[4];
  assign o[2488] = i[4];
  assign o[2489] = i[4];
  assign o[2490] = i[4];
  assign o[2491] = i[4];
  assign o[2492] = i[4];
  assign o[2493] = i[4];
  assign o[2494] = i[4];
  assign o[2495] = i[4];
  assign o[2496] = i[4];
  assign o[2497] = i[4];
  assign o[2498] = i[4];
  assign o[2499] = i[4];
  assign o[2500] = i[4];
  assign o[2501] = i[4];
  assign o[2502] = i[4];
  assign o[2503] = i[4];
  assign o[2504] = i[4];
  assign o[2505] = i[4];
  assign o[2506] = i[4];
  assign o[2507] = i[4];
  assign o[2508] = i[4];
  assign o[2509] = i[4];
  assign o[2510] = i[4];
  assign o[2511] = i[4];
  assign o[2512] = i[4];
  assign o[2513] = i[4];
  assign o[2514] = i[4];
  assign o[2515] = i[4];
  assign o[2516] = i[4];
  assign o[2517] = i[4];
  assign o[2518] = i[4];
  assign o[2519] = i[4];
  assign o[2520] = i[4];
  assign o[2521] = i[4];
  assign o[2522] = i[4];
  assign o[2523] = i[4];
  assign o[2524] = i[4];
  assign o[2525] = i[4];
  assign o[2526] = i[4];
  assign o[2527] = i[4];
  assign o[2528] = i[4];
  assign o[2529] = i[4];
  assign o[2530] = i[4];
  assign o[2531] = i[4];
  assign o[2532] = i[4];
  assign o[2533] = i[4];
  assign o[2534] = i[4];
  assign o[2535] = i[4];
  assign o[2536] = i[4];
  assign o[2537] = i[4];
  assign o[2538] = i[4];
  assign o[2539] = i[4];
  assign o[2540] = i[4];
  assign o[2541] = i[4];
  assign o[2542] = i[4];
  assign o[2543] = i[4];
  assign o[2544] = i[4];
  assign o[2545] = i[4];
  assign o[2546] = i[4];
  assign o[2547] = i[4];
  assign o[2548] = i[4];
  assign o[2549] = i[4];
  assign o[2550] = i[4];
  assign o[2551] = i[4];
  assign o[2552] = i[4];
  assign o[2553] = i[4];
  assign o[2554] = i[4];
  assign o[2555] = i[4];
  assign o[2556] = i[4];
  assign o[2557] = i[4];
  assign o[2558] = i[4];
  assign o[2559] = i[4];
  assign o[1536] = i[3];
  assign o[1537] = i[3];
  assign o[1538] = i[3];
  assign o[1539] = i[3];
  assign o[1540] = i[3];
  assign o[1541] = i[3];
  assign o[1542] = i[3];
  assign o[1543] = i[3];
  assign o[1544] = i[3];
  assign o[1545] = i[3];
  assign o[1546] = i[3];
  assign o[1547] = i[3];
  assign o[1548] = i[3];
  assign o[1549] = i[3];
  assign o[1550] = i[3];
  assign o[1551] = i[3];
  assign o[1552] = i[3];
  assign o[1553] = i[3];
  assign o[1554] = i[3];
  assign o[1555] = i[3];
  assign o[1556] = i[3];
  assign o[1557] = i[3];
  assign o[1558] = i[3];
  assign o[1559] = i[3];
  assign o[1560] = i[3];
  assign o[1561] = i[3];
  assign o[1562] = i[3];
  assign o[1563] = i[3];
  assign o[1564] = i[3];
  assign o[1565] = i[3];
  assign o[1566] = i[3];
  assign o[1567] = i[3];
  assign o[1568] = i[3];
  assign o[1569] = i[3];
  assign o[1570] = i[3];
  assign o[1571] = i[3];
  assign o[1572] = i[3];
  assign o[1573] = i[3];
  assign o[1574] = i[3];
  assign o[1575] = i[3];
  assign o[1576] = i[3];
  assign o[1577] = i[3];
  assign o[1578] = i[3];
  assign o[1579] = i[3];
  assign o[1580] = i[3];
  assign o[1581] = i[3];
  assign o[1582] = i[3];
  assign o[1583] = i[3];
  assign o[1584] = i[3];
  assign o[1585] = i[3];
  assign o[1586] = i[3];
  assign o[1587] = i[3];
  assign o[1588] = i[3];
  assign o[1589] = i[3];
  assign o[1590] = i[3];
  assign o[1591] = i[3];
  assign o[1592] = i[3];
  assign o[1593] = i[3];
  assign o[1594] = i[3];
  assign o[1595] = i[3];
  assign o[1596] = i[3];
  assign o[1597] = i[3];
  assign o[1598] = i[3];
  assign o[1599] = i[3];
  assign o[1600] = i[3];
  assign o[1601] = i[3];
  assign o[1602] = i[3];
  assign o[1603] = i[3];
  assign o[1604] = i[3];
  assign o[1605] = i[3];
  assign o[1606] = i[3];
  assign o[1607] = i[3];
  assign o[1608] = i[3];
  assign o[1609] = i[3];
  assign o[1610] = i[3];
  assign o[1611] = i[3];
  assign o[1612] = i[3];
  assign o[1613] = i[3];
  assign o[1614] = i[3];
  assign o[1615] = i[3];
  assign o[1616] = i[3];
  assign o[1617] = i[3];
  assign o[1618] = i[3];
  assign o[1619] = i[3];
  assign o[1620] = i[3];
  assign o[1621] = i[3];
  assign o[1622] = i[3];
  assign o[1623] = i[3];
  assign o[1624] = i[3];
  assign o[1625] = i[3];
  assign o[1626] = i[3];
  assign o[1627] = i[3];
  assign o[1628] = i[3];
  assign o[1629] = i[3];
  assign o[1630] = i[3];
  assign o[1631] = i[3];
  assign o[1632] = i[3];
  assign o[1633] = i[3];
  assign o[1634] = i[3];
  assign o[1635] = i[3];
  assign o[1636] = i[3];
  assign o[1637] = i[3];
  assign o[1638] = i[3];
  assign o[1639] = i[3];
  assign o[1640] = i[3];
  assign o[1641] = i[3];
  assign o[1642] = i[3];
  assign o[1643] = i[3];
  assign o[1644] = i[3];
  assign o[1645] = i[3];
  assign o[1646] = i[3];
  assign o[1647] = i[3];
  assign o[1648] = i[3];
  assign o[1649] = i[3];
  assign o[1650] = i[3];
  assign o[1651] = i[3];
  assign o[1652] = i[3];
  assign o[1653] = i[3];
  assign o[1654] = i[3];
  assign o[1655] = i[3];
  assign o[1656] = i[3];
  assign o[1657] = i[3];
  assign o[1658] = i[3];
  assign o[1659] = i[3];
  assign o[1660] = i[3];
  assign o[1661] = i[3];
  assign o[1662] = i[3];
  assign o[1663] = i[3];
  assign o[1664] = i[3];
  assign o[1665] = i[3];
  assign o[1666] = i[3];
  assign o[1667] = i[3];
  assign o[1668] = i[3];
  assign o[1669] = i[3];
  assign o[1670] = i[3];
  assign o[1671] = i[3];
  assign o[1672] = i[3];
  assign o[1673] = i[3];
  assign o[1674] = i[3];
  assign o[1675] = i[3];
  assign o[1676] = i[3];
  assign o[1677] = i[3];
  assign o[1678] = i[3];
  assign o[1679] = i[3];
  assign o[1680] = i[3];
  assign o[1681] = i[3];
  assign o[1682] = i[3];
  assign o[1683] = i[3];
  assign o[1684] = i[3];
  assign o[1685] = i[3];
  assign o[1686] = i[3];
  assign o[1687] = i[3];
  assign o[1688] = i[3];
  assign o[1689] = i[3];
  assign o[1690] = i[3];
  assign o[1691] = i[3];
  assign o[1692] = i[3];
  assign o[1693] = i[3];
  assign o[1694] = i[3];
  assign o[1695] = i[3];
  assign o[1696] = i[3];
  assign o[1697] = i[3];
  assign o[1698] = i[3];
  assign o[1699] = i[3];
  assign o[1700] = i[3];
  assign o[1701] = i[3];
  assign o[1702] = i[3];
  assign o[1703] = i[3];
  assign o[1704] = i[3];
  assign o[1705] = i[3];
  assign o[1706] = i[3];
  assign o[1707] = i[3];
  assign o[1708] = i[3];
  assign o[1709] = i[3];
  assign o[1710] = i[3];
  assign o[1711] = i[3];
  assign o[1712] = i[3];
  assign o[1713] = i[3];
  assign o[1714] = i[3];
  assign o[1715] = i[3];
  assign o[1716] = i[3];
  assign o[1717] = i[3];
  assign o[1718] = i[3];
  assign o[1719] = i[3];
  assign o[1720] = i[3];
  assign o[1721] = i[3];
  assign o[1722] = i[3];
  assign o[1723] = i[3];
  assign o[1724] = i[3];
  assign o[1725] = i[3];
  assign o[1726] = i[3];
  assign o[1727] = i[3];
  assign o[1728] = i[3];
  assign o[1729] = i[3];
  assign o[1730] = i[3];
  assign o[1731] = i[3];
  assign o[1732] = i[3];
  assign o[1733] = i[3];
  assign o[1734] = i[3];
  assign o[1735] = i[3];
  assign o[1736] = i[3];
  assign o[1737] = i[3];
  assign o[1738] = i[3];
  assign o[1739] = i[3];
  assign o[1740] = i[3];
  assign o[1741] = i[3];
  assign o[1742] = i[3];
  assign o[1743] = i[3];
  assign o[1744] = i[3];
  assign o[1745] = i[3];
  assign o[1746] = i[3];
  assign o[1747] = i[3];
  assign o[1748] = i[3];
  assign o[1749] = i[3];
  assign o[1750] = i[3];
  assign o[1751] = i[3];
  assign o[1752] = i[3];
  assign o[1753] = i[3];
  assign o[1754] = i[3];
  assign o[1755] = i[3];
  assign o[1756] = i[3];
  assign o[1757] = i[3];
  assign o[1758] = i[3];
  assign o[1759] = i[3];
  assign o[1760] = i[3];
  assign o[1761] = i[3];
  assign o[1762] = i[3];
  assign o[1763] = i[3];
  assign o[1764] = i[3];
  assign o[1765] = i[3];
  assign o[1766] = i[3];
  assign o[1767] = i[3];
  assign o[1768] = i[3];
  assign o[1769] = i[3];
  assign o[1770] = i[3];
  assign o[1771] = i[3];
  assign o[1772] = i[3];
  assign o[1773] = i[3];
  assign o[1774] = i[3];
  assign o[1775] = i[3];
  assign o[1776] = i[3];
  assign o[1777] = i[3];
  assign o[1778] = i[3];
  assign o[1779] = i[3];
  assign o[1780] = i[3];
  assign o[1781] = i[3];
  assign o[1782] = i[3];
  assign o[1783] = i[3];
  assign o[1784] = i[3];
  assign o[1785] = i[3];
  assign o[1786] = i[3];
  assign o[1787] = i[3];
  assign o[1788] = i[3];
  assign o[1789] = i[3];
  assign o[1790] = i[3];
  assign o[1791] = i[3];
  assign o[1792] = i[3];
  assign o[1793] = i[3];
  assign o[1794] = i[3];
  assign o[1795] = i[3];
  assign o[1796] = i[3];
  assign o[1797] = i[3];
  assign o[1798] = i[3];
  assign o[1799] = i[3];
  assign o[1800] = i[3];
  assign o[1801] = i[3];
  assign o[1802] = i[3];
  assign o[1803] = i[3];
  assign o[1804] = i[3];
  assign o[1805] = i[3];
  assign o[1806] = i[3];
  assign o[1807] = i[3];
  assign o[1808] = i[3];
  assign o[1809] = i[3];
  assign o[1810] = i[3];
  assign o[1811] = i[3];
  assign o[1812] = i[3];
  assign o[1813] = i[3];
  assign o[1814] = i[3];
  assign o[1815] = i[3];
  assign o[1816] = i[3];
  assign o[1817] = i[3];
  assign o[1818] = i[3];
  assign o[1819] = i[3];
  assign o[1820] = i[3];
  assign o[1821] = i[3];
  assign o[1822] = i[3];
  assign o[1823] = i[3];
  assign o[1824] = i[3];
  assign o[1825] = i[3];
  assign o[1826] = i[3];
  assign o[1827] = i[3];
  assign o[1828] = i[3];
  assign o[1829] = i[3];
  assign o[1830] = i[3];
  assign o[1831] = i[3];
  assign o[1832] = i[3];
  assign o[1833] = i[3];
  assign o[1834] = i[3];
  assign o[1835] = i[3];
  assign o[1836] = i[3];
  assign o[1837] = i[3];
  assign o[1838] = i[3];
  assign o[1839] = i[3];
  assign o[1840] = i[3];
  assign o[1841] = i[3];
  assign o[1842] = i[3];
  assign o[1843] = i[3];
  assign o[1844] = i[3];
  assign o[1845] = i[3];
  assign o[1846] = i[3];
  assign o[1847] = i[3];
  assign o[1848] = i[3];
  assign o[1849] = i[3];
  assign o[1850] = i[3];
  assign o[1851] = i[3];
  assign o[1852] = i[3];
  assign o[1853] = i[3];
  assign o[1854] = i[3];
  assign o[1855] = i[3];
  assign o[1856] = i[3];
  assign o[1857] = i[3];
  assign o[1858] = i[3];
  assign o[1859] = i[3];
  assign o[1860] = i[3];
  assign o[1861] = i[3];
  assign o[1862] = i[3];
  assign o[1863] = i[3];
  assign o[1864] = i[3];
  assign o[1865] = i[3];
  assign o[1866] = i[3];
  assign o[1867] = i[3];
  assign o[1868] = i[3];
  assign o[1869] = i[3];
  assign o[1870] = i[3];
  assign o[1871] = i[3];
  assign o[1872] = i[3];
  assign o[1873] = i[3];
  assign o[1874] = i[3];
  assign o[1875] = i[3];
  assign o[1876] = i[3];
  assign o[1877] = i[3];
  assign o[1878] = i[3];
  assign o[1879] = i[3];
  assign o[1880] = i[3];
  assign o[1881] = i[3];
  assign o[1882] = i[3];
  assign o[1883] = i[3];
  assign o[1884] = i[3];
  assign o[1885] = i[3];
  assign o[1886] = i[3];
  assign o[1887] = i[3];
  assign o[1888] = i[3];
  assign o[1889] = i[3];
  assign o[1890] = i[3];
  assign o[1891] = i[3];
  assign o[1892] = i[3];
  assign o[1893] = i[3];
  assign o[1894] = i[3];
  assign o[1895] = i[3];
  assign o[1896] = i[3];
  assign o[1897] = i[3];
  assign o[1898] = i[3];
  assign o[1899] = i[3];
  assign o[1900] = i[3];
  assign o[1901] = i[3];
  assign o[1902] = i[3];
  assign o[1903] = i[3];
  assign o[1904] = i[3];
  assign o[1905] = i[3];
  assign o[1906] = i[3];
  assign o[1907] = i[3];
  assign o[1908] = i[3];
  assign o[1909] = i[3];
  assign o[1910] = i[3];
  assign o[1911] = i[3];
  assign o[1912] = i[3];
  assign o[1913] = i[3];
  assign o[1914] = i[3];
  assign o[1915] = i[3];
  assign o[1916] = i[3];
  assign o[1917] = i[3];
  assign o[1918] = i[3];
  assign o[1919] = i[3];
  assign o[1920] = i[3];
  assign o[1921] = i[3];
  assign o[1922] = i[3];
  assign o[1923] = i[3];
  assign o[1924] = i[3];
  assign o[1925] = i[3];
  assign o[1926] = i[3];
  assign o[1927] = i[3];
  assign o[1928] = i[3];
  assign o[1929] = i[3];
  assign o[1930] = i[3];
  assign o[1931] = i[3];
  assign o[1932] = i[3];
  assign o[1933] = i[3];
  assign o[1934] = i[3];
  assign o[1935] = i[3];
  assign o[1936] = i[3];
  assign o[1937] = i[3];
  assign o[1938] = i[3];
  assign o[1939] = i[3];
  assign o[1940] = i[3];
  assign o[1941] = i[3];
  assign o[1942] = i[3];
  assign o[1943] = i[3];
  assign o[1944] = i[3];
  assign o[1945] = i[3];
  assign o[1946] = i[3];
  assign o[1947] = i[3];
  assign o[1948] = i[3];
  assign o[1949] = i[3];
  assign o[1950] = i[3];
  assign o[1951] = i[3];
  assign o[1952] = i[3];
  assign o[1953] = i[3];
  assign o[1954] = i[3];
  assign o[1955] = i[3];
  assign o[1956] = i[3];
  assign o[1957] = i[3];
  assign o[1958] = i[3];
  assign o[1959] = i[3];
  assign o[1960] = i[3];
  assign o[1961] = i[3];
  assign o[1962] = i[3];
  assign o[1963] = i[3];
  assign o[1964] = i[3];
  assign o[1965] = i[3];
  assign o[1966] = i[3];
  assign o[1967] = i[3];
  assign o[1968] = i[3];
  assign o[1969] = i[3];
  assign o[1970] = i[3];
  assign o[1971] = i[3];
  assign o[1972] = i[3];
  assign o[1973] = i[3];
  assign o[1974] = i[3];
  assign o[1975] = i[3];
  assign o[1976] = i[3];
  assign o[1977] = i[3];
  assign o[1978] = i[3];
  assign o[1979] = i[3];
  assign o[1980] = i[3];
  assign o[1981] = i[3];
  assign o[1982] = i[3];
  assign o[1983] = i[3];
  assign o[1984] = i[3];
  assign o[1985] = i[3];
  assign o[1986] = i[3];
  assign o[1987] = i[3];
  assign o[1988] = i[3];
  assign o[1989] = i[3];
  assign o[1990] = i[3];
  assign o[1991] = i[3];
  assign o[1992] = i[3];
  assign o[1993] = i[3];
  assign o[1994] = i[3];
  assign o[1995] = i[3];
  assign o[1996] = i[3];
  assign o[1997] = i[3];
  assign o[1998] = i[3];
  assign o[1999] = i[3];
  assign o[2000] = i[3];
  assign o[2001] = i[3];
  assign o[2002] = i[3];
  assign o[2003] = i[3];
  assign o[2004] = i[3];
  assign o[2005] = i[3];
  assign o[2006] = i[3];
  assign o[2007] = i[3];
  assign o[2008] = i[3];
  assign o[2009] = i[3];
  assign o[2010] = i[3];
  assign o[2011] = i[3];
  assign o[2012] = i[3];
  assign o[2013] = i[3];
  assign o[2014] = i[3];
  assign o[2015] = i[3];
  assign o[2016] = i[3];
  assign o[2017] = i[3];
  assign o[2018] = i[3];
  assign o[2019] = i[3];
  assign o[2020] = i[3];
  assign o[2021] = i[3];
  assign o[2022] = i[3];
  assign o[2023] = i[3];
  assign o[2024] = i[3];
  assign o[2025] = i[3];
  assign o[2026] = i[3];
  assign o[2027] = i[3];
  assign o[2028] = i[3];
  assign o[2029] = i[3];
  assign o[2030] = i[3];
  assign o[2031] = i[3];
  assign o[2032] = i[3];
  assign o[2033] = i[3];
  assign o[2034] = i[3];
  assign o[2035] = i[3];
  assign o[2036] = i[3];
  assign o[2037] = i[3];
  assign o[2038] = i[3];
  assign o[2039] = i[3];
  assign o[2040] = i[3];
  assign o[2041] = i[3];
  assign o[2042] = i[3];
  assign o[2043] = i[3];
  assign o[2044] = i[3];
  assign o[2045] = i[3];
  assign o[2046] = i[3];
  assign o[2047] = i[3];
  assign o[1024] = i[2];
  assign o[1025] = i[2];
  assign o[1026] = i[2];
  assign o[1027] = i[2];
  assign o[1028] = i[2];
  assign o[1029] = i[2];
  assign o[1030] = i[2];
  assign o[1031] = i[2];
  assign o[1032] = i[2];
  assign o[1033] = i[2];
  assign o[1034] = i[2];
  assign o[1035] = i[2];
  assign o[1036] = i[2];
  assign o[1037] = i[2];
  assign o[1038] = i[2];
  assign o[1039] = i[2];
  assign o[1040] = i[2];
  assign o[1041] = i[2];
  assign o[1042] = i[2];
  assign o[1043] = i[2];
  assign o[1044] = i[2];
  assign o[1045] = i[2];
  assign o[1046] = i[2];
  assign o[1047] = i[2];
  assign o[1048] = i[2];
  assign o[1049] = i[2];
  assign o[1050] = i[2];
  assign o[1051] = i[2];
  assign o[1052] = i[2];
  assign o[1053] = i[2];
  assign o[1054] = i[2];
  assign o[1055] = i[2];
  assign o[1056] = i[2];
  assign o[1057] = i[2];
  assign o[1058] = i[2];
  assign o[1059] = i[2];
  assign o[1060] = i[2];
  assign o[1061] = i[2];
  assign o[1062] = i[2];
  assign o[1063] = i[2];
  assign o[1064] = i[2];
  assign o[1065] = i[2];
  assign o[1066] = i[2];
  assign o[1067] = i[2];
  assign o[1068] = i[2];
  assign o[1069] = i[2];
  assign o[1070] = i[2];
  assign o[1071] = i[2];
  assign o[1072] = i[2];
  assign o[1073] = i[2];
  assign o[1074] = i[2];
  assign o[1075] = i[2];
  assign o[1076] = i[2];
  assign o[1077] = i[2];
  assign o[1078] = i[2];
  assign o[1079] = i[2];
  assign o[1080] = i[2];
  assign o[1081] = i[2];
  assign o[1082] = i[2];
  assign o[1083] = i[2];
  assign o[1084] = i[2];
  assign o[1085] = i[2];
  assign o[1086] = i[2];
  assign o[1087] = i[2];
  assign o[1088] = i[2];
  assign o[1089] = i[2];
  assign o[1090] = i[2];
  assign o[1091] = i[2];
  assign o[1092] = i[2];
  assign o[1093] = i[2];
  assign o[1094] = i[2];
  assign o[1095] = i[2];
  assign o[1096] = i[2];
  assign o[1097] = i[2];
  assign o[1098] = i[2];
  assign o[1099] = i[2];
  assign o[1100] = i[2];
  assign o[1101] = i[2];
  assign o[1102] = i[2];
  assign o[1103] = i[2];
  assign o[1104] = i[2];
  assign o[1105] = i[2];
  assign o[1106] = i[2];
  assign o[1107] = i[2];
  assign o[1108] = i[2];
  assign o[1109] = i[2];
  assign o[1110] = i[2];
  assign o[1111] = i[2];
  assign o[1112] = i[2];
  assign o[1113] = i[2];
  assign o[1114] = i[2];
  assign o[1115] = i[2];
  assign o[1116] = i[2];
  assign o[1117] = i[2];
  assign o[1118] = i[2];
  assign o[1119] = i[2];
  assign o[1120] = i[2];
  assign o[1121] = i[2];
  assign o[1122] = i[2];
  assign o[1123] = i[2];
  assign o[1124] = i[2];
  assign o[1125] = i[2];
  assign o[1126] = i[2];
  assign o[1127] = i[2];
  assign o[1128] = i[2];
  assign o[1129] = i[2];
  assign o[1130] = i[2];
  assign o[1131] = i[2];
  assign o[1132] = i[2];
  assign o[1133] = i[2];
  assign o[1134] = i[2];
  assign o[1135] = i[2];
  assign o[1136] = i[2];
  assign o[1137] = i[2];
  assign o[1138] = i[2];
  assign o[1139] = i[2];
  assign o[1140] = i[2];
  assign o[1141] = i[2];
  assign o[1142] = i[2];
  assign o[1143] = i[2];
  assign o[1144] = i[2];
  assign o[1145] = i[2];
  assign o[1146] = i[2];
  assign o[1147] = i[2];
  assign o[1148] = i[2];
  assign o[1149] = i[2];
  assign o[1150] = i[2];
  assign o[1151] = i[2];
  assign o[1152] = i[2];
  assign o[1153] = i[2];
  assign o[1154] = i[2];
  assign o[1155] = i[2];
  assign o[1156] = i[2];
  assign o[1157] = i[2];
  assign o[1158] = i[2];
  assign o[1159] = i[2];
  assign o[1160] = i[2];
  assign o[1161] = i[2];
  assign o[1162] = i[2];
  assign o[1163] = i[2];
  assign o[1164] = i[2];
  assign o[1165] = i[2];
  assign o[1166] = i[2];
  assign o[1167] = i[2];
  assign o[1168] = i[2];
  assign o[1169] = i[2];
  assign o[1170] = i[2];
  assign o[1171] = i[2];
  assign o[1172] = i[2];
  assign o[1173] = i[2];
  assign o[1174] = i[2];
  assign o[1175] = i[2];
  assign o[1176] = i[2];
  assign o[1177] = i[2];
  assign o[1178] = i[2];
  assign o[1179] = i[2];
  assign o[1180] = i[2];
  assign o[1181] = i[2];
  assign o[1182] = i[2];
  assign o[1183] = i[2];
  assign o[1184] = i[2];
  assign o[1185] = i[2];
  assign o[1186] = i[2];
  assign o[1187] = i[2];
  assign o[1188] = i[2];
  assign o[1189] = i[2];
  assign o[1190] = i[2];
  assign o[1191] = i[2];
  assign o[1192] = i[2];
  assign o[1193] = i[2];
  assign o[1194] = i[2];
  assign o[1195] = i[2];
  assign o[1196] = i[2];
  assign o[1197] = i[2];
  assign o[1198] = i[2];
  assign o[1199] = i[2];
  assign o[1200] = i[2];
  assign o[1201] = i[2];
  assign o[1202] = i[2];
  assign o[1203] = i[2];
  assign o[1204] = i[2];
  assign o[1205] = i[2];
  assign o[1206] = i[2];
  assign o[1207] = i[2];
  assign o[1208] = i[2];
  assign o[1209] = i[2];
  assign o[1210] = i[2];
  assign o[1211] = i[2];
  assign o[1212] = i[2];
  assign o[1213] = i[2];
  assign o[1214] = i[2];
  assign o[1215] = i[2];
  assign o[1216] = i[2];
  assign o[1217] = i[2];
  assign o[1218] = i[2];
  assign o[1219] = i[2];
  assign o[1220] = i[2];
  assign o[1221] = i[2];
  assign o[1222] = i[2];
  assign o[1223] = i[2];
  assign o[1224] = i[2];
  assign o[1225] = i[2];
  assign o[1226] = i[2];
  assign o[1227] = i[2];
  assign o[1228] = i[2];
  assign o[1229] = i[2];
  assign o[1230] = i[2];
  assign o[1231] = i[2];
  assign o[1232] = i[2];
  assign o[1233] = i[2];
  assign o[1234] = i[2];
  assign o[1235] = i[2];
  assign o[1236] = i[2];
  assign o[1237] = i[2];
  assign o[1238] = i[2];
  assign o[1239] = i[2];
  assign o[1240] = i[2];
  assign o[1241] = i[2];
  assign o[1242] = i[2];
  assign o[1243] = i[2];
  assign o[1244] = i[2];
  assign o[1245] = i[2];
  assign o[1246] = i[2];
  assign o[1247] = i[2];
  assign o[1248] = i[2];
  assign o[1249] = i[2];
  assign o[1250] = i[2];
  assign o[1251] = i[2];
  assign o[1252] = i[2];
  assign o[1253] = i[2];
  assign o[1254] = i[2];
  assign o[1255] = i[2];
  assign o[1256] = i[2];
  assign o[1257] = i[2];
  assign o[1258] = i[2];
  assign o[1259] = i[2];
  assign o[1260] = i[2];
  assign o[1261] = i[2];
  assign o[1262] = i[2];
  assign o[1263] = i[2];
  assign o[1264] = i[2];
  assign o[1265] = i[2];
  assign o[1266] = i[2];
  assign o[1267] = i[2];
  assign o[1268] = i[2];
  assign o[1269] = i[2];
  assign o[1270] = i[2];
  assign o[1271] = i[2];
  assign o[1272] = i[2];
  assign o[1273] = i[2];
  assign o[1274] = i[2];
  assign o[1275] = i[2];
  assign o[1276] = i[2];
  assign o[1277] = i[2];
  assign o[1278] = i[2];
  assign o[1279] = i[2];
  assign o[1280] = i[2];
  assign o[1281] = i[2];
  assign o[1282] = i[2];
  assign o[1283] = i[2];
  assign o[1284] = i[2];
  assign o[1285] = i[2];
  assign o[1286] = i[2];
  assign o[1287] = i[2];
  assign o[1288] = i[2];
  assign o[1289] = i[2];
  assign o[1290] = i[2];
  assign o[1291] = i[2];
  assign o[1292] = i[2];
  assign o[1293] = i[2];
  assign o[1294] = i[2];
  assign o[1295] = i[2];
  assign o[1296] = i[2];
  assign o[1297] = i[2];
  assign o[1298] = i[2];
  assign o[1299] = i[2];
  assign o[1300] = i[2];
  assign o[1301] = i[2];
  assign o[1302] = i[2];
  assign o[1303] = i[2];
  assign o[1304] = i[2];
  assign o[1305] = i[2];
  assign o[1306] = i[2];
  assign o[1307] = i[2];
  assign o[1308] = i[2];
  assign o[1309] = i[2];
  assign o[1310] = i[2];
  assign o[1311] = i[2];
  assign o[1312] = i[2];
  assign o[1313] = i[2];
  assign o[1314] = i[2];
  assign o[1315] = i[2];
  assign o[1316] = i[2];
  assign o[1317] = i[2];
  assign o[1318] = i[2];
  assign o[1319] = i[2];
  assign o[1320] = i[2];
  assign o[1321] = i[2];
  assign o[1322] = i[2];
  assign o[1323] = i[2];
  assign o[1324] = i[2];
  assign o[1325] = i[2];
  assign o[1326] = i[2];
  assign o[1327] = i[2];
  assign o[1328] = i[2];
  assign o[1329] = i[2];
  assign o[1330] = i[2];
  assign o[1331] = i[2];
  assign o[1332] = i[2];
  assign o[1333] = i[2];
  assign o[1334] = i[2];
  assign o[1335] = i[2];
  assign o[1336] = i[2];
  assign o[1337] = i[2];
  assign o[1338] = i[2];
  assign o[1339] = i[2];
  assign o[1340] = i[2];
  assign o[1341] = i[2];
  assign o[1342] = i[2];
  assign o[1343] = i[2];
  assign o[1344] = i[2];
  assign o[1345] = i[2];
  assign o[1346] = i[2];
  assign o[1347] = i[2];
  assign o[1348] = i[2];
  assign o[1349] = i[2];
  assign o[1350] = i[2];
  assign o[1351] = i[2];
  assign o[1352] = i[2];
  assign o[1353] = i[2];
  assign o[1354] = i[2];
  assign o[1355] = i[2];
  assign o[1356] = i[2];
  assign o[1357] = i[2];
  assign o[1358] = i[2];
  assign o[1359] = i[2];
  assign o[1360] = i[2];
  assign o[1361] = i[2];
  assign o[1362] = i[2];
  assign o[1363] = i[2];
  assign o[1364] = i[2];
  assign o[1365] = i[2];
  assign o[1366] = i[2];
  assign o[1367] = i[2];
  assign o[1368] = i[2];
  assign o[1369] = i[2];
  assign o[1370] = i[2];
  assign o[1371] = i[2];
  assign o[1372] = i[2];
  assign o[1373] = i[2];
  assign o[1374] = i[2];
  assign o[1375] = i[2];
  assign o[1376] = i[2];
  assign o[1377] = i[2];
  assign o[1378] = i[2];
  assign o[1379] = i[2];
  assign o[1380] = i[2];
  assign o[1381] = i[2];
  assign o[1382] = i[2];
  assign o[1383] = i[2];
  assign o[1384] = i[2];
  assign o[1385] = i[2];
  assign o[1386] = i[2];
  assign o[1387] = i[2];
  assign o[1388] = i[2];
  assign o[1389] = i[2];
  assign o[1390] = i[2];
  assign o[1391] = i[2];
  assign o[1392] = i[2];
  assign o[1393] = i[2];
  assign o[1394] = i[2];
  assign o[1395] = i[2];
  assign o[1396] = i[2];
  assign o[1397] = i[2];
  assign o[1398] = i[2];
  assign o[1399] = i[2];
  assign o[1400] = i[2];
  assign o[1401] = i[2];
  assign o[1402] = i[2];
  assign o[1403] = i[2];
  assign o[1404] = i[2];
  assign o[1405] = i[2];
  assign o[1406] = i[2];
  assign o[1407] = i[2];
  assign o[1408] = i[2];
  assign o[1409] = i[2];
  assign o[1410] = i[2];
  assign o[1411] = i[2];
  assign o[1412] = i[2];
  assign o[1413] = i[2];
  assign o[1414] = i[2];
  assign o[1415] = i[2];
  assign o[1416] = i[2];
  assign o[1417] = i[2];
  assign o[1418] = i[2];
  assign o[1419] = i[2];
  assign o[1420] = i[2];
  assign o[1421] = i[2];
  assign o[1422] = i[2];
  assign o[1423] = i[2];
  assign o[1424] = i[2];
  assign o[1425] = i[2];
  assign o[1426] = i[2];
  assign o[1427] = i[2];
  assign o[1428] = i[2];
  assign o[1429] = i[2];
  assign o[1430] = i[2];
  assign o[1431] = i[2];
  assign o[1432] = i[2];
  assign o[1433] = i[2];
  assign o[1434] = i[2];
  assign o[1435] = i[2];
  assign o[1436] = i[2];
  assign o[1437] = i[2];
  assign o[1438] = i[2];
  assign o[1439] = i[2];
  assign o[1440] = i[2];
  assign o[1441] = i[2];
  assign o[1442] = i[2];
  assign o[1443] = i[2];
  assign o[1444] = i[2];
  assign o[1445] = i[2];
  assign o[1446] = i[2];
  assign o[1447] = i[2];
  assign o[1448] = i[2];
  assign o[1449] = i[2];
  assign o[1450] = i[2];
  assign o[1451] = i[2];
  assign o[1452] = i[2];
  assign o[1453] = i[2];
  assign o[1454] = i[2];
  assign o[1455] = i[2];
  assign o[1456] = i[2];
  assign o[1457] = i[2];
  assign o[1458] = i[2];
  assign o[1459] = i[2];
  assign o[1460] = i[2];
  assign o[1461] = i[2];
  assign o[1462] = i[2];
  assign o[1463] = i[2];
  assign o[1464] = i[2];
  assign o[1465] = i[2];
  assign o[1466] = i[2];
  assign o[1467] = i[2];
  assign o[1468] = i[2];
  assign o[1469] = i[2];
  assign o[1470] = i[2];
  assign o[1471] = i[2];
  assign o[1472] = i[2];
  assign o[1473] = i[2];
  assign o[1474] = i[2];
  assign o[1475] = i[2];
  assign o[1476] = i[2];
  assign o[1477] = i[2];
  assign o[1478] = i[2];
  assign o[1479] = i[2];
  assign o[1480] = i[2];
  assign o[1481] = i[2];
  assign o[1482] = i[2];
  assign o[1483] = i[2];
  assign o[1484] = i[2];
  assign o[1485] = i[2];
  assign o[1486] = i[2];
  assign o[1487] = i[2];
  assign o[1488] = i[2];
  assign o[1489] = i[2];
  assign o[1490] = i[2];
  assign o[1491] = i[2];
  assign o[1492] = i[2];
  assign o[1493] = i[2];
  assign o[1494] = i[2];
  assign o[1495] = i[2];
  assign o[1496] = i[2];
  assign o[1497] = i[2];
  assign o[1498] = i[2];
  assign o[1499] = i[2];
  assign o[1500] = i[2];
  assign o[1501] = i[2];
  assign o[1502] = i[2];
  assign o[1503] = i[2];
  assign o[1504] = i[2];
  assign o[1505] = i[2];
  assign o[1506] = i[2];
  assign o[1507] = i[2];
  assign o[1508] = i[2];
  assign o[1509] = i[2];
  assign o[1510] = i[2];
  assign o[1511] = i[2];
  assign o[1512] = i[2];
  assign o[1513] = i[2];
  assign o[1514] = i[2];
  assign o[1515] = i[2];
  assign o[1516] = i[2];
  assign o[1517] = i[2];
  assign o[1518] = i[2];
  assign o[1519] = i[2];
  assign o[1520] = i[2];
  assign o[1521] = i[2];
  assign o[1522] = i[2];
  assign o[1523] = i[2];
  assign o[1524] = i[2];
  assign o[1525] = i[2];
  assign o[1526] = i[2];
  assign o[1527] = i[2];
  assign o[1528] = i[2];
  assign o[1529] = i[2];
  assign o[1530] = i[2];
  assign o[1531] = i[2];
  assign o[1532] = i[2];
  assign o[1533] = i[2];
  assign o[1534] = i[2];
  assign o[1535] = i[2];
  assign o[512] = i[1];
  assign o[513] = i[1];
  assign o[514] = i[1];
  assign o[515] = i[1];
  assign o[516] = i[1];
  assign o[517] = i[1];
  assign o[518] = i[1];
  assign o[519] = i[1];
  assign o[520] = i[1];
  assign o[521] = i[1];
  assign o[522] = i[1];
  assign o[523] = i[1];
  assign o[524] = i[1];
  assign o[525] = i[1];
  assign o[526] = i[1];
  assign o[527] = i[1];
  assign o[528] = i[1];
  assign o[529] = i[1];
  assign o[530] = i[1];
  assign o[531] = i[1];
  assign o[532] = i[1];
  assign o[533] = i[1];
  assign o[534] = i[1];
  assign o[535] = i[1];
  assign o[536] = i[1];
  assign o[537] = i[1];
  assign o[538] = i[1];
  assign o[539] = i[1];
  assign o[540] = i[1];
  assign o[541] = i[1];
  assign o[542] = i[1];
  assign o[543] = i[1];
  assign o[544] = i[1];
  assign o[545] = i[1];
  assign o[546] = i[1];
  assign o[547] = i[1];
  assign o[548] = i[1];
  assign o[549] = i[1];
  assign o[550] = i[1];
  assign o[551] = i[1];
  assign o[552] = i[1];
  assign o[553] = i[1];
  assign o[554] = i[1];
  assign o[555] = i[1];
  assign o[556] = i[1];
  assign o[557] = i[1];
  assign o[558] = i[1];
  assign o[559] = i[1];
  assign o[560] = i[1];
  assign o[561] = i[1];
  assign o[562] = i[1];
  assign o[563] = i[1];
  assign o[564] = i[1];
  assign o[565] = i[1];
  assign o[566] = i[1];
  assign o[567] = i[1];
  assign o[568] = i[1];
  assign o[569] = i[1];
  assign o[570] = i[1];
  assign o[571] = i[1];
  assign o[572] = i[1];
  assign o[573] = i[1];
  assign o[574] = i[1];
  assign o[575] = i[1];
  assign o[576] = i[1];
  assign o[577] = i[1];
  assign o[578] = i[1];
  assign o[579] = i[1];
  assign o[580] = i[1];
  assign o[581] = i[1];
  assign o[582] = i[1];
  assign o[583] = i[1];
  assign o[584] = i[1];
  assign o[585] = i[1];
  assign o[586] = i[1];
  assign o[587] = i[1];
  assign o[588] = i[1];
  assign o[589] = i[1];
  assign o[590] = i[1];
  assign o[591] = i[1];
  assign o[592] = i[1];
  assign o[593] = i[1];
  assign o[594] = i[1];
  assign o[595] = i[1];
  assign o[596] = i[1];
  assign o[597] = i[1];
  assign o[598] = i[1];
  assign o[599] = i[1];
  assign o[600] = i[1];
  assign o[601] = i[1];
  assign o[602] = i[1];
  assign o[603] = i[1];
  assign o[604] = i[1];
  assign o[605] = i[1];
  assign o[606] = i[1];
  assign o[607] = i[1];
  assign o[608] = i[1];
  assign o[609] = i[1];
  assign o[610] = i[1];
  assign o[611] = i[1];
  assign o[612] = i[1];
  assign o[613] = i[1];
  assign o[614] = i[1];
  assign o[615] = i[1];
  assign o[616] = i[1];
  assign o[617] = i[1];
  assign o[618] = i[1];
  assign o[619] = i[1];
  assign o[620] = i[1];
  assign o[621] = i[1];
  assign o[622] = i[1];
  assign o[623] = i[1];
  assign o[624] = i[1];
  assign o[625] = i[1];
  assign o[626] = i[1];
  assign o[627] = i[1];
  assign o[628] = i[1];
  assign o[629] = i[1];
  assign o[630] = i[1];
  assign o[631] = i[1];
  assign o[632] = i[1];
  assign o[633] = i[1];
  assign o[634] = i[1];
  assign o[635] = i[1];
  assign o[636] = i[1];
  assign o[637] = i[1];
  assign o[638] = i[1];
  assign o[639] = i[1];
  assign o[640] = i[1];
  assign o[641] = i[1];
  assign o[642] = i[1];
  assign o[643] = i[1];
  assign o[644] = i[1];
  assign o[645] = i[1];
  assign o[646] = i[1];
  assign o[647] = i[1];
  assign o[648] = i[1];
  assign o[649] = i[1];
  assign o[650] = i[1];
  assign o[651] = i[1];
  assign o[652] = i[1];
  assign o[653] = i[1];
  assign o[654] = i[1];
  assign o[655] = i[1];
  assign o[656] = i[1];
  assign o[657] = i[1];
  assign o[658] = i[1];
  assign o[659] = i[1];
  assign o[660] = i[1];
  assign o[661] = i[1];
  assign o[662] = i[1];
  assign o[663] = i[1];
  assign o[664] = i[1];
  assign o[665] = i[1];
  assign o[666] = i[1];
  assign o[667] = i[1];
  assign o[668] = i[1];
  assign o[669] = i[1];
  assign o[670] = i[1];
  assign o[671] = i[1];
  assign o[672] = i[1];
  assign o[673] = i[1];
  assign o[674] = i[1];
  assign o[675] = i[1];
  assign o[676] = i[1];
  assign o[677] = i[1];
  assign o[678] = i[1];
  assign o[679] = i[1];
  assign o[680] = i[1];
  assign o[681] = i[1];
  assign o[682] = i[1];
  assign o[683] = i[1];
  assign o[684] = i[1];
  assign o[685] = i[1];
  assign o[686] = i[1];
  assign o[687] = i[1];
  assign o[688] = i[1];
  assign o[689] = i[1];
  assign o[690] = i[1];
  assign o[691] = i[1];
  assign o[692] = i[1];
  assign o[693] = i[1];
  assign o[694] = i[1];
  assign o[695] = i[1];
  assign o[696] = i[1];
  assign o[697] = i[1];
  assign o[698] = i[1];
  assign o[699] = i[1];
  assign o[700] = i[1];
  assign o[701] = i[1];
  assign o[702] = i[1];
  assign o[703] = i[1];
  assign o[704] = i[1];
  assign o[705] = i[1];
  assign o[706] = i[1];
  assign o[707] = i[1];
  assign o[708] = i[1];
  assign o[709] = i[1];
  assign o[710] = i[1];
  assign o[711] = i[1];
  assign o[712] = i[1];
  assign o[713] = i[1];
  assign o[714] = i[1];
  assign o[715] = i[1];
  assign o[716] = i[1];
  assign o[717] = i[1];
  assign o[718] = i[1];
  assign o[719] = i[1];
  assign o[720] = i[1];
  assign o[721] = i[1];
  assign o[722] = i[1];
  assign o[723] = i[1];
  assign o[724] = i[1];
  assign o[725] = i[1];
  assign o[726] = i[1];
  assign o[727] = i[1];
  assign o[728] = i[1];
  assign o[729] = i[1];
  assign o[730] = i[1];
  assign o[731] = i[1];
  assign o[732] = i[1];
  assign o[733] = i[1];
  assign o[734] = i[1];
  assign o[735] = i[1];
  assign o[736] = i[1];
  assign o[737] = i[1];
  assign o[738] = i[1];
  assign o[739] = i[1];
  assign o[740] = i[1];
  assign o[741] = i[1];
  assign o[742] = i[1];
  assign o[743] = i[1];
  assign o[744] = i[1];
  assign o[745] = i[1];
  assign o[746] = i[1];
  assign o[747] = i[1];
  assign o[748] = i[1];
  assign o[749] = i[1];
  assign o[750] = i[1];
  assign o[751] = i[1];
  assign o[752] = i[1];
  assign o[753] = i[1];
  assign o[754] = i[1];
  assign o[755] = i[1];
  assign o[756] = i[1];
  assign o[757] = i[1];
  assign o[758] = i[1];
  assign o[759] = i[1];
  assign o[760] = i[1];
  assign o[761] = i[1];
  assign o[762] = i[1];
  assign o[763] = i[1];
  assign o[764] = i[1];
  assign o[765] = i[1];
  assign o[766] = i[1];
  assign o[767] = i[1];
  assign o[768] = i[1];
  assign o[769] = i[1];
  assign o[770] = i[1];
  assign o[771] = i[1];
  assign o[772] = i[1];
  assign o[773] = i[1];
  assign o[774] = i[1];
  assign o[775] = i[1];
  assign o[776] = i[1];
  assign o[777] = i[1];
  assign o[778] = i[1];
  assign o[779] = i[1];
  assign o[780] = i[1];
  assign o[781] = i[1];
  assign o[782] = i[1];
  assign o[783] = i[1];
  assign o[784] = i[1];
  assign o[785] = i[1];
  assign o[786] = i[1];
  assign o[787] = i[1];
  assign o[788] = i[1];
  assign o[789] = i[1];
  assign o[790] = i[1];
  assign o[791] = i[1];
  assign o[792] = i[1];
  assign o[793] = i[1];
  assign o[794] = i[1];
  assign o[795] = i[1];
  assign o[796] = i[1];
  assign o[797] = i[1];
  assign o[798] = i[1];
  assign o[799] = i[1];
  assign o[800] = i[1];
  assign o[801] = i[1];
  assign o[802] = i[1];
  assign o[803] = i[1];
  assign o[804] = i[1];
  assign o[805] = i[1];
  assign o[806] = i[1];
  assign o[807] = i[1];
  assign o[808] = i[1];
  assign o[809] = i[1];
  assign o[810] = i[1];
  assign o[811] = i[1];
  assign o[812] = i[1];
  assign o[813] = i[1];
  assign o[814] = i[1];
  assign o[815] = i[1];
  assign o[816] = i[1];
  assign o[817] = i[1];
  assign o[818] = i[1];
  assign o[819] = i[1];
  assign o[820] = i[1];
  assign o[821] = i[1];
  assign o[822] = i[1];
  assign o[823] = i[1];
  assign o[824] = i[1];
  assign o[825] = i[1];
  assign o[826] = i[1];
  assign o[827] = i[1];
  assign o[828] = i[1];
  assign o[829] = i[1];
  assign o[830] = i[1];
  assign o[831] = i[1];
  assign o[832] = i[1];
  assign o[833] = i[1];
  assign o[834] = i[1];
  assign o[835] = i[1];
  assign o[836] = i[1];
  assign o[837] = i[1];
  assign o[838] = i[1];
  assign o[839] = i[1];
  assign o[840] = i[1];
  assign o[841] = i[1];
  assign o[842] = i[1];
  assign o[843] = i[1];
  assign o[844] = i[1];
  assign o[845] = i[1];
  assign o[846] = i[1];
  assign o[847] = i[1];
  assign o[848] = i[1];
  assign o[849] = i[1];
  assign o[850] = i[1];
  assign o[851] = i[1];
  assign o[852] = i[1];
  assign o[853] = i[1];
  assign o[854] = i[1];
  assign o[855] = i[1];
  assign o[856] = i[1];
  assign o[857] = i[1];
  assign o[858] = i[1];
  assign o[859] = i[1];
  assign o[860] = i[1];
  assign o[861] = i[1];
  assign o[862] = i[1];
  assign o[863] = i[1];
  assign o[864] = i[1];
  assign o[865] = i[1];
  assign o[866] = i[1];
  assign o[867] = i[1];
  assign o[868] = i[1];
  assign o[869] = i[1];
  assign o[870] = i[1];
  assign o[871] = i[1];
  assign o[872] = i[1];
  assign o[873] = i[1];
  assign o[874] = i[1];
  assign o[875] = i[1];
  assign o[876] = i[1];
  assign o[877] = i[1];
  assign o[878] = i[1];
  assign o[879] = i[1];
  assign o[880] = i[1];
  assign o[881] = i[1];
  assign o[882] = i[1];
  assign o[883] = i[1];
  assign o[884] = i[1];
  assign o[885] = i[1];
  assign o[886] = i[1];
  assign o[887] = i[1];
  assign o[888] = i[1];
  assign o[889] = i[1];
  assign o[890] = i[1];
  assign o[891] = i[1];
  assign o[892] = i[1];
  assign o[893] = i[1];
  assign o[894] = i[1];
  assign o[895] = i[1];
  assign o[896] = i[1];
  assign o[897] = i[1];
  assign o[898] = i[1];
  assign o[899] = i[1];
  assign o[900] = i[1];
  assign o[901] = i[1];
  assign o[902] = i[1];
  assign o[903] = i[1];
  assign o[904] = i[1];
  assign o[905] = i[1];
  assign o[906] = i[1];
  assign o[907] = i[1];
  assign o[908] = i[1];
  assign o[909] = i[1];
  assign o[910] = i[1];
  assign o[911] = i[1];
  assign o[912] = i[1];
  assign o[913] = i[1];
  assign o[914] = i[1];
  assign o[915] = i[1];
  assign o[916] = i[1];
  assign o[917] = i[1];
  assign o[918] = i[1];
  assign o[919] = i[1];
  assign o[920] = i[1];
  assign o[921] = i[1];
  assign o[922] = i[1];
  assign o[923] = i[1];
  assign o[924] = i[1];
  assign o[925] = i[1];
  assign o[926] = i[1];
  assign o[927] = i[1];
  assign o[928] = i[1];
  assign o[929] = i[1];
  assign o[930] = i[1];
  assign o[931] = i[1];
  assign o[932] = i[1];
  assign o[933] = i[1];
  assign o[934] = i[1];
  assign o[935] = i[1];
  assign o[936] = i[1];
  assign o[937] = i[1];
  assign o[938] = i[1];
  assign o[939] = i[1];
  assign o[940] = i[1];
  assign o[941] = i[1];
  assign o[942] = i[1];
  assign o[943] = i[1];
  assign o[944] = i[1];
  assign o[945] = i[1];
  assign o[946] = i[1];
  assign o[947] = i[1];
  assign o[948] = i[1];
  assign o[949] = i[1];
  assign o[950] = i[1];
  assign o[951] = i[1];
  assign o[952] = i[1];
  assign o[953] = i[1];
  assign o[954] = i[1];
  assign o[955] = i[1];
  assign o[956] = i[1];
  assign o[957] = i[1];
  assign o[958] = i[1];
  assign o[959] = i[1];
  assign o[960] = i[1];
  assign o[961] = i[1];
  assign o[962] = i[1];
  assign o[963] = i[1];
  assign o[964] = i[1];
  assign o[965] = i[1];
  assign o[966] = i[1];
  assign o[967] = i[1];
  assign o[968] = i[1];
  assign o[969] = i[1];
  assign o[970] = i[1];
  assign o[971] = i[1];
  assign o[972] = i[1];
  assign o[973] = i[1];
  assign o[974] = i[1];
  assign o[975] = i[1];
  assign o[976] = i[1];
  assign o[977] = i[1];
  assign o[978] = i[1];
  assign o[979] = i[1];
  assign o[980] = i[1];
  assign o[981] = i[1];
  assign o[982] = i[1];
  assign o[983] = i[1];
  assign o[984] = i[1];
  assign o[985] = i[1];
  assign o[986] = i[1];
  assign o[987] = i[1];
  assign o[988] = i[1];
  assign o[989] = i[1];
  assign o[990] = i[1];
  assign o[991] = i[1];
  assign o[992] = i[1];
  assign o[993] = i[1];
  assign o[994] = i[1];
  assign o[995] = i[1];
  assign o[996] = i[1];
  assign o[997] = i[1];
  assign o[998] = i[1];
  assign o[999] = i[1];
  assign o[1000] = i[1];
  assign o[1001] = i[1];
  assign o[1002] = i[1];
  assign o[1003] = i[1];
  assign o[1004] = i[1];
  assign o[1005] = i[1];
  assign o[1006] = i[1];
  assign o[1007] = i[1];
  assign o[1008] = i[1];
  assign o[1009] = i[1];
  assign o[1010] = i[1];
  assign o[1011] = i[1];
  assign o[1012] = i[1];
  assign o[1013] = i[1];
  assign o[1014] = i[1];
  assign o[1015] = i[1];
  assign o[1016] = i[1];
  assign o[1017] = i[1];
  assign o[1018] = i[1];
  assign o[1019] = i[1];
  assign o[1020] = i[1];
  assign o[1021] = i[1];
  assign o[1022] = i[1];
  assign o[1023] = i[1];
  assign o[0] = i[0];
  assign o[1] = i[0];
  assign o[2] = i[0];
  assign o[3] = i[0];
  assign o[4] = i[0];
  assign o[5] = i[0];
  assign o[6] = i[0];
  assign o[7] = i[0];
  assign o[8] = i[0];
  assign o[9] = i[0];
  assign o[10] = i[0];
  assign o[11] = i[0];
  assign o[12] = i[0];
  assign o[13] = i[0];
  assign o[14] = i[0];
  assign o[15] = i[0];
  assign o[16] = i[0];
  assign o[17] = i[0];
  assign o[18] = i[0];
  assign o[19] = i[0];
  assign o[20] = i[0];
  assign o[21] = i[0];
  assign o[22] = i[0];
  assign o[23] = i[0];
  assign o[24] = i[0];
  assign o[25] = i[0];
  assign o[26] = i[0];
  assign o[27] = i[0];
  assign o[28] = i[0];
  assign o[29] = i[0];
  assign o[30] = i[0];
  assign o[31] = i[0];
  assign o[32] = i[0];
  assign o[33] = i[0];
  assign o[34] = i[0];
  assign o[35] = i[0];
  assign o[36] = i[0];
  assign o[37] = i[0];
  assign o[38] = i[0];
  assign o[39] = i[0];
  assign o[40] = i[0];
  assign o[41] = i[0];
  assign o[42] = i[0];
  assign o[43] = i[0];
  assign o[44] = i[0];
  assign o[45] = i[0];
  assign o[46] = i[0];
  assign o[47] = i[0];
  assign o[48] = i[0];
  assign o[49] = i[0];
  assign o[50] = i[0];
  assign o[51] = i[0];
  assign o[52] = i[0];
  assign o[53] = i[0];
  assign o[54] = i[0];
  assign o[55] = i[0];
  assign o[56] = i[0];
  assign o[57] = i[0];
  assign o[58] = i[0];
  assign o[59] = i[0];
  assign o[60] = i[0];
  assign o[61] = i[0];
  assign o[62] = i[0];
  assign o[63] = i[0];
  assign o[64] = i[0];
  assign o[65] = i[0];
  assign o[66] = i[0];
  assign o[67] = i[0];
  assign o[68] = i[0];
  assign o[69] = i[0];
  assign o[70] = i[0];
  assign o[71] = i[0];
  assign o[72] = i[0];
  assign o[73] = i[0];
  assign o[74] = i[0];
  assign o[75] = i[0];
  assign o[76] = i[0];
  assign o[77] = i[0];
  assign o[78] = i[0];
  assign o[79] = i[0];
  assign o[80] = i[0];
  assign o[81] = i[0];
  assign o[82] = i[0];
  assign o[83] = i[0];
  assign o[84] = i[0];
  assign o[85] = i[0];
  assign o[86] = i[0];
  assign o[87] = i[0];
  assign o[88] = i[0];
  assign o[89] = i[0];
  assign o[90] = i[0];
  assign o[91] = i[0];
  assign o[92] = i[0];
  assign o[93] = i[0];
  assign o[94] = i[0];
  assign o[95] = i[0];
  assign o[96] = i[0];
  assign o[97] = i[0];
  assign o[98] = i[0];
  assign o[99] = i[0];
  assign o[100] = i[0];
  assign o[101] = i[0];
  assign o[102] = i[0];
  assign o[103] = i[0];
  assign o[104] = i[0];
  assign o[105] = i[0];
  assign o[106] = i[0];
  assign o[107] = i[0];
  assign o[108] = i[0];
  assign o[109] = i[0];
  assign o[110] = i[0];
  assign o[111] = i[0];
  assign o[112] = i[0];
  assign o[113] = i[0];
  assign o[114] = i[0];
  assign o[115] = i[0];
  assign o[116] = i[0];
  assign o[117] = i[0];
  assign o[118] = i[0];
  assign o[119] = i[0];
  assign o[120] = i[0];
  assign o[121] = i[0];
  assign o[122] = i[0];
  assign o[123] = i[0];
  assign o[124] = i[0];
  assign o[125] = i[0];
  assign o[126] = i[0];
  assign o[127] = i[0];
  assign o[128] = i[0];
  assign o[129] = i[0];
  assign o[130] = i[0];
  assign o[131] = i[0];
  assign o[132] = i[0];
  assign o[133] = i[0];
  assign o[134] = i[0];
  assign o[135] = i[0];
  assign o[136] = i[0];
  assign o[137] = i[0];
  assign o[138] = i[0];
  assign o[139] = i[0];
  assign o[140] = i[0];
  assign o[141] = i[0];
  assign o[142] = i[0];
  assign o[143] = i[0];
  assign o[144] = i[0];
  assign o[145] = i[0];
  assign o[146] = i[0];
  assign o[147] = i[0];
  assign o[148] = i[0];
  assign o[149] = i[0];
  assign o[150] = i[0];
  assign o[151] = i[0];
  assign o[152] = i[0];
  assign o[153] = i[0];
  assign o[154] = i[0];
  assign o[155] = i[0];
  assign o[156] = i[0];
  assign o[157] = i[0];
  assign o[158] = i[0];
  assign o[159] = i[0];
  assign o[160] = i[0];
  assign o[161] = i[0];
  assign o[162] = i[0];
  assign o[163] = i[0];
  assign o[164] = i[0];
  assign o[165] = i[0];
  assign o[166] = i[0];
  assign o[167] = i[0];
  assign o[168] = i[0];
  assign o[169] = i[0];
  assign o[170] = i[0];
  assign o[171] = i[0];
  assign o[172] = i[0];
  assign o[173] = i[0];
  assign o[174] = i[0];
  assign o[175] = i[0];
  assign o[176] = i[0];
  assign o[177] = i[0];
  assign o[178] = i[0];
  assign o[179] = i[0];
  assign o[180] = i[0];
  assign o[181] = i[0];
  assign o[182] = i[0];
  assign o[183] = i[0];
  assign o[184] = i[0];
  assign o[185] = i[0];
  assign o[186] = i[0];
  assign o[187] = i[0];
  assign o[188] = i[0];
  assign o[189] = i[0];
  assign o[190] = i[0];
  assign o[191] = i[0];
  assign o[192] = i[0];
  assign o[193] = i[0];
  assign o[194] = i[0];
  assign o[195] = i[0];
  assign o[196] = i[0];
  assign o[197] = i[0];
  assign o[198] = i[0];
  assign o[199] = i[0];
  assign o[200] = i[0];
  assign o[201] = i[0];
  assign o[202] = i[0];
  assign o[203] = i[0];
  assign o[204] = i[0];
  assign o[205] = i[0];
  assign o[206] = i[0];
  assign o[207] = i[0];
  assign o[208] = i[0];
  assign o[209] = i[0];
  assign o[210] = i[0];
  assign o[211] = i[0];
  assign o[212] = i[0];
  assign o[213] = i[0];
  assign o[214] = i[0];
  assign o[215] = i[0];
  assign o[216] = i[0];
  assign o[217] = i[0];
  assign o[218] = i[0];
  assign o[219] = i[0];
  assign o[220] = i[0];
  assign o[221] = i[0];
  assign o[222] = i[0];
  assign o[223] = i[0];
  assign o[224] = i[0];
  assign o[225] = i[0];
  assign o[226] = i[0];
  assign o[227] = i[0];
  assign o[228] = i[0];
  assign o[229] = i[0];
  assign o[230] = i[0];
  assign o[231] = i[0];
  assign o[232] = i[0];
  assign o[233] = i[0];
  assign o[234] = i[0];
  assign o[235] = i[0];
  assign o[236] = i[0];
  assign o[237] = i[0];
  assign o[238] = i[0];
  assign o[239] = i[0];
  assign o[240] = i[0];
  assign o[241] = i[0];
  assign o[242] = i[0];
  assign o[243] = i[0];
  assign o[244] = i[0];
  assign o[245] = i[0];
  assign o[246] = i[0];
  assign o[247] = i[0];
  assign o[248] = i[0];
  assign o[249] = i[0];
  assign o[250] = i[0];
  assign o[251] = i[0];
  assign o[252] = i[0];
  assign o[253] = i[0];
  assign o[254] = i[0];
  assign o[255] = i[0];
  assign o[256] = i[0];
  assign o[257] = i[0];
  assign o[258] = i[0];
  assign o[259] = i[0];
  assign o[260] = i[0];
  assign o[261] = i[0];
  assign o[262] = i[0];
  assign o[263] = i[0];
  assign o[264] = i[0];
  assign o[265] = i[0];
  assign o[266] = i[0];
  assign o[267] = i[0];
  assign o[268] = i[0];
  assign o[269] = i[0];
  assign o[270] = i[0];
  assign o[271] = i[0];
  assign o[272] = i[0];
  assign o[273] = i[0];
  assign o[274] = i[0];
  assign o[275] = i[0];
  assign o[276] = i[0];
  assign o[277] = i[0];
  assign o[278] = i[0];
  assign o[279] = i[0];
  assign o[280] = i[0];
  assign o[281] = i[0];
  assign o[282] = i[0];
  assign o[283] = i[0];
  assign o[284] = i[0];
  assign o[285] = i[0];
  assign o[286] = i[0];
  assign o[287] = i[0];
  assign o[288] = i[0];
  assign o[289] = i[0];
  assign o[290] = i[0];
  assign o[291] = i[0];
  assign o[292] = i[0];
  assign o[293] = i[0];
  assign o[294] = i[0];
  assign o[295] = i[0];
  assign o[296] = i[0];
  assign o[297] = i[0];
  assign o[298] = i[0];
  assign o[299] = i[0];
  assign o[300] = i[0];
  assign o[301] = i[0];
  assign o[302] = i[0];
  assign o[303] = i[0];
  assign o[304] = i[0];
  assign o[305] = i[0];
  assign o[306] = i[0];
  assign o[307] = i[0];
  assign o[308] = i[0];
  assign o[309] = i[0];
  assign o[310] = i[0];
  assign o[311] = i[0];
  assign o[312] = i[0];
  assign o[313] = i[0];
  assign o[314] = i[0];
  assign o[315] = i[0];
  assign o[316] = i[0];
  assign o[317] = i[0];
  assign o[318] = i[0];
  assign o[319] = i[0];
  assign o[320] = i[0];
  assign o[321] = i[0];
  assign o[322] = i[0];
  assign o[323] = i[0];
  assign o[324] = i[0];
  assign o[325] = i[0];
  assign o[326] = i[0];
  assign o[327] = i[0];
  assign o[328] = i[0];
  assign o[329] = i[0];
  assign o[330] = i[0];
  assign o[331] = i[0];
  assign o[332] = i[0];
  assign o[333] = i[0];
  assign o[334] = i[0];
  assign o[335] = i[0];
  assign o[336] = i[0];
  assign o[337] = i[0];
  assign o[338] = i[0];
  assign o[339] = i[0];
  assign o[340] = i[0];
  assign o[341] = i[0];
  assign o[342] = i[0];
  assign o[343] = i[0];
  assign o[344] = i[0];
  assign o[345] = i[0];
  assign o[346] = i[0];
  assign o[347] = i[0];
  assign o[348] = i[0];
  assign o[349] = i[0];
  assign o[350] = i[0];
  assign o[351] = i[0];
  assign o[352] = i[0];
  assign o[353] = i[0];
  assign o[354] = i[0];
  assign o[355] = i[0];
  assign o[356] = i[0];
  assign o[357] = i[0];
  assign o[358] = i[0];
  assign o[359] = i[0];
  assign o[360] = i[0];
  assign o[361] = i[0];
  assign o[362] = i[0];
  assign o[363] = i[0];
  assign o[364] = i[0];
  assign o[365] = i[0];
  assign o[366] = i[0];
  assign o[367] = i[0];
  assign o[368] = i[0];
  assign o[369] = i[0];
  assign o[370] = i[0];
  assign o[371] = i[0];
  assign o[372] = i[0];
  assign o[373] = i[0];
  assign o[374] = i[0];
  assign o[375] = i[0];
  assign o[376] = i[0];
  assign o[377] = i[0];
  assign o[378] = i[0];
  assign o[379] = i[0];
  assign o[380] = i[0];
  assign o[381] = i[0];
  assign o[382] = i[0];
  assign o[383] = i[0];
  assign o[384] = i[0];
  assign o[385] = i[0];
  assign o[386] = i[0];
  assign o[387] = i[0];
  assign o[388] = i[0];
  assign o[389] = i[0];
  assign o[390] = i[0];
  assign o[391] = i[0];
  assign o[392] = i[0];
  assign o[393] = i[0];
  assign o[394] = i[0];
  assign o[395] = i[0];
  assign o[396] = i[0];
  assign o[397] = i[0];
  assign o[398] = i[0];
  assign o[399] = i[0];
  assign o[400] = i[0];
  assign o[401] = i[0];
  assign o[402] = i[0];
  assign o[403] = i[0];
  assign o[404] = i[0];
  assign o[405] = i[0];
  assign o[406] = i[0];
  assign o[407] = i[0];
  assign o[408] = i[0];
  assign o[409] = i[0];
  assign o[410] = i[0];
  assign o[411] = i[0];
  assign o[412] = i[0];
  assign o[413] = i[0];
  assign o[414] = i[0];
  assign o[415] = i[0];
  assign o[416] = i[0];
  assign o[417] = i[0];
  assign o[418] = i[0];
  assign o[419] = i[0];
  assign o[420] = i[0];
  assign o[421] = i[0];
  assign o[422] = i[0];
  assign o[423] = i[0];
  assign o[424] = i[0];
  assign o[425] = i[0];
  assign o[426] = i[0];
  assign o[427] = i[0];
  assign o[428] = i[0];
  assign o[429] = i[0];
  assign o[430] = i[0];
  assign o[431] = i[0];
  assign o[432] = i[0];
  assign o[433] = i[0];
  assign o[434] = i[0];
  assign o[435] = i[0];
  assign o[436] = i[0];
  assign o[437] = i[0];
  assign o[438] = i[0];
  assign o[439] = i[0];
  assign o[440] = i[0];
  assign o[441] = i[0];
  assign o[442] = i[0];
  assign o[443] = i[0];
  assign o[444] = i[0];
  assign o[445] = i[0];
  assign o[446] = i[0];
  assign o[447] = i[0];
  assign o[448] = i[0];
  assign o[449] = i[0];
  assign o[450] = i[0];
  assign o[451] = i[0];
  assign o[452] = i[0];
  assign o[453] = i[0];
  assign o[454] = i[0];
  assign o[455] = i[0];
  assign o[456] = i[0];
  assign o[457] = i[0];
  assign o[458] = i[0];
  assign o[459] = i[0];
  assign o[460] = i[0];
  assign o[461] = i[0];
  assign o[462] = i[0];
  assign o[463] = i[0];
  assign o[464] = i[0];
  assign o[465] = i[0];
  assign o[466] = i[0];
  assign o[467] = i[0];
  assign o[468] = i[0];
  assign o[469] = i[0];
  assign o[470] = i[0];
  assign o[471] = i[0];
  assign o[472] = i[0];
  assign o[473] = i[0];
  assign o[474] = i[0];
  assign o[475] = i[0];
  assign o[476] = i[0];
  assign o[477] = i[0];
  assign o[478] = i[0];
  assign o[479] = i[0];
  assign o[480] = i[0];
  assign o[481] = i[0];
  assign o[482] = i[0];
  assign o[483] = i[0];
  assign o[484] = i[0];
  assign o[485] = i[0];
  assign o[486] = i[0];
  assign o[487] = i[0];
  assign o[488] = i[0];
  assign o[489] = i[0];
  assign o[490] = i[0];
  assign o[491] = i[0];
  assign o[492] = i[0];
  assign o[493] = i[0];
  assign o[494] = i[0];
  assign o[495] = i[0];
  assign o[496] = i[0];
  assign o[497] = i[0];
  assign o[498] = i[0];
  assign o[499] = i[0];
  assign o[500] = i[0];
  assign o[501] = i[0];
  assign o[502] = i[0];
  assign o[503] = i[0];
  assign o[504] = i[0];
  assign o[505] = i[0];
  assign o[506] = i[0];
  assign o[507] = i[0];
  assign o[508] = i[0];
  assign o[509] = i[0];
  assign o[510] = i[0];
  assign o[511] = i[0];

endmodule

