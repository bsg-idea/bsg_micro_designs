

module top
(
  i,
  o
);

  input [31:0] i;
  output [2047:0] o;

  bsg_expand_bitmask
  wrapper
  (
    .i(i),
    .o(o)
  );


endmodule



module bsg_expand_bitmask
(
  i,
  o
);

  input [31:0] i;
  output [2047:0] o;
  wire [2047:0] o;
  assign o[1984] = i[31];
  assign o[1985] = i[31];
  assign o[1986] = i[31];
  assign o[1987] = i[31];
  assign o[1988] = i[31];
  assign o[1989] = i[31];
  assign o[1990] = i[31];
  assign o[1991] = i[31];
  assign o[1992] = i[31];
  assign o[1993] = i[31];
  assign o[1994] = i[31];
  assign o[1995] = i[31];
  assign o[1996] = i[31];
  assign o[1997] = i[31];
  assign o[1998] = i[31];
  assign o[1999] = i[31];
  assign o[2000] = i[31];
  assign o[2001] = i[31];
  assign o[2002] = i[31];
  assign o[2003] = i[31];
  assign o[2004] = i[31];
  assign o[2005] = i[31];
  assign o[2006] = i[31];
  assign o[2007] = i[31];
  assign o[2008] = i[31];
  assign o[2009] = i[31];
  assign o[2010] = i[31];
  assign o[2011] = i[31];
  assign o[2012] = i[31];
  assign o[2013] = i[31];
  assign o[2014] = i[31];
  assign o[2015] = i[31];
  assign o[2016] = i[31];
  assign o[2017] = i[31];
  assign o[2018] = i[31];
  assign o[2019] = i[31];
  assign o[2020] = i[31];
  assign o[2021] = i[31];
  assign o[2022] = i[31];
  assign o[2023] = i[31];
  assign o[2024] = i[31];
  assign o[2025] = i[31];
  assign o[2026] = i[31];
  assign o[2027] = i[31];
  assign o[2028] = i[31];
  assign o[2029] = i[31];
  assign o[2030] = i[31];
  assign o[2031] = i[31];
  assign o[2032] = i[31];
  assign o[2033] = i[31];
  assign o[2034] = i[31];
  assign o[2035] = i[31];
  assign o[2036] = i[31];
  assign o[2037] = i[31];
  assign o[2038] = i[31];
  assign o[2039] = i[31];
  assign o[2040] = i[31];
  assign o[2041] = i[31];
  assign o[2042] = i[31];
  assign o[2043] = i[31];
  assign o[2044] = i[31];
  assign o[2045] = i[31];
  assign o[2046] = i[31];
  assign o[2047] = i[31];
  assign o[1920] = i[30];
  assign o[1921] = i[30];
  assign o[1922] = i[30];
  assign o[1923] = i[30];
  assign o[1924] = i[30];
  assign o[1925] = i[30];
  assign o[1926] = i[30];
  assign o[1927] = i[30];
  assign o[1928] = i[30];
  assign o[1929] = i[30];
  assign o[1930] = i[30];
  assign o[1931] = i[30];
  assign o[1932] = i[30];
  assign o[1933] = i[30];
  assign o[1934] = i[30];
  assign o[1935] = i[30];
  assign o[1936] = i[30];
  assign o[1937] = i[30];
  assign o[1938] = i[30];
  assign o[1939] = i[30];
  assign o[1940] = i[30];
  assign o[1941] = i[30];
  assign o[1942] = i[30];
  assign o[1943] = i[30];
  assign o[1944] = i[30];
  assign o[1945] = i[30];
  assign o[1946] = i[30];
  assign o[1947] = i[30];
  assign o[1948] = i[30];
  assign o[1949] = i[30];
  assign o[1950] = i[30];
  assign o[1951] = i[30];
  assign o[1952] = i[30];
  assign o[1953] = i[30];
  assign o[1954] = i[30];
  assign o[1955] = i[30];
  assign o[1956] = i[30];
  assign o[1957] = i[30];
  assign o[1958] = i[30];
  assign o[1959] = i[30];
  assign o[1960] = i[30];
  assign o[1961] = i[30];
  assign o[1962] = i[30];
  assign o[1963] = i[30];
  assign o[1964] = i[30];
  assign o[1965] = i[30];
  assign o[1966] = i[30];
  assign o[1967] = i[30];
  assign o[1968] = i[30];
  assign o[1969] = i[30];
  assign o[1970] = i[30];
  assign o[1971] = i[30];
  assign o[1972] = i[30];
  assign o[1973] = i[30];
  assign o[1974] = i[30];
  assign o[1975] = i[30];
  assign o[1976] = i[30];
  assign o[1977] = i[30];
  assign o[1978] = i[30];
  assign o[1979] = i[30];
  assign o[1980] = i[30];
  assign o[1981] = i[30];
  assign o[1982] = i[30];
  assign o[1983] = i[30];
  assign o[1856] = i[29];
  assign o[1857] = i[29];
  assign o[1858] = i[29];
  assign o[1859] = i[29];
  assign o[1860] = i[29];
  assign o[1861] = i[29];
  assign o[1862] = i[29];
  assign o[1863] = i[29];
  assign o[1864] = i[29];
  assign o[1865] = i[29];
  assign o[1866] = i[29];
  assign o[1867] = i[29];
  assign o[1868] = i[29];
  assign o[1869] = i[29];
  assign o[1870] = i[29];
  assign o[1871] = i[29];
  assign o[1872] = i[29];
  assign o[1873] = i[29];
  assign o[1874] = i[29];
  assign o[1875] = i[29];
  assign o[1876] = i[29];
  assign o[1877] = i[29];
  assign o[1878] = i[29];
  assign o[1879] = i[29];
  assign o[1880] = i[29];
  assign o[1881] = i[29];
  assign o[1882] = i[29];
  assign o[1883] = i[29];
  assign o[1884] = i[29];
  assign o[1885] = i[29];
  assign o[1886] = i[29];
  assign o[1887] = i[29];
  assign o[1888] = i[29];
  assign o[1889] = i[29];
  assign o[1890] = i[29];
  assign o[1891] = i[29];
  assign o[1892] = i[29];
  assign o[1893] = i[29];
  assign o[1894] = i[29];
  assign o[1895] = i[29];
  assign o[1896] = i[29];
  assign o[1897] = i[29];
  assign o[1898] = i[29];
  assign o[1899] = i[29];
  assign o[1900] = i[29];
  assign o[1901] = i[29];
  assign o[1902] = i[29];
  assign o[1903] = i[29];
  assign o[1904] = i[29];
  assign o[1905] = i[29];
  assign o[1906] = i[29];
  assign o[1907] = i[29];
  assign o[1908] = i[29];
  assign o[1909] = i[29];
  assign o[1910] = i[29];
  assign o[1911] = i[29];
  assign o[1912] = i[29];
  assign o[1913] = i[29];
  assign o[1914] = i[29];
  assign o[1915] = i[29];
  assign o[1916] = i[29];
  assign o[1917] = i[29];
  assign o[1918] = i[29];
  assign o[1919] = i[29];
  assign o[1792] = i[28];
  assign o[1793] = i[28];
  assign o[1794] = i[28];
  assign o[1795] = i[28];
  assign o[1796] = i[28];
  assign o[1797] = i[28];
  assign o[1798] = i[28];
  assign o[1799] = i[28];
  assign o[1800] = i[28];
  assign o[1801] = i[28];
  assign o[1802] = i[28];
  assign o[1803] = i[28];
  assign o[1804] = i[28];
  assign o[1805] = i[28];
  assign o[1806] = i[28];
  assign o[1807] = i[28];
  assign o[1808] = i[28];
  assign o[1809] = i[28];
  assign o[1810] = i[28];
  assign o[1811] = i[28];
  assign o[1812] = i[28];
  assign o[1813] = i[28];
  assign o[1814] = i[28];
  assign o[1815] = i[28];
  assign o[1816] = i[28];
  assign o[1817] = i[28];
  assign o[1818] = i[28];
  assign o[1819] = i[28];
  assign o[1820] = i[28];
  assign o[1821] = i[28];
  assign o[1822] = i[28];
  assign o[1823] = i[28];
  assign o[1824] = i[28];
  assign o[1825] = i[28];
  assign o[1826] = i[28];
  assign o[1827] = i[28];
  assign o[1828] = i[28];
  assign o[1829] = i[28];
  assign o[1830] = i[28];
  assign o[1831] = i[28];
  assign o[1832] = i[28];
  assign o[1833] = i[28];
  assign o[1834] = i[28];
  assign o[1835] = i[28];
  assign o[1836] = i[28];
  assign o[1837] = i[28];
  assign o[1838] = i[28];
  assign o[1839] = i[28];
  assign o[1840] = i[28];
  assign o[1841] = i[28];
  assign o[1842] = i[28];
  assign o[1843] = i[28];
  assign o[1844] = i[28];
  assign o[1845] = i[28];
  assign o[1846] = i[28];
  assign o[1847] = i[28];
  assign o[1848] = i[28];
  assign o[1849] = i[28];
  assign o[1850] = i[28];
  assign o[1851] = i[28];
  assign o[1852] = i[28];
  assign o[1853] = i[28];
  assign o[1854] = i[28];
  assign o[1855] = i[28];
  assign o[1728] = i[27];
  assign o[1729] = i[27];
  assign o[1730] = i[27];
  assign o[1731] = i[27];
  assign o[1732] = i[27];
  assign o[1733] = i[27];
  assign o[1734] = i[27];
  assign o[1735] = i[27];
  assign o[1736] = i[27];
  assign o[1737] = i[27];
  assign o[1738] = i[27];
  assign o[1739] = i[27];
  assign o[1740] = i[27];
  assign o[1741] = i[27];
  assign o[1742] = i[27];
  assign o[1743] = i[27];
  assign o[1744] = i[27];
  assign o[1745] = i[27];
  assign o[1746] = i[27];
  assign o[1747] = i[27];
  assign o[1748] = i[27];
  assign o[1749] = i[27];
  assign o[1750] = i[27];
  assign o[1751] = i[27];
  assign o[1752] = i[27];
  assign o[1753] = i[27];
  assign o[1754] = i[27];
  assign o[1755] = i[27];
  assign o[1756] = i[27];
  assign o[1757] = i[27];
  assign o[1758] = i[27];
  assign o[1759] = i[27];
  assign o[1760] = i[27];
  assign o[1761] = i[27];
  assign o[1762] = i[27];
  assign o[1763] = i[27];
  assign o[1764] = i[27];
  assign o[1765] = i[27];
  assign o[1766] = i[27];
  assign o[1767] = i[27];
  assign o[1768] = i[27];
  assign o[1769] = i[27];
  assign o[1770] = i[27];
  assign o[1771] = i[27];
  assign o[1772] = i[27];
  assign o[1773] = i[27];
  assign o[1774] = i[27];
  assign o[1775] = i[27];
  assign o[1776] = i[27];
  assign o[1777] = i[27];
  assign o[1778] = i[27];
  assign o[1779] = i[27];
  assign o[1780] = i[27];
  assign o[1781] = i[27];
  assign o[1782] = i[27];
  assign o[1783] = i[27];
  assign o[1784] = i[27];
  assign o[1785] = i[27];
  assign o[1786] = i[27];
  assign o[1787] = i[27];
  assign o[1788] = i[27];
  assign o[1789] = i[27];
  assign o[1790] = i[27];
  assign o[1791] = i[27];
  assign o[1664] = i[26];
  assign o[1665] = i[26];
  assign o[1666] = i[26];
  assign o[1667] = i[26];
  assign o[1668] = i[26];
  assign o[1669] = i[26];
  assign o[1670] = i[26];
  assign o[1671] = i[26];
  assign o[1672] = i[26];
  assign o[1673] = i[26];
  assign o[1674] = i[26];
  assign o[1675] = i[26];
  assign o[1676] = i[26];
  assign o[1677] = i[26];
  assign o[1678] = i[26];
  assign o[1679] = i[26];
  assign o[1680] = i[26];
  assign o[1681] = i[26];
  assign o[1682] = i[26];
  assign o[1683] = i[26];
  assign o[1684] = i[26];
  assign o[1685] = i[26];
  assign o[1686] = i[26];
  assign o[1687] = i[26];
  assign o[1688] = i[26];
  assign o[1689] = i[26];
  assign o[1690] = i[26];
  assign o[1691] = i[26];
  assign o[1692] = i[26];
  assign o[1693] = i[26];
  assign o[1694] = i[26];
  assign o[1695] = i[26];
  assign o[1696] = i[26];
  assign o[1697] = i[26];
  assign o[1698] = i[26];
  assign o[1699] = i[26];
  assign o[1700] = i[26];
  assign o[1701] = i[26];
  assign o[1702] = i[26];
  assign o[1703] = i[26];
  assign o[1704] = i[26];
  assign o[1705] = i[26];
  assign o[1706] = i[26];
  assign o[1707] = i[26];
  assign o[1708] = i[26];
  assign o[1709] = i[26];
  assign o[1710] = i[26];
  assign o[1711] = i[26];
  assign o[1712] = i[26];
  assign o[1713] = i[26];
  assign o[1714] = i[26];
  assign o[1715] = i[26];
  assign o[1716] = i[26];
  assign o[1717] = i[26];
  assign o[1718] = i[26];
  assign o[1719] = i[26];
  assign o[1720] = i[26];
  assign o[1721] = i[26];
  assign o[1722] = i[26];
  assign o[1723] = i[26];
  assign o[1724] = i[26];
  assign o[1725] = i[26];
  assign o[1726] = i[26];
  assign o[1727] = i[26];
  assign o[1600] = i[25];
  assign o[1601] = i[25];
  assign o[1602] = i[25];
  assign o[1603] = i[25];
  assign o[1604] = i[25];
  assign o[1605] = i[25];
  assign o[1606] = i[25];
  assign o[1607] = i[25];
  assign o[1608] = i[25];
  assign o[1609] = i[25];
  assign o[1610] = i[25];
  assign o[1611] = i[25];
  assign o[1612] = i[25];
  assign o[1613] = i[25];
  assign o[1614] = i[25];
  assign o[1615] = i[25];
  assign o[1616] = i[25];
  assign o[1617] = i[25];
  assign o[1618] = i[25];
  assign o[1619] = i[25];
  assign o[1620] = i[25];
  assign o[1621] = i[25];
  assign o[1622] = i[25];
  assign o[1623] = i[25];
  assign o[1624] = i[25];
  assign o[1625] = i[25];
  assign o[1626] = i[25];
  assign o[1627] = i[25];
  assign o[1628] = i[25];
  assign o[1629] = i[25];
  assign o[1630] = i[25];
  assign o[1631] = i[25];
  assign o[1632] = i[25];
  assign o[1633] = i[25];
  assign o[1634] = i[25];
  assign o[1635] = i[25];
  assign o[1636] = i[25];
  assign o[1637] = i[25];
  assign o[1638] = i[25];
  assign o[1639] = i[25];
  assign o[1640] = i[25];
  assign o[1641] = i[25];
  assign o[1642] = i[25];
  assign o[1643] = i[25];
  assign o[1644] = i[25];
  assign o[1645] = i[25];
  assign o[1646] = i[25];
  assign o[1647] = i[25];
  assign o[1648] = i[25];
  assign o[1649] = i[25];
  assign o[1650] = i[25];
  assign o[1651] = i[25];
  assign o[1652] = i[25];
  assign o[1653] = i[25];
  assign o[1654] = i[25];
  assign o[1655] = i[25];
  assign o[1656] = i[25];
  assign o[1657] = i[25];
  assign o[1658] = i[25];
  assign o[1659] = i[25];
  assign o[1660] = i[25];
  assign o[1661] = i[25];
  assign o[1662] = i[25];
  assign o[1663] = i[25];
  assign o[1536] = i[24];
  assign o[1537] = i[24];
  assign o[1538] = i[24];
  assign o[1539] = i[24];
  assign o[1540] = i[24];
  assign o[1541] = i[24];
  assign o[1542] = i[24];
  assign o[1543] = i[24];
  assign o[1544] = i[24];
  assign o[1545] = i[24];
  assign o[1546] = i[24];
  assign o[1547] = i[24];
  assign o[1548] = i[24];
  assign o[1549] = i[24];
  assign o[1550] = i[24];
  assign o[1551] = i[24];
  assign o[1552] = i[24];
  assign o[1553] = i[24];
  assign o[1554] = i[24];
  assign o[1555] = i[24];
  assign o[1556] = i[24];
  assign o[1557] = i[24];
  assign o[1558] = i[24];
  assign o[1559] = i[24];
  assign o[1560] = i[24];
  assign o[1561] = i[24];
  assign o[1562] = i[24];
  assign o[1563] = i[24];
  assign o[1564] = i[24];
  assign o[1565] = i[24];
  assign o[1566] = i[24];
  assign o[1567] = i[24];
  assign o[1568] = i[24];
  assign o[1569] = i[24];
  assign o[1570] = i[24];
  assign o[1571] = i[24];
  assign o[1572] = i[24];
  assign o[1573] = i[24];
  assign o[1574] = i[24];
  assign o[1575] = i[24];
  assign o[1576] = i[24];
  assign o[1577] = i[24];
  assign o[1578] = i[24];
  assign o[1579] = i[24];
  assign o[1580] = i[24];
  assign o[1581] = i[24];
  assign o[1582] = i[24];
  assign o[1583] = i[24];
  assign o[1584] = i[24];
  assign o[1585] = i[24];
  assign o[1586] = i[24];
  assign o[1587] = i[24];
  assign o[1588] = i[24];
  assign o[1589] = i[24];
  assign o[1590] = i[24];
  assign o[1591] = i[24];
  assign o[1592] = i[24];
  assign o[1593] = i[24];
  assign o[1594] = i[24];
  assign o[1595] = i[24];
  assign o[1596] = i[24];
  assign o[1597] = i[24];
  assign o[1598] = i[24];
  assign o[1599] = i[24];
  assign o[1472] = i[23];
  assign o[1473] = i[23];
  assign o[1474] = i[23];
  assign o[1475] = i[23];
  assign o[1476] = i[23];
  assign o[1477] = i[23];
  assign o[1478] = i[23];
  assign o[1479] = i[23];
  assign o[1480] = i[23];
  assign o[1481] = i[23];
  assign o[1482] = i[23];
  assign o[1483] = i[23];
  assign o[1484] = i[23];
  assign o[1485] = i[23];
  assign o[1486] = i[23];
  assign o[1487] = i[23];
  assign o[1488] = i[23];
  assign o[1489] = i[23];
  assign o[1490] = i[23];
  assign o[1491] = i[23];
  assign o[1492] = i[23];
  assign o[1493] = i[23];
  assign o[1494] = i[23];
  assign o[1495] = i[23];
  assign o[1496] = i[23];
  assign o[1497] = i[23];
  assign o[1498] = i[23];
  assign o[1499] = i[23];
  assign o[1500] = i[23];
  assign o[1501] = i[23];
  assign o[1502] = i[23];
  assign o[1503] = i[23];
  assign o[1504] = i[23];
  assign o[1505] = i[23];
  assign o[1506] = i[23];
  assign o[1507] = i[23];
  assign o[1508] = i[23];
  assign o[1509] = i[23];
  assign o[1510] = i[23];
  assign o[1511] = i[23];
  assign o[1512] = i[23];
  assign o[1513] = i[23];
  assign o[1514] = i[23];
  assign o[1515] = i[23];
  assign o[1516] = i[23];
  assign o[1517] = i[23];
  assign o[1518] = i[23];
  assign o[1519] = i[23];
  assign o[1520] = i[23];
  assign o[1521] = i[23];
  assign o[1522] = i[23];
  assign o[1523] = i[23];
  assign o[1524] = i[23];
  assign o[1525] = i[23];
  assign o[1526] = i[23];
  assign o[1527] = i[23];
  assign o[1528] = i[23];
  assign o[1529] = i[23];
  assign o[1530] = i[23];
  assign o[1531] = i[23];
  assign o[1532] = i[23];
  assign o[1533] = i[23];
  assign o[1534] = i[23];
  assign o[1535] = i[23];
  assign o[1408] = i[22];
  assign o[1409] = i[22];
  assign o[1410] = i[22];
  assign o[1411] = i[22];
  assign o[1412] = i[22];
  assign o[1413] = i[22];
  assign o[1414] = i[22];
  assign o[1415] = i[22];
  assign o[1416] = i[22];
  assign o[1417] = i[22];
  assign o[1418] = i[22];
  assign o[1419] = i[22];
  assign o[1420] = i[22];
  assign o[1421] = i[22];
  assign o[1422] = i[22];
  assign o[1423] = i[22];
  assign o[1424] = i[22];
  assign o[1425] = i[22];
  assign o[1426] = i[22];
  assign o[1427] = i[22];
  assign o[1428] = i[22];
  assign o[1429] = i[22];
  assign o[1430] = i[22];
  assign o[1431] = i[22];
  assign o[1432] = i[22];
  assign o[1433] = i[22];
  assign o[1434] = i[22];
  assign o[1435] = i[22];
  assign o[1436] = i[22];
  assign o[1437] = i[22];
  assign o[1438] = i[22];
  assign o[1439] = i[22];
  assign o[1440] = i[22];
  assign o[1441] = i[22];
  assign o[1442] = i[22];
  assign o[1443] = i[22];
  assign o[1444] = i[22];
  assign o[1445] = i[22];
  assign o[1446] = i[22];
  assign o[1447] = i[22];
  assign o[1448] = i[22];
  assign o[1449] = i[22];
  assign o[1450] = i[22];
  assign o[1451] = i[22];
  assign o[1452] = i[22];
  assign o[1453] = i[22];
  assign o[1454] = i[22];
  assign o[1455] = i[22];
  assign o[1456] = i[22];
  assign o[1457] = i[22];
  assign o[1458] = i[22];
  assign o[1459] = i[22];
  assign o[1460] = i[22];
  assign o[1461] = i[22];
  assign o[1462] = i[22];
  assign o[1463] = i[22];
  assign o[1464] = i[22];
  assign o[1465] = i[22];
  assign o[1466] = i[22];
  assign o[1467] = i[22];
  assign o[1468] = i[22];
  assign o[1469] = i[22];
  assign o[1470] = i[22];
  assign o[1471] = i[22];
  assign o[1344] = i[21];
  assign o[1345] = i[21];
  assign o[1346] = i[21];
  assign o[1347] = i[21];
  assign o[1348] = i[21];
  assign o[1349] = i[21];
  assign o[1350] = i[21];
  assign o[1351] = i[21];
  assign o[1352] = i[21];
  assign o[1353] = i[21];
  assign o[1354] = i[21];
  assign o[1355] = i[21];
  assign o[1356] = i[21];
  assign o[1357] = i[21];
  assign o[1358] = i[21];
  assign o[1359] = i[21];
  assign o[1360] = i[21];
  assign o[1361] = i[21];
  assign o[1362] = i[21];
  assign o[1363] = i[21];
  assign o[1364] = i[21];
  assign o[1365] = i[21];
  assign o[1366] = i[21];
  assign o[1367] = i[21];
  assign o[1368] = i[21];
  assign o[1369] = i[21];
  assign o[1370] = i[21];
  assign o[1371] = i[21];
  assign o[1372] = i[21];
  assign o[1373] = i[21];
  assign o[1374] = i[21];
  assign o[1375] = i[21];
  assign o[1376] = i[21];
  assign o[1377] = i[21];
  assign o[1378] = i[21];
  assign o[1379] = i[21];
  assign o[1380] = i[21];
  assign o[1381] = i[21];
  assign o[1382] = i[21];
  assign o[1383] = i[21];
  assign o[1384] = i[21];
  assign o[1385] = i[21];
  assign o[1386] = i[21];
  assign o[1387] = i[21];
  assign o[1388] = i[21];
  assign o[1389] = i[21];
  assign o[1390] = i[21];
  assign o[1391] = i[21];
  assign o[1392] = i[21];
  assign o[1393] = i[21];
  assign o[1394] = i[21];
  assign o[1395] = i[21];
  assign o[1396] = i[21];
  assign o[1397] = i[21];
  assign o[1398] = i[21];
  assign o[1399] = i[21];
  assign o[1400] = i[21];
  assign o[1401] = i[21];
  assign o[1402] = i[21];
  assign o[1403] = i[21];
  assign o[1404] = i[21];
  assign o[1405] = i[21];
  assign o[1406] = i[21];
  assign o[1407] = i[21];
  assign o[1280] = i[20];
  assign o[1281] = i[20];
  assign o[1282] = i[20];
  assign o[1283] = i[20];
  assign o[1284] = i[20];
  assign o[1285] = i[20];
  assign o[1286] = i[20];
  assign o[1287] = i[20];
  assign o[1288] = i[20];
  assign o[1289] = i[20];
  assign o[1290] = i[20];
  assign o[1291] = i[20];
  assign o[1292] = i[20];
  assign o[1293] = i[20];
  assign o[1294] = i[20];
  assign o[1295] = i[20];
  assign o[1296] = i[20];
  assign o[1297] = i[20];
  assign o[1298] = i[20];
  assign o[1299] = i[20];
  assign o[1300] = i[20];
  assign o[1301] = i[20];
  assign o[1302] = i[20];
  assign o[1303] = i[20];
  assign o[1304] = i[20];
  assign o[1305] = i[20];
  assign o[1306] = i[20];
  assign o[1307] = i[20];
  assign o[1308] = i[20];
  assign o[1309] = i[20];
  assign o[1310] = i[20];
  assign o[1311] = i[20];
  assign o[1312] = i[20];
  assign o[1313] = i[20];
  assign o[1314] = i[20];
  assign o[1315] = i[20];
  assign o[1316] = i[20];
  assign o[1317] = i[20];
  assign o[1318] = i[20];
  assign o[1319] = i[20];
  assign o[1320] = i[20];
  assign o[1321] = i[20];
  assign o[1322] = i[20];
  assign o[1323] = i[20];
  assign o[1324] = i[20];
  assign o[1325] = i[20];
  assign o[1326] = i[20];
  assign o[1327] = i[20];
  assign o[1328] = i[20];
  assign o[1329] = i[20];
  assign o[1330] = i[20];
  assign o[1331] = i[20];
  assign o[1332] = i[20];
  assign o[1333] = i[20];
  assign o[1334] = i[20];
  assign o[1335] = i[20];
  assign o[1336] = i[20];
  assign o[1337] = i[20];
  assign o[1338] = i[20];
  assign o[1339] = i[20];
  assign o[1340] = i[20];
  assign o[1341] = i[20];
  assign o[1342] = i[20];
  assign o[1343] = i[20];
  assign o[1216] = i[19];
  assign o[1217] = i[19];
  assign o[1218] = i[19];
  assign o[1219] = i[19];
  assign o[1220] = i[19];
  assign o[1221] = i[19];
  assign o[1222] = i[19];
  assign o[1223] = i[19];
  assign o[1224] = i[19];
  assign o[1225] = i[19];
  assign o[1226] = i[19];
  assign o[1227] = i[19];
  assign o[1228] = i[19];
  assign o[1229] = i[19];
  assign o[1230] = i[19];
  assign o[1231] = i[19];
  assign o[1232] = i[19];
  assign o[1233] = i[19];
  assign o[1234] = i[19];
  assign o[1235] = i[19];
  assign o[1236] = i[19];
  assign o[1237] = i[19];
  assign o[1238] = i[19];
  assign o[1239] = i[19];
  assign o[1240] = i[19];
  assign o[1241] = i[19];
  assign o[1242] = i[19];
  assign o[1243] = i[19];
  assign o[1244] = i[19];
  assign o[1245] = i[19];
  assign o[1246] = i[19];
  assign o[1247] = i[19];
  assign o[1248] = i[19];
  assign o[1249] = i[19];
  assign o[1250] = i[19];
  assign o[1251] = i[19];
  assign o[1252] = i[19];
  assign o[1253] = i[19];
  assign o[1254] = i[19];
  assign o[1255] = i[19];
  assign o[1256] = i[19];
  assign o[1257] = i[19];
  assign o[1258] = i[19];
  assign o[1259] = i[19];
  assign o[1260] = i[19];
  assign o[1261] = i[19];
  assign o[1262] = i[19];
  assign o[1263] = i[19];
  assign o[1264] = i[19];
  assign o[1265] = i[19];
  assign o[1266] = i[19];
  assign o[1267] = i[19];
  assign o[1268] = i[19];
  assign o[1269] = i[19];
  assign o[1270] = i[19];
  assign o[1271] = i[19];
  assign o[1272] = i[19];
  assign o[1273] = i[19];
  assign o[1274] = i[19];
  assign o[1275] = i[19];
  assign o[1276] = i[19];
  assign o[1277] = i[19];
  assign o[1278] = i[19];
  assign o[1279] = i[19];
  assign o[1152] = i[18];
  assign o[1153] = i[18];
  assign o[1154] = i[18];
  assign o[1155] = i[18];
  assign o[1156] = i[18];
  assign o[1157] = i[18];
  assign o[1158] = i[18];
  assign o[1159] = i[18];
  assign o[1160] = i[18];
  assign o[1161] = i[18];
  assign o[1162] = i[18];
  assign o[1163] = i[18];
  assign o[1164] = i[18];
  assign o[1165] = i[18];
  assign o[1166] = i[18];
  assign o[1167] = i[18];
  assign o[1168] = i[18];
  assign o[1169] = i[18];
  assign o[1170] = i[18];
  assign o[1171] = i[18];
  assign o[1172] = i[18];
  assign o[1173] = i[18];
  assign o[1174] = i[18];
  assign o[1175] = i[18];
  assign o[1176] = i[18];
  assign o[1177] = i[18];
  assign o[1178] = i[18];
  assign o[1179] = i[18];
  assign o[1180] = i[18];
  assign o[1181] = i[18];
  assign o[1182] = i[18];
  assign o[1183] = i[18];
  assign o[1184] = i[18];
  assign o[1185] = i[18];
  assign o[1186] = i[18];
  assign o[1187] = i[18];
  assign o[1188] = i[18];
  assign o[1189] = i[18];
  assign o[1190] = i[18];
  assign o[1191] = i[18];
  assign o[1192] = i[18];
  assign o[1193] = i[18];
  assign o[1194] = i[18];
  assign o[1195] = i[18];
  assign o[1196] = i[18];
  assign o[1197] = i[18];
  assign o[1198] = i[18];
  assign o[1199] = i[18];
  assign o[1200] = i[18];
  assign o[1201] = i[18];
  assign o[1202] = i[18];
  assign o[1203] = i[18];
  assign o[1204] = i[18];
  assign o[1205] = i[18];
  assign o[1206] = i[18];
  assign o[1207] = i[18];
  assign o[1208] = i[18];
  assign o[1209] = i[18];
  assign o[1210] = i[18];
  assign o[1211] = i[18];
  assign o[1212] = i[18];
  assign o[1213] = i[18];
  assign o[1214] = i[18];
  assign o[1215] = i[18];
  assign o[1088] = i[17];
  assign o[1089] = i[17];
  assign o[1090] = i[17];
  assign o[1091] = i[17];
  assign o[1092] = i[17];
  assign o[1093] = i[17];
  assign o[1094] = i[17];
  assign o[1095] = i[17];
  assign o[1096] = i[17];
  assign o[1097] = i[17];
  assign o[1098] = i[17];
  assign o[1099] = i[17];
  assign o[1100] = i[17];
  assign o[1101] = i[17];
  assign o[1102] = i[17];
  assign o[1103] = i[17];
  assign o[1104] = i[17];
  assign o[1105] = i[17];
  assign o[1106] = i[17];
  assign o[1107] = i[17];
  assign o[1108] = i[17];
  assign o[1109] = i[17];
  assign o[1110] = i[17];
  assign o[1111] = i[17];
  assign o[1112] = i[17];
  assign o[1113] = i[17];
  assign o[1114] = i[17];
  assign o[1115] = i[17];
  assign o[1116] = i[17];
  assign o[1117] = i[17];
  assign o[1118] = i[17];
  assign o[1119] = i[17];
  assign o[1120] = i[17];
  assign o[1121] = i[17];
  assign o[1122] = i[17];
  assign o[1123] = i[17];
  assign o[1124] = i[17];
  assign o[1125] = i[17];
  assign o[1126] = i[17];
  assign o[1127] = i[17];
  assign o[1128] = i[17];
  assign o[1129] = i[17];
  assign o[1130] = i[17];
  assign o[1131] = i[17];
  assign o[1132] = i[17];
  assign o[1133] = i[17];
  assign o[1134] = i[17];
  assign o[1135] = i[17];
  assign o[1136] = i[17];
  assign o[1137] = i[17];
  assign o[1138] = i[17];
  assign o[1139] = i[17];
  assign o[1140] = i[17];
  assign o[1141] = i[17];
  assign o[1142] = i[17];
  assign o[1143] = i[17];
  assign o[1144] = i[17];
  assign o[1145] = i[17];
  assign o[1146] = i[17];
  assign o[1147] = i[17];
  assign o[1148] = i[17];
  assign o[1149] = i[17];
  assign o[1150] = i[17];
  assign o[1151] = i[17];
  assign o[1024] = i[16];
  assign o[1025] = i[16];
  assign o[1026] = i[16];
  assign o[1027] = i[16];
  assign o[1028] = i[16];
  assign o[1029] = i[16];
  assign o[1030] = i[16];
  assign o[1031] = i[16];
  assign o[1032] = i[16];
  assign o[1033] = i[16];
  assign o[1034] = i[16];
  assign o[1035] = i[16];
  assign o[1036] = i[16];
  assign o[1037] = i[16];
  assign o[1038] = i[16];
  assign o[1039] = i[16];
  assign o[1040] = i[16];
  assign o[1041] = i[16];
  assign o[1042] = i[16];
  assign o[1043] = i[16];
  assign o[1044] = i[16];
  assign o[1045] = i[16];
  assign o[1046] = i[16];
  assign o[1047] = i[16];
  assign o[1048] = i[16];
  assign o[1049] = i[16];
  assign o[1050] = i[16];
  assign o[1051] = i[16];
  assign o[1052] = i[16];
  assign o[1053] = i[16];
  assign o[1054] = i[16];
  assign o[1055] = i[16];
  assign o[1056] = i[16];
  assign o[1057] = i[16];
  assign o[1058] = i[16];
  assign o[1059] = i[16];
  assign o[1060] = i[16];
  assign o[1061] = i[16];
  assign o[1062] = i[16];
  assign o[1063] = i[16];
  assign o[1064] = i[16];
  assign o[1065] = i[16];
  assign o[1066] = i[16];
  assign o[1067] = i[16];
  assign o[1068] = i[16];
  assign o[1069] = i[16];
  assign o[1070] = i[16];
  assign o[1071] = i[16];
  assign o[1072] = i[16];
  assign o[1073] = i[16];
  assign o[1074] = i[16];
  assign o[1075] = i[16];
  assign o[1076] = i[16];
  assign o[1077] = i[16];
  assign o[1078] = i[16];
  assign o[1079] = i[16];
  assign o[1080] = i[16];
  assign o[1081] = i[16];
  assign o[1082] = i[16];
  assign o[1083] = i[16];
  assign o[1084] = i[16];
  assign o[1085] = i[16];
  assign o[1086] = i[16];
  assign o[1087] = i[16];
  assign o[960] = i[15];
  assign o[961] = i[15];
  assign o[962] = i[15];
  assign o[963] = i[15];
  assign o[964] = i[15];
  assign o[965] = i[15];
  assign o[966] = i[15];
  assign o[967] = i[15];
  assign o[968] = i[15];
  assign o[969] = i[15];
  assign o[970] = i[15];
  assign o[971] = i[15];
  assign o[972] = i[15];
  assign o[973] = i[15];
  assign o[974] = i[15];
  assign o[975] = i[15];
  assign o[976] = i[15];
  assign o[977] = i[15];
  assign o[978] = i[15];
  assign o[979] = i[15];
  assign o[980] = i[15];
  assign o[981] = i[15];
  assign o[982] = i[15];
  assign o[983] = i[15];
  assign o[984] = i[15];
  assign o[985] = i[15];
  assign o[986] = i[15];
  assign o[987] = i[15];
  assign o[988] = i[15];
  assign o[989] = i[15];
  assign o[990] = i[15];
  assign o[991] = i[15];
  assign o[992] = i[15];
  assign o[993] = i[15];
  assign o[994] = i[15];
  assign o[995] = i[15];
  assign o[996] = i[15];
  assign o[997] = i[15];
  assign o[998] = i[15];
  assign o[999] = i[15];
  assign o[1000] = i[15];
  assign o[1001] = i[15];
  assign o[1002] = i[15];
  assign o[1003] = i[15];
  assign o[1004] = i[15];
  assign o[1005] = i[15];
  assign o[1006] = i[15];
  assign o[1007] = i[15];
  assign o[1008] = i[15];
  assign o[1009] = i[15];
  assign o[1010] = i[15];
  assign o[1011] = i[15];
  assign o[1012] = i[15];
  assign o[1013] = i[15];
  assign o[1014] = i[15];
  assign o[1015] = i[15];
  assign o[1016] = i[15];
  assign o[1017] = i[15];
  assign o[1018] = i[15];
  assign o[1019] = i[15];
  assign o[1020] = i[15];
  assign o[1021] = i[15];
  assign o[1022] = i[15];
  assign o[1023] = i[15];
  assign o[896] = i[14];
  assign o[897] = i[14];
  assign o[898] = i[14];
  assign o[899] = i[14];
  assign o[900] = i[14];
  assign o[901] = i[14];
  assign o[902] = i[14];
  assign o[903] = i[14];
  assign o[904] = i[14];
  assign o[905] = i[14];
  assign o[906] = i[14];
  assign o[907] = i[14];
  assign o[908] = i[14];
  assign o[909] = i[14];
  assign o[910] = i[14];
  assign o[911] = i[14];
  assign o[912] = i[14];
  assign o[913] = i[14];
  assign o[914] = i[14];
  assign o[915] = i[14];
  assign o[916] = i[14];
  assign o[917] = i[14];
  assign o[918] = i[14];
  assign o[919] = i[14];
  assign o[920] = i[14];
  assign o[921] = i[14];
  assign o[922] = i[14];
  assign o[923] = i[14];
  assign o[924] = i[14];
  assign o[925] = i[14];
  assign o[926] = i[14];
  assign o[927] = i[14];
  assign o[928] = i[14];
  assign o[929] = i[14];
  assign o[930] = i[14];
  assign o[931] = i[14];
  assign o[932] = i[14];
  assign o[933] = i[14];
  assign o[934] = i[14];
  assign o[935] = i[14];
  assign o[936] = i[14];
  assign o[937] = i[14];
  assign o[938] = i[14];
  assign o[939] = i[14];
  assign o[940] = i[14];
  assign o[941] = i[14];
  assign o[942] = i[14];
  assign o[943] = i[14];
  assign o[944] = i[14];
  assign o[945] = i[14];
  assign o[946] = i[14];
  assign o[947] = i[14];
  assign o[948] = i[14];
  assign o[949] = i[14];
  assign o[950] = i[14];
  assign o[951] = i[14];
  assign o[952] = i[14];
  assign o[953] = i[14];
  assign o[954] = i[14];
  assign o[955] = i[14];
  assign o[956] = i[14];
  assign o[957] = i[14];
  assign o[958] = i[14];
  assign o[959] = i[14];
  assign o[832] = i[13];
  assign o[833] = i[13];
  assign o[834] = i[13];
  assign o[835] = i[13];
  assign o[836] = i[13];
  assign o[837] = i[13];
  assign o[838] = i[13];
  assign o[839] = i[13];
  assign o[840] = i[13];
  assign o[841] = i[13];
  assign o[842] = i[13];
  assign o[843] = i[13];
  assign o[844] = i[13];
  assign o[845] = i[13];
  assign o[846] = i[13];
  assign o[847] = i[13];
  assign o[848] = i[13];
  assign o[849] = i[13];
  assign o[850] = i[13];
  assign o[851] = i[13];
  assign o[852] = i[13];
  assign o[853] = i[13];
  assign o[854] = i[13];
  assign o[855] = i[13];
  assign o[856] = i[13];
  assign o[857] = i[13];
  assign o[858] = i[13];
  assign o[859] = i[13];
  assign o[860] = i[13];
  assign o[861] = i[13];
  assign o[862] = i[13];
  assign o[863] = i[13];
  assign o[864] = i[13];
  assign o[865] = i[13];
  assign o[866] = i[13];
  assign o[867] = i[13];
  assign o[868] = i[13];
  assign o[869] = i[13];
  assign o[870] = i[13];
  assign o[871] = i[13];
  assign o[872] = i[13];
  assign o[873] = i[13];
  assign o[874] = i[13];
  assign o[875] = i[13];
  assign o[876] = i[13];
  assign o[877] = i[13];
  assign o[878] = i[13];
  assign o[879] = i[13];
  assign o[880] = i[13];
  assign o[881] = i[13];
  assign o[882] = i[13];
  assign o[883] = i[13];
  assign o[884] = i[13];
  assign o[885] = i[13];
  assign o[886] = i[13];
  assign o[887] = i[13];
  assign o[888] = i[13];
  assign o[889] = i[13];
  assign o[890] = i[13];
  assign o[891] = i[13];
  assign o[892] = i[13];
  assign o[893] = i[13];
  assign o[894] = i[13];
  assign o[895] = i[13];
  assign o[768] = i[12];
  assign o[769] = i[12];
  assign o[770] = i[12];
  assign o[771] = i[12];
  assign o[772] = i[12];
  assign o[773] = i[12];
  assign o[774] = i[12];
  assign o[775] = i[12];
  assign o[776] = i[12];
  assign o[777] = i[12];
  assign o[778] = i[12];
  assign o[779] = i[12];
  assign o[780] = i[12];
  assign o[781] = i[12];
  assign o[782] = i[12];
  assign o[783] = i[12];
  assign o[784] = i[12];
  assign o[785] = i[12];
  assign o[786] = i[12];
  assign o[787] = i[12];
  assign o[788] = i[12];
  assign o[789] = i[12];
  assign o[790] = i[12];
  assign o[791] = i[12];
  assign o[792] = i[12];
  assign o[793] = i[12];
  assign o[794] = i[12];
  assign o[795] = i[12];
  assign o[796] = i[12];
  assign o[797] = i[12];
  assign o[798] = i[12];
  assign o[799] = i[12];
  assign o[800] = i[12];
  assign o[801] = i[12];
  assign o[802] = i[12];
  assign o[803] = i[12];
  assign o[804] = i[12];
  assign o[805] = i[12];
  assign o[806] = i[12];
  assign o[807] = i[12];
  assign o[808] = i[12];
  assign o[809] = i[12];
  assign o[810] = i[12];
  assign o[811] = i[12];
  assign o[812] = i[12];
  assign o[813] = i[12];
  assign o[814] = i[12];
  assign o[815] = i[12];
  assign o[816] = i[12];
  assign o[817] = i[12];
  assign o[818] = i[12];
  assign o[819] = i[12];
  assign o[820] = i[12];
  assign o[821] = i[12];
  assign o[822] = i[12];
  assign o[823] = i[12];
  assign o[824] = i[12];
  assign o[825] = i[12];
  assign o[826] = i[12];
  assign o[827] = i[12];
  assign o[828] = i[12];
  assign o[829] = i[12];
  assign o[830] = i[12];
  assign o[831] = i[12];
  assign o[704] = i[11];
  assign o[705] = i[11];
  assign o[706] = i[11];
  assign o[707] = i[11];
  assign o[708] = i[11];
  assign o[709] = i[11];
  assign o[710] = i[11];
  assign o[711] = i[11];
  assign o[712] = i[11];
  assign o[713] = i[11];
  assign o[714] = i[11];
  assign o[715] = i[11];
  assign o[716] = i[11];
  assign o[717] = i[11];
  assign o[718] = i[11];
  assign o[719] = i[11];
  assign o[720] = i[11];
  assign o[721] = i[11];
  assign o[722] = i[11];
  assign o[723] = i[11];
  assign o[724] = i[11];
  assign o[725] = i[11];
  assign o[726] = i[11];
  assign o[727] = i[11];
  assign o[728] = i[11];
  assign o[729] = i[11];
  assign o[730] = i[11];
  assign o[731] = i[11];
  assign o[732] = i[11];
  assign o[733] = i[11];
  assign o[734] = i[11];
  assign o[735] = i[11];
  assign o[736] = i[11];
  assign o[737] = i[11];
  assign o[738] = i[11];
  assign o[739] = i[11];
  assign o[740] = i[11];
  assign o[741] = i[11];
  assign o[742] = i[11];
  assign o[743] = i[11];
  assign o[744] = i[11];
  assign o[745] = i[11];
  assign o[746] = i[11];
  assign o[747] = i[11];
  assign o[748] = i[11];
  assign o[749] = i[11];
  assign o[750] = i[11];
  assign o[751] = i[11];
  assign o[752] = i[11];
  assign o[753] = i[11];
  assign o[754] = i[11];
  assign o[755] = i[11];
  assign o[756] = i[11];
  assign o[757] = i[11];
  assign o[758] = i[11];
  assign o[759] = i[11];
  assign o[760] = i[11];
  assign o[761] = i[11];
  assign o[762] = i[11];
  assign o[763] = i[11];
  assign o[764] = i[11];
  assign o[765] = i[11];
  assign o[766] = i[11];
  assign o[767] = i[11];
  assign o[640] = i[10];
  assign o[641] = i[10];
  assign o[642] = i[10];
  assign o[643] = i[10];
  assign o[644] = i[10];
  assign o[645] = i[10];
  assign o[646] = i[10];
  assign o[647] = i[10];
  assign o[648] = i[10];
  assign o[649] = i[10];
  assign o[650] = i[10];
  assign o[651] = i[10];
  assign o[652] = i[10];
  assign o[653] = i[10];
  assign o[654] = i[10];
  assign o[655] = i[10];
  assign o[656] = i[10];
  assign o[657] = i[10];
  assign o[658] = i[10];
  assign o[659] = i[10];
  assign o[660] = i[10];
  assign o[661] = i[10];
  assign o[662] = i[10];
  assign o[663] = i[10];
  assign o[664] = i[10];
  assign o[665] = i[10];
  assign o[666] = i[10];
  assign o[667] = i[10];
  assign o[668] = i[10];
  assign o[669] = i[10];
  assign o[670] = i[10];
  assign o[671] = i[10];
  assign o[672] = i[10];
  assign o[673] = i[10];
  assign o[674] = i[10];
  assign o[675] = i[10];
  assign o[676] = i[10];
  assign o[677] = i[10];
  assign o[678] = i[10];
  assign o[679] = i[10];
  assign o[680] = i[10];
  assign o[681] = i[10];
  assign o[682] = i[10];
  assign o[683] = i[10];
  assign o[684] = i[10];
  assign o[685] = i[10];
  assign o[686] = i[10];
  assign o[687] = i[10];
  assign o[688] = i[10];
  assign o[689] = i[10];
  assign o[690] = i[10];
  assign o[691] = i[10];
  assign o[692] = i[10];
  assign o[693] = i[10];
  assign o[694] = i[10];
  assign o[695] = i[10];
  assign o[696] = i[10];
  assign o[697] = i[10];
  assign o[698] = i[10];
  assign o[699] = i[10];
  assign o[700] = i[10];
  assign o[701] = i[10];
  assign o[702] = i[10];
  assign o[703] = i[10];
  assign o[576] = i[9];
  assign o[577] = i[9];
  assign o[578] = i[9];
  assign o[579] = i[9];
  assign o[580] = i[9];
  assign o[581] = i[9];
  assign o[582] = i[9];
  assign o[583] = i[9];
  assign o[584] = i[9];
  assign o[585] = i[9];
  assign o[586] = i[9];
  assign o[587] = i[9];
  assign o[588] = i[9];
  assign o[589] = i[9];
  assign o[590] = i[9];
  assign o[591] = i[9];
  assign o[592] = i[9];
  assign o[593] = i[9];
  assign o[594] = i[9];
  assign o[595] = i[9];
  assign o[596] = i[9];
  assign o[597] = i[9];
  assign o[598] = i[9];
  assign o[599] = i[9];
  assign o[600] = i[9];
  assign o[601] = i[9];
  assign o[602] = i[9];
  assign o[603] = i[9];
  assign o[604] = i[9];
  assign o[605] = i[9];
  assign o[606] = i[9];
  assign o[607] = i[9];
  assign o[608] = i[9];
  assign o[609] = i[9];
  assign o[610] = i[9];
  assign o[611] = i[9];
  assign o[612] = i[9];
  assign o[613] = i[9];
  assign o[614] = i[9];
  assign o[615] = i[9];
  assign o[616] = i[9];
  assign o[617] = i[9];
  assign o[618] = i[9];
  assign o[619] = i[9];
  assign o[620] = i[9];
  assign o[621] = i[9];
  assign o[622] = i[9];
  assign o[623] = i[9];
  assign o[624] = i[9];
  assign o[625] = i[9];
  assign o[626] = i[9];
  assign o[627] = i[9];
  assign o[628] = i[9];
  assign o[629] = i[9];
  assign o[630] = i[9];
  assign o[631] = i[9];
  assign o[632] = i[9];
  assign o[633] = i[9];
  assign o[634] = i[9];
  assign o[635] = i[9];
  assign o[636] = i[9];
  assign o[637] = i[9];
  assign o[638] = i[9];
  assign o[639] = i[9];
  assign o[512] = i[8];
  assign o[513] = i[8];
  assign o[514] = i[8];
  assign o[515] = i[8];
  assign o[516] = i[8];
  assign o[517] = i[8];
  assign o[518] = i[8];
  assign o[519] = i[8];
  assign o[520] = i[8];
  assign o[521] = i[8];
  assign o[522] = i[8];
  assign o[523] = i[8];
  assign o[524] = i[8];
  assign o[525] = i[8];
  assign o[526] = i[8];
  assign o[527] = i[8];
  assign o[528] = i[8];
  assign o[529] = i[8];
  assign o[530] = i[8];
  assign o[531] = i[8];
  assign o[532] = i[8];
  assign o[533] = i[8];
  assign o[534] = i[8];
  assign o[535] = i[8];
  assign o[536] = i[8];
  assign o[537] = i[8];
  assign o[538] = i[8];
  assign o[539] = i[8];
  assign o[540] = i[8];
  assign o[541] = i[8];
  assign o[542] = i[8];
  assign o[543] = i[8];
  assign o[544] = i[8];
  assign o[545] = i[8];
  assign o[546] = i[8];
  assign o[547] = i[8];
  assign o[548] = i[8];
  assign o[549] = i[8];
  assign o[550] = i[8];
  assign o[551] = i[8];
  assign o[552] = i[8];
  assign o[553] = i[8];
  assign o[554] = i[8];
  assign o[555] = i[8];
  assign o[556] = i[8];
  assign o[557] = i[8];
  assign o[558] = i[8];
  assign o[559] = i[8];
  assign o[560] = i[8];
  assign o[561] = i[8];
  assign o[562] = i[8];
  assign o[563] = i[8];
  assign o[564] = i[8];
  assign o[565] = i[8];
  assign o[566] = i[8];
  assign o[567] = i[8];
  assign o[568] = i[8];
  assign o[569] = i[8];
  assign o[570] = i[8];
  assign o[571] = i[8];
  assign o[572] = i[8];
  assign o[573] = i[8];
  assign o[574] = i[8];
  assign o[575] = i[8];
  assign o[448] = i[7];
  assign o[449] = i[7];
  assign o[450] = i[7];
  assign o[451] = i[7];
  assign o[452] = i[7];
  assign o[453] = i[7];
  assign o[454] = i[7];
  assign o[455] = i[7];
  assign o[456] = i[7];
  assign o[457] = i[7];
  assign o[458] = i[7];
  assign o[459] = i[7];
  assign o[460] = i[7];
  assign o[461] = i[7];
  assign o[462] = i[7];
  assign o[463] = i[7];
  assign o[464] = i[7];
  assign o[465] = i[7];
  assign o[466] = i[7];
  assign o[467] = i[7];
  assign o[468] = i[7];
  assign o[469] = i[7];
  assign o[470] = i[7];
  assign o[471] = i[7];
  assign o[472] = i[7];
  assign o[473] = i[7];
  assign o[474] = i[7];
  assign o[475] = i[7];
  assign o[476] = i[7];
  assign o[477] = i[7];
  assign o[478] = i[7];
  assign o[479] = i[7];
  assign o[480] = i[7];
  assign o[481] = i[7];
  assign o[482] = i[7];
  assign o[483] = i[7];
  assign o[484] = i[7];
  assign o[485] = i[7];
  assign o[486] = i[7];
  assign o[487] = i[7];
  assign o[488] = i[7];
  assign o[489] = i[7];
  assign o[490] = i[7];
  assign o[491] = i[7];
  assign o[492] = i[7];
  assign o[493] = i[7];
  assign o[494] = i[7];
  assign o[495] = i[7];
  assign o[496] = i[7];
  assign o[497] = i[7];
  assign o[498] = i[7];
  assign o[499] = i[7];
  assign o[500] = i[7];
  assign o[501] = i[7];
  assign o[502] = i[7];
  assign o[503] = i[7];
  assign o[504] = i[7];
  assign o[505] = i[7];
  assign o[506] = i[7];
  assign o[507] = i[7];
  assign o[508] = i[7];
  assign o[509] = i[7];
  assign o[510] = i[7];
  assign o[511] = i[7];
  assign o[384] = i[6];
  assign o[385] = i[6];
  assign o[386] = i[6];
  assign o[387] = i[6];
  assign o[388] = i[6];
  assign o[389] = i[6];
  assign o[390] = i[6];
  assign o[391] = i[6];
  assign o[392] = i[6];
  assign o[393] = i[6];
  assign o[394] = i[6];
  assign o[395] = i[6];
  assign o[396] = i[6];
  assign o[397] = i[6];
  assign o[398] = i[6];
  assign o[399] = i[6];
  assign o[400] = i[6];
  assign o[401] = i[6];
  assign o[402] = i[6];
  assign o[403] = i[6];
  assign o[404] = i[6];
  assign o[405] = i[6];
  assign o[406] = i[6];
  assign o[407] = i[6];
  assign o[408] = i[6];
  assign o[409] = i[6];
  assign o[410] = i[6];
  assign o[411] = i[6];
  assign o[412] = i[6];
  assign o[413] = i[6];
  assign o[414] = i[6];
  assign o[415] = i[6];
  assign o[416] = i[6];
  assign o[417] = i[6];
  assign o[418] = i[6];
  assign o[419] = i[6];
  assign o[420] = i[6];
  assign o[421] = i[6];
  assign o[422] = i[6];
  assign o[423] = i[6];
  assign o[424] = i[6];
  assign o[425] = i[6];
  assign o[426] = i[6];
  assign o[427] = i[6];
  assign o[428] = i[6];
  assign o[429] = i[6];
  assign o[430] = i[6];
  assign o[431] = i[6];
  assign o[432] = i[6];
  assign o[433] = i[6];
  assign o[434] = i[6];
  assign o[435] = i[6];
  assign o[436] = i[6];
  assign o[437] = i[6];
  assign o[438] = i[6];
  assign o[439] = i[6];
  assign o[440] = i[6];
  assign o[441] = i[6];
  assign o[442] = i[6];
  assign o[443] = i[6];
  assign o[444] = i[6];
  assign o[445] = i[6];
  assign o[446] = i[6];
  assign o[447] = i[6];
  assign o[320] = i[5];
  assign o[321] = i[5];
  assign o[322] = i[5];
  assign o[323] = i[5];
  assign o[324] = i[5];
  assign o[325] = i[5];
  assign o[326] = i[5];
  assign o[327] = i[5];
  assign o[328] = i[5];
  assign o[329] = i[5];
  assign o[330] = i[5];
  assign o[331] = i[5];
  assign o[332] = i[5];
  assign o[333] = i[5];
  assign o[334] = i[5];
  assign o[335] = i[5];
  assign o[336] = i[5];
  assign o[337] = i[5];
  assign o[338] = i[5];
  assign o[339] = i[5];
  assign o[340] = i[5];
  assign o[341] = i[5];
  assign o[342] = i[5];
  assign o[343] = i[5];
  assign o[344] = i[5];
  assign o[345] = i[5];
  assign o[346] = i[5];
  assign o[347] = i[5];
  assign o[348] = i[5];
  assign o[349] = i[5];
  assign o[350] = i[5];
  assign o[351] = i[5];
  assign o[352] = i[5];
  assign o[353] = i[5];
  assign o[354] = i[5];
  assign o[355] = i[5];
  assign o[356] = i[5];
  assign o[357] = i[5];
  assign o[358] = i[5];
  assign o[359] = i[5];
  assign o[360] = i[5];
  assign o[361] = i[5];
  assign o[362] = i[5];
  assign o[363] = i[5];
  assign o[364] = i[5];
  assign o[365] = i[5];
  assign o[366] = i[5];
  assign o[367] = i[5];
  assign o[368] = i[5];
  assign o[369] = i[5];
  assign o[370] = i[5];
  assign o[371] = i[5];
  assign o[372] = i[5];
  assign o[373] = i[5];
  assign o[374] = i[5];
  assign o[375] = i[5];
  assign o[376] = i[5];
  assign o[377] = i[5];
  assign o[378] = i[5];
  assign o[379] = i[5];
  assign o[380] = i[5];
  assign o[381] = i[5];
  assign o[382] = i[5];
  assign o[383] = i[5];
  assign o[256] = i[4];
  assign o[257] = i[4];
  assign o[258] = i[4];
  assign o[259] = i[4];
  assign o[260] = i[4];
  assign o[261] = i[4];
  assign o[262] = i[4];
  assign o[263] = i[4];
  assign o[264] = i[4];
  assign o[265] = i[4];
  assign o[266] = i[4];
  assign o[267] = i[4];
  assign o[268] = i[4];
  assign o[269] = i[4];
  assign o[270] = i[4];
  assign o[271] = i[4];
  assign o[272] = i[4];
  assign o[273] = i[4];
  assign o[274] = i[4];
  assign o[275] = i[4];
  assign o[276] = i[4];
  assign o[277] = i[4];
  assign o[278] = i[4];
  assign o[279] = i[4];
  assign o[280] = i[4];
  assign o[281] = i[4];
  assign o[282] = i[4];
  assign o[283] = i[4];
  assign o[284] = i[4];
  assign o[285] = i[4];
  assign o[286] = i[4];
  assign o[287] = i[4];
  assign o[288] = i[4];
  assign o[289] = i[4];
  assign o[290] = i[4];
  assign o[291] = i[4];
  assign o[292] = i[4];
  assign o[293] = i[4];
  assign o[294] = i[4];
  assign o[295] = i[4];
  assign o[296] = i[4];
  assign o[297] = i[4];
  assign o[298] = i[4];
  assign o[299] = i[4];
  assign o[300] = i[4];
  assign o[301] = i[4];
  assign o[302] = i[4];
  assign o[303] = i[4];
  assign o[304] = i[4];
  assign o[305] = i[4];
  assign o[306] = i[4];
  assign o[307] = i[4];
  assign o[308] = i[4];
  assign o[309] = i[4];
  assign o[310] = i[4];
  assign o[311] = i[4];
  assign o[312] = i[4];
  assign o[313] = i[4];
  assign o[314] = i[4];
  assign o[315] = i[4];
  assign o[316] = i[4];
  assign o[317] = i[4];
  assign o[318] = i[4];
  assign o[319] = i[4];
  assign o[192] = i[3];
  assign o[193] = i[3];
  assign o[194] = i[3];
  assign o[195] = i[3];
  assign o[196] = i[3];
  assign o[197] = i[3];
  assign o[198] = i[3];
  assign o[199] = i[3];
  assign o[200] = i[3];
  assign o[201] = i[3];
  assign o[202] = i[3];
  assign o[203] = i[3];
  assign o[204] = i[3];
  assign o[205] = i[3];
  assign o[206] = i[3];
  assign o[207] = i[3];
  assign o[208] = i[3];
  assign o[209] = i[3];
  assign o[210] = i[3];
  assign o[211] = i[3];
  assign o[212] = i[3];
  assign o[213] = i[3];
  assign o[214] = i[3];
  assign o[215] = i[3];
  assign o[216] = i[3];
  assign o[217] = i[3];
  assign o[218] = i[3];
  assign o[219] = i[3];
  assign o[220] = i[3];
  assign o[221] = i[3];
  assign o[222] = i[3];
  assign o[223] = i[3];
  assign o[224] = i[3];
  assign o[225] = i[3];
  assign o[226] = i[3];
  assign o[227] = i[3];
  assign o[228] = i[3];
  assign o[229] = i[3];
  assign o[230] = i[3];
  assign o[231] = i[3];
  assign o[232] = i[3];
  assign o[233] = i[3];
  assign o[234] = i[3];
  assign o[235] = i[3];
  assign o[236] = i[3];
  assign o[237] = i[3];
  assign o[238] = i[3];
  assign o[239] = i[3];
  assign o[240] = i[3];
  assign o[241] = i[3];
  assign o[242] = i[3];
  assign o[243] = i[3];
  assign o[244] = i[3];
  assign o[245] = i[3];
  assign o[246] = i[3];
  assign o[247] = i[3];
  assign o[248] = i[3];
  assign o[249] = i[3];
  assign o[250] = i[3];
  assign o[251] = i[3];
  assign o[252] = i[3];
  assign o[253] = i[3];
  assign o[254] = i[3];
  assign o[255] = i[3];
  assign o[128] = i[2];
  assign o[129] = i[2];
  assign o[130] = i[2];
  assign o[131] = i[2];
  assign o[132] = i[2];
  assign o[133] = i[2];
  assign o[134] = i[2];
  assign o[135] = i[2];
  assign o[136] = i[2];
  assign o[137] = i[2];
  assign o[138] = i[2];
  assign o[139] = i[2];
  assign o[140] = i[2];
  assign o[141] = i[2];
  assign o[142] = i[2];
  assign o[143] = i[2];
  assign o[144] = i[2];
  assign o[145] = i[2];
  assign o[146] = i[2];
  assign o[147] = i[2];
  assign o[148] = i[2];
  assign o[149] = i[2];
  assign o[150] = i[2];
  assign o[151] = i[2];
  assign o[152] = i[2];
  assign o[153] = i[2];
  assign o[154] = i[2];
  assign o[155] = i[2];
  assign o[156] = i[2];
  assign o[157] = i[2];
  assign o[158] = i[2];
  assign o[159] = i[2];
  assign o[160] = i[2];
  assign o[161] = i[2];
  assign o[162] = i[2];
  assign o[163] = i[2];
  assign o[164] = i[2];
  assign o[165] = i[2];
  assign o[166] = i[2];
  assign o[167] = i[2];
  assign o[168] = i[2];
  assign o[169] = i[2];
  assign o[170] = i[2];
  assign o[171] = i[2];
  assign o[172] = i[2];
  assign o[173] = i[2];
  assign o[174] = i[2];
  assign o[175] = i[2];
  assign o[176] = i[2];
  assign o[177] = i[2];
  assign o[178] = i[2];
  assign o[179] = i[2];
  assign o[180] = i[2];
  assign o[181] = i[2];
  assign o[182] = i[2];
  assign o[183] = i[2];
  assign o[184] = i[2];
  assign o[185] = i[2];
  assign o[186] = i[2];
  assign o[187] = i[2];
  assign o[188] = i[2];
  assign o[189] = i[2];
  assign o[190] = i[2];
  assign o[191] = i[2];
  assign o[64] = i[1];
  assign o[65] = i[1];
  assign o[66] = i[1];
  assign o[67] = i[1];
  assign o[68] = i[1];
  assign o[69] = i[1];
  assign o[70] = i[1];
  assign o[71] = i[1];
  assign o[72] = i[1];
  assign o[73] = i[1];
  assign o[74] = i[1];
  assign o[75] = i[1];
  assign o[76] = i[1];
  assign o[77] = i[1];
  assign o[78] = i[1];
  assign o[79] = i[1];
  assign o[80] = i[1];
  assign o[81] = i[1];
  assign o[82] = i[1];
  assign o[83] = i[1];
  assign o[84] = i[1];
  assign o[85] = i[1];
  assign o[86] = i[1];
  assign o[87] = i[1];
  assign o[88] = i[1];
  assign o[89] = i[1];
  assign o[90] = i[1];
  assign o[91] = i[1];
  assign o[92] = i[1];
  assign o[93] = i[1];
  assign o[94] = i[1];
  assign o[95] = i[1];
  assign o[96] = i[1];
  assign o[97] = i[1];
  assign o[98] = i[1];
  assign o[99] = i[1];
  assign o[100] = i[1];
  assign o[101] = i[1];
  assign o[102] = i[1];
  assign o[103] = i[1];
  assign o[104] = i[1];
  assign o[105] = i[1];
  assign o[106] = i[1];
  assign o[107] = i[1];
  assign o[108] = i[1];
  assign o[109] = i[1];
  assign o[110] = i[1];
  assign o[111] = i[1];
  assign o[112] = i[1];
  assign o[113] = i[1];
  assign o[114] = i[1];
  assign o[115] = i[1];
  assign o[116] = i[1];
  assign o[117] = i[1];
  assign o[118] = i[1];
  assign o[119] = i[1];
  assign o[120] = i[1];
  assign o[121] = i[1];
  assign o[122] = i[1];
  assign o[123] = i[1];
  assign o[124] = i[1];
  assign o[125] = i[1];
  assign o[126] = i[1];
  assign o[127] = i[1];
  assign o[0] = i[0];
  assign o[1] = i[0];
  assign o[2] = i[0];
  assign o[3] = i[0];
  assign o[4] = i[0];
  assign o[5] = i[0];
  assign o[6] = i[0];
  assign o[7] = i[0];
  assign o[8] = i[0];
  assign o[9] = i[0];
  assign o[10] = i[0];
  assign o[11] = i[0];
  assign o[12] = i[0];
  assign o[13] = i[0];
  assign o[14] = i[0];
  assign o[15] = i[0];
  assign o[16] = i[0];
  assign o[17] = i[0];
  assign o[18] = i[0];
  assign o[19] = i[0];
  assign o[20] = i[0];
  assign o[21] = i[0];
  assign o[22] = i[0];
  assign o[23] = i[0];
  assign o[24] = i[0];
  assign o[25] = i[0];
  assign o[26] = i[0];
  assign o[27] = i[0];
  assign o[28] = i[0];
  assign o[29] = i[0];
  assign o[30] = i[0];
  assign o[31] = i[0];
  assign o[32] = i[0];
  assign o[33] = i[0];
  assign o[34] = i[0];
  assign o[35] = i[0];
  assign o[36] = i[0];
  assign o[37] = i[0];
  assign o[38] = i[0];
  assign o[39] = i[0];
  assign o[40] = i[0];
  assign o[41] = i[0];
  assign o[42] = i[0];
  assign o[43] = i[0];
  assign o[44] = i[0];
  assign o[45] = i[0];
  assign o[46] = i[0];
  assign o[47] = i[0];
  assign o[48] = i[0];
  assign o[49] = i[0];
  assign o[50] = i[0];
  assign o[51] = i[0];
  assign o[52] = i[0];
  assign o[53] = i[0];
  assign o[54] = i[0];
  assign o[55] = i[0];
  assign o[56] = i[0];
  assign o[57] = i[0];
  assign o[58] = i[0];
  assign o[59] = i[0];
  assign o[60] = i[0];
  assign o[61] = i[0];
  assign o[62] = i[0];
  assign o[63] = i[0];

endmodule

