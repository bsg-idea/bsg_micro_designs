

module top
(
  i,
  o
);

  input [31:0] i;
  output [2047:0] o;

  bsg_expand_bitmask
  wrapper
  (
    .i(i),
    .o(o)
  );


endmodule



module bsg_expand_bitmask
(
  i,
  o
);

  input [31:0] i;
  output [2047:0] o;
  wire [2047:0] o;
  wire o_2047_,o_1983_,o_1919_,o_1855_,o_1791_,o_1727_,o_1663_,o_1599_,o_1535_,o_1471_,
  o_1407_,o_1343_,o_1279_,o_1215_,o_1151_,o_1087_,o_1023_,o_959_,o_895_,o_831_,
  o_767_,o_703_,o_639_,o_575_,o_511_,o_447_,o_383_,o_319_,o_255_,o_191_,o_127_,o_63_;
  assign o_2047_ = i[31];
  assign o[1984] = o_2047_;
  assign o[1985] = o_2047_;
  assign o[1986] = o_2047_;
  assign o[1987] = o_2047_;
  assign o[1988] = o_2047_;
  assign o[1989] = o_2047_;
  assign o[1990] = o_2047_;
  assign o[1991] = o_2047_;
  assign o[1992] = o_2047_;
  assign o[1993] = o_2047_;
  assign o[1994] = o_2047_;
  assign o[1995] = o_2047_;
  assign o[1996] = o_2047_;
  assign o[1997] = o_2047_;
  assign o[1998] = o_2047_;
  assign o[1999] = o_2047_;
  assign o[2000] = o_2047_;
  assign o[2001] = o_2047_;
  assign o[2002] = o_2047_;
  assign o[2003] = o_2047_;
  assign o[2004] = o_2047_;
  assign o[2005] = o_2047_;
  assign o[2006] = o_2047_;
  assign o[2007] = o_2047_;
  assign o[2008] = o_2047_;
  assign o[2009] = o_2047_;
  assign o[2010] = o_2047_;
  assign o[2011] = o_2047_;
  assign o[2012] = o_2047_;
  assign o[2013] = o_2047_;
  assign o[2014] = o_2047_;
  assign o[2015] = o_2047_;
  assign o[2016] = o_2047_;
  assign o[2017] = o_2047_;
  assign o[2018] = o_2047_;
  assign o[2019] = o_2047_;
  assign o[2020] = o_2047_;
  assign o[2021] = o_2047_;
  assign o[2022] = o_2047_;
  assign o[2023] = o_2047_;
  assign o[2024] = o_2047_;
  assign o[2025] = o_2047_;
  assign o[2026] = o_2047_;
  assign o[2027] = o_2047_;
  assign o[2028] = o_2047_;
  assign o[2029] = o_2047_;
  assign o[2030] = o_2047_;
  assign o[2031] = o_2047_;
  assign o[2032] = o_2047_;
  assign o[2033] = o_2047_;
  assign o[2034] = o_2047_;
  assign o[2035] = o_2047_;
  assign o[2036] = o_2047_;
  assign o[2037] = o_2047_;
  assign o[2038] = o_2047_;
  assign o[2039] = o_2047_;
  assign o[2040] = o_2047_;
  assign o[2041] = o_2047_;
  assign o[2042] = o_2047_;
  assign o[2043] = o_2047_;
  assign o[2044] = o_2047_;
  assign o[2045] = o_2047_;
  assign o[2046] = o_2047_;
  assign o[2047] = o_2047_;
  assign o_1983_ = i[30];
  assign o[1920] = o_1983_;
  assign o[1921] = o_1983_;
  assign o[1922] = o_1983_;
  assign o[1923] = o_1983_;
  assign o[1924] = o_1983_;
  assign o[1925] = o_1983_;
  assign o[1926] = o_1983_;
  assign o[1927] = o_1983_;
  assign o[1928] = o_1983_;
  assign o[1929] = o_1983_;
  assign o[1930] = o_1983_;
  assign o[1931] = o_1983_;
  assign o[1932] = o_1983_;
  assign o[1933] = o_1983_;
  assign o[1934] = o_1983_;
  assign o[1935] = o_1983_;
  assign o[1936] = o_1983_;
  assign o[1937] = o_1983_;
  assign o[1938] = o_1983_;
  assign o[1939] = o_1983_;
  assign o[1940] = o_1983_;
  assign o[1941] = o_1983_;
  assign o[1942] = o_1983_;
  assign o[1943] = o_1983_;
  assign o[1944] = o_1983_;
  assign o[1945] = o_1983_;
  assign o[1946] = o_1983_;
  assign o[1947] = o_1983_;
  assign o[1948] = o_1983_;
  assign o[1949] = o_1983_;
  assign o[1950] = o_1983_;
  assign o[1951] = o_1983_;
  assign o[1952] = o_1983_;
  assign o[1953] = o_1983_;
  assign o[1954] = o_1983_;
  assign o[1955] = o_1983_;
  assign o[1956] = o_1983_;
  assign o[1957] = o_1983_;
  assign o[1958] = o_1983_;
  assign o[1959] = o_1983_;
  assign o[1960] = o_1983_;
  assign o[1961] = o_1983_;
  assign o[1962] = o_1983_;
  assign o[1963] = o_1983_;
  assign o[1964] = o_1983_;
  assign o[1965] = o_1983_;
  assign o[1966] = o_1983_;
  assign o[1967] = o_1983_;
  assign o[1968] = o_1983_;
  assign o[1969] = o_1983_;
  assign o[1970] = o_1983_;
  assign o[1971] = o_1983_;
  assign o[1972] = o_1983_;
  assign o[1973] = o_1983_;
  assign o[1974] = o_1983_;
  assign o[1975] = o_1983_;
  assign o[1976] = o_1983_;
  assign o[1977] = o_1983_;
  assign o[1978] = o_1983_;
  assign o[1979] = o_1983_;
  assign o[1980] = o_1983_;
  assign o[1981] = o_1983_;
  assign o[1982] = o_1983_;
  assign o[1983] = o_1983_;
  assign o_1919_ = i[29];
  assign o[1856] = o_1919_;
  assign o[1857] = o_1919_;
  assign o[1858] = o_1919_;
  assign o[1859] = o_1919_;
  assign o[1860] = o_1919_;
  assign o[1861] = o_1919_;
  assign o[1862] = o_1919_;
  assign o[1863] = o_1919_;
  assign o[1864] = o_1919_;
  assign o[1865] = o_1919_;
  assign o[1866] = o_1919_;
  assign o[1867] = o_1919_;
  assign o[1868] = o_1919_;
  assign o[1869] = o_1919_;
  assign o[1870] = o_1919_;
  assign o[1871] = o_1919_;
  assign o[1872] = o_1919_;
  assign o[1873] = o_1919_;
  assign o[1874] = o_1919_;
  assign o[1875] = o_1919_;
  assign o[1876] = o_1919_;
  assign o[1877] = o_1919_;
  assign o[1878] = o_1919_;
  assign o[1879] = o_1919_;
  assign o[1880] = o_1919_;
  assign o[1881] = o_1919_;
  assign o[1882] = o_1919_;
  assign o[1883] = o_1919_;
  assign o[1884] = o_1919_;
  assign o[1885] = o_1919_;
  assign o[1886] = o_1919_;
  assign o[1887] = o_1919_;
  assign o[1888] = o_1919_;
  assign o[1889] = o_1919_;
  assign o[1890] = o_1919_;
  assign o[1891] = o_1919_;
  assign o[1892] = o_1919_;
  assign o[1893] = o_1919_;
  assign o[1894] = o_1919_;
  assign o[1895] = o_1919_;
  assign o[1896] = o_1919_;
  assign o[1897] = o_1919_;
  assign o[1898] = o_1919_;
  assign o[1899] = o_1919_;
  assign o[1900] = o_1919_;
  assign o[1901] = o_1919_;
  assign o[1902] = o_1919_;
  assign o[1903] = o_1919_;
  assign o[1904] = o_1919_;
  assign o[1905] = o_1919_;
  assign o[1906] = o_1919_;
  assign o[1907] = o_1919_;
  assign o[1908] = o_1919_;
  assign o[1909] = o_1919_;
  assign o[1910] = o_1919_;
  assign o[1911] = o_1919_;
  assign o[1912] = o_1919_;
  assign o[1913] = o_1919_;
  assign o[1914] = o_1919_;
  assign o[1915] = o_1919_;
  assign o[1916] = o_1919_;
  assign o[1917] = o_1919_;
  assign o[1918] = o_1919_;
  assign o[1919] = o_1919_;
  assign o_1855_ = i[28];
  assign o[1792] = o_1855_;
  assign o[1793] = o_1855_;
  assign o[1794] = o_1855_;
  assign o[1795] = o_1855_;
  assign o[1796] = o_1855_;
  assign o[1797] = o_1855_;
  assign o[1798] = o_1855_;
  assign o[1799] = o_1855_;
  assign o[1800] = o_1855_;
  assign o[1801] = o_1855_;
  assign o[1802] = o_1855_;
  assign o[1803] = o_1855_;
  assign o[1804] = o_1855_;
  assign o[1805] = o_1855_;
  assign o[1806] = o_1855_;
  assign o[1807] = o_1855_;
  assign o[1808] = o_1855_;
  assign o[1809] = o_1855_;
  assign o[1810] = o_1855_;
  assign o[1811] = o_1855_;
  assign o[1812] = o_1855_;
  assign o[1813] = o_1855_;
  assign o[1814] = o_1855_;
  assign o[1815] = o_1855_;
  assign o[1816] = o_1855_;
  assign o[1817] = o_1855_;
  assign o[1818] = o_1855_;
  assign o[1819] = o_1855_;
  assign o[1820] = o_1855_;
  assign o[1821] = o_1855_;
  assign o[1822] = o_1855_;
  assign o[1823] = o_1855_;
  assign o[1824] = o_1855_;
  assign o[1825] = o_1855_;
  assign o[1826] = o_1855_;
  assign o[1827] = o_1855_;
  assign o[1828] = o_1855_;
  assign o[1829] = o_1855_;
  assign o[1830] = o_1855_;
  assign o[1831] = o_1855_;
  assign o[1832] = o_1855_;
  assign o[1833] = o_1855_;
  assign o[1834] = o_1855_;
  assign o[1835] = o_1855_;
  assign o[1836] = o_1855_;
  assign o[1837] = o_1855_;
  assign o[1838] = o_1855_;
  assign o[1839] = o_1855_;
  assign o[1840] = o_1855_;
  assign o[1841] = o_1855_;
  assign o[1842] = o_1855_;
  assign o[1843] = o_1855_;
  assign o[1844] = o_1855_;
  assign o[1845] = o_1855_;
  assign o[1846] = o_1855_;
  assign o[1847] = o_1855_;
  assign o[1848] = o_1855_;
  assign o[1849] = o_1855_;
  assign o[1850] = o_1855_;
  assign o[1851] = o_1855_;
  assign o[1852] = o_1855_;
  assign o[1853] = o_1855_;
  assign o[1854] = o_1855_;
  assign o[1855] = o_1855_;
  assign o_1791_ = i[27];
  assign o[1728] = o_1791_;
  assign o[1729] = o_1791_;
  assign o[1730] = o_1791_;
  assign o[1731] = o_1791_;
  assign o[1732] = o_1791_;
  assign o[1733] = o_1791_;
  assign o[1734] = o_1791_;
  assign o[1735] = o_1791_;
  assign o[1736] = o_1791_;
  assign o[1737] = o_1791_;
  assign o[1738] = o_1791_;
  assign o[1739] = o_1791_;
  assign o[1740] = o_1791_;
  assign o[1741] = o_1791_;
  assign o[1742] = o_1791_;
  assign o[1743] = o_1791_;
  assign o[1744] = o_1791_;
  assign o[1745] = o_1791_;
  assign o[1746] = o_1791_;
  assign o[1747] = o_1791_;
  assign o[1748] = o_1791_;
  assign o[1749] = o_1791_;
  assign o[1750] = o_1791_;
  assign o[1751] = o_1791_;
  assign o[1752] = o_1791_;
  assign o[1753] = o_1791_;
  assign o[1754] = o_1791_;
  assign o[1755] = o_1791_;
  assign o[1756] = o_1791_;
  assign o[1757] = o_1791_;
  assign o[1758] = o_1791_;
  assign o[1759] = o_1791_;
  assign o[1760] = o_1791_;
  assign o[1761] = o_1791_;
  assign o[1762] = o_1791_;
  assign o[1763] = o_1791_;
  assign o[1764] = o_1791_;
  assign o[1765] = o_1791_;
  assign o[1766] = o_1791_;
  assign o[1767] = o_1791_;
  assign o[1768] = o_1791_;
  assign o[1769] = o_1791_;
  assign o[1770] = o_1791_;
  assign o[1771] = o_1791_;
  assign o[1772] = o_1791_;
  assign o[1773] = o_1791_;
  assign o[1774] = o_1791_;
  assign o[1775] = o_1791_;
  assign o[1776] = o_1791_;
  assign o[1777] = o_1791_;
  assign o[1778] = o_1791_;
  assign o[1779] = o_1791_;
  assign o[1780] = o_1791_;
  assign o[1781] = o_1791_;
  assign o[1782] = o_1791_;
  assign o[1783] = o_1791_;
  assign o[1784] = o_1791_;
  assign o[1785] = o_1791_;
  assign o[1786] = o_1791_;
  assign o[1787] = o_1791_;
  assign o[1788] = o_1791_;
  assign o[1789] = o_1791_;
  assign o[1790] = o_1791_;
  assign o[1791] = o_1791_;
  assign o_1727_ = i[26];
  assign o[1664] = o_1727_;
  assign o[1665] = o_1727_;
  assign o[1666] = o_1727_;
  assign o[1667] = o_1727_;
  assign o[1668] = o_1727_;
  assign o[1669] = o_1727_;
  assign o[1670] = o_1727_;
  assign o[1671] = o_1727_;
  assign o[1672] = o_1727_;
  assign o[1673] = o_1727_;
  assign o[1674] = o_1727_;
  assign o[1675] = o_1727_;
  assign o[1676] = o_1727_;
  assign o[1677] = o_1727_;
  assign o[1678] = o_1727_;
  assign o[1679] = o_1727_;
  assign o[1680] = o_1727_;
  assign o[1681] = o_1727_;
  assign o[1682] = o_1727_;
  assign o[1683] = o_1727_;
  assign o[1684] = o_1727_;
  assign o[1685] = o_1727_;
  assign o[1686] = o_1727_;
  assign o[1687] = o_1727_;
  assign o[1688] = o_1727_;
  assign o[1689] = o_1727_;
  assign o[1690] = o_1727_;
  assign o[1691] = o_1727_;
  assign o[1692] = o_1727_;
  assign o[1693] = o_1727_;
  assign o[1694] = o_1727_;
  assign o[1695] = o_1727_;
  assign o[1696] = o_1727_;
  assign o[1697] = o_1727_;
  assign o[1698] = o_1727_;
  assign o[1699] = o_1727_;
  assign o[1700] = o_1727_;
  assign o[1701] = o_1727_;
  assign o[1702] = o_1727_;
  assign o[1703] = o_1727_;
  assign o[1704] = o_1727_;
  assign o[1705] = o_1727_;
  assign o[1706] = o_1727_;
  assign o[1707] = o_1727_;
  assign o[1708] = o_1727_;
  assign o[1709] = o_1727_;
  assign o[1710] = o_1727_;
  assign o[1711] = o_1727_;
  assign o[1712] = o_1727_;
  assign o[1713] = o_1727_;
  assign o[1714] = o_1727_;
  assign o[1715] = o_1727_;
  assign o[1716] = o_1727_;
  assign o[1717] = o_1727_;
  assign o[1718] = o_1727_;
  assign o[1719] = o_1727_;
  assign o[1720] = o_1727_;
  assign o[1721] = o_1727_;
  assign o[1722] = o_1727_;
  assign o[1723] = o_1727_;
  assign o[1724] = o_1727_;
  assign o[1725] = o_1727_;
  assign o[1726] = o_1727_;
  assign o[1727] = o_1727_;
  assign o_1663_ = i[25];
  assign o[1600] = o_1663_;
  assign o[1601] = o_1663_;
  assign o[1602] = o_1663_;
  assign o[1603] = o_1663_;
  assign o[1604] = o_1663_;
  assign o[1605] = o_1663_;
  assign o[1606] = o_1663_;
  assign o[1607] = o_1663_;
  assign o[1608] = o_1663_;
  assign o[1609] = o_1663_;
  assign o[1610] = o_1663_;
  assign o[1611] = o_1663_;
  assign o[1612] = o_1663_;
  assign o[1613] = o_1663_;
  assign o[1614] = o_1663_;
  assign o[1615] = o_1663_;
  assign o[1616] = o_1663_;
  assign o[1617] = o_1663_;
  assign o[1618] = o_1663_;
  assign o[1619] = o_1663_;
  assign o[1620] = o_1663_;
  assign o[1621] = o_1663_;
  assign o[1622] = o_1663_;
  assign o[1623] = o_1663_;
  assign o[1624] = o_1663_;
  assign o[1625] = o_1663_;
  assign o[1626] = o_1663_;
  assign o[1627] = o_1663_;
  assign o[1628] = o_1663_;
  assign o[1629] = o_1663_;
  assign o[1630] = o_1663_;
  assign o[1631] = o_1663_;
  assign o[1632] = o_1663_;
  assign o[1633] = o_1663_;
  assign o[1634] = o_1663_;
  assign o[1635] = o_1663_;
  assign o[1636] = o_1663_;
  assign o[1637] = o_1663_;
  assign o[1638] = o_1663_;
  assign o[1639] = o_1663_;
  assign o[1640] = o_1663_;
  assign o[1641] = o_1663_;
  assign o[1642] = o_1663_;
  assign o[1643] = o_1663_;
  assign o[1644] = o_1663_;
  assign o[1645] = o_1663_;
  assign o[1646] = o_1663_;
  assign o[1647] = o_1663_;
  assign o[1648] = o_1663_;
  assign o[1649] = o_1663_;
  assign o[1650] = o_1663_;
  assign o[1651] = o_1663_;
  assign o[1652] = o_1663_;
  assign o[1653] = o_1663_;
  assign o[1654] = o_1663_;
  assign o[1655] = o_1663_;
  assign o[1656] = o_1663_;
  assign o[1657] = o_1663_;
  assign o[1658] = o_1663_;
  assign o[1659] = o_1663_;
  assign o[1660] = o_1663_;
  assign o[1661] = o_1663_;
  assign o[1662] = o_1663_;
  assign o[1663] = o_1663_;
  assign o_1599_ = i[24];
  assign o[1536] = o_1599_;
  assign o[1537] = o_1599_;
  assign o[1538] = o_1599_;
  assign o[1539] = o_1599_;
  assign o[1540] = o_1599_;
  assign o[1541] = o_1599_;
  assign o[1542] = o_1599_;
  assign o[1543] = o_1599_;
  assign o[1544] = o_1599_;
  assign o[1545] = o_1599_;
  assign o[1546] = o_1599_;
  assign o[1547] = o_1599_;
  assign o[1548] = o_1599_;
  assign o[1549] = o_1599_;
  assign o[1550] = o_1599_;
  assign o[1551] = o_1599_;
  assign o[1552] = o_1599_;
  assign o[1553] = o_1599_;
  assign o[1554] = o_1599_;
  assign o[1555] = o_1599_;
  assign o[1556] = o_1599_;
  assign o[1557] = o_1599_;
  assign o[1558] = o_1599_;
  assign o[1559] = o_1599_;
  assign o[1560] = o_1599_;
  assign o[1561] = o_1599_;
  assign o[1562] = o_1599_;
  assign o[1563] = o_1599_;
  assign o[1564] = o_1599_;
  assign o[1565] = o_1599_;
  assign o[1566] = o_1599_;
  assign o[1567] = o_1599_;
  assign o[1568] = o_1599_;
  assign o[1569] = o_1599_;
  assign o[1570] = o_1599_;
  assign o[1571] = o_1599_;
  assign o[1572] = o_1599_;
  assign o[1573] = o_1599_;
  assign o[1574] = o_1599_;
  assign o[1575] = o_1599_;
  assign o[1576] = o_1599_;
  assign o[1577] = o_1599_;
  assign o[1578] = o_1599_;
  assign o[1579] = o_1599_;
  assign o[1580] = o_1599_;
  assign o[1581] = o_1599_;
  assign o[1582] = o_1599_;
  assign o[1583] = o_1599_;
  assign o[1584] = o_1599_;
  assign o[1585] = o_1599_;
  assign o[1586] = o_1599_;
  assign o[1587] = o_1599_;
  assign o[1588] = o_1599_;
  assign o[1589] = o_1599_;
  assign o[1590] = o_1599_;
  assign o[1591] = o_1599_;
  assign o[1592] = o_1599_;
  assign o[1593] = o_1599_;
  assign o[1594] = o_1599_;
  assign o[1595] = o_1599_;
  assign o[1596] = o_1599_;
  assign o[1597] = o_1599_;
  assign o[1598] = o_1599_;
  assign o[1599] = o_1599_;
  assign o_1535_ = i[23];
  assign o[1472] = o_1535_;
  assign o[1473] = o_1535_;
  assign o[1474] = o_1535_;
  assign o[1475] = o_1535_;
  assign o[1476] = o_1535_;
  assign o[1477] = o_1535_;
  assign o[1478] = o_1535_;
  assign o[1479] = o_1535_;
  assign o[1480] = o_1535_;
  assign o[1481] = o_1535_;
  assign o[1482] = o_1535_;
  assign o[1483] = o_1535_;
  assign o[1484] = o_1535_;
  assign o[1485] = o_1535_;
  assign o[1486] = o_1535_;
  assign o[1487] = o_1535_;
  assign o[1488] = o_1535_;
  assign o[1489] = o_1535_;
  assign o[1490] = o_1535_;
  assign o[1491] = o_1535_;
  assign o[1492] = o_1535_;
  assign o[1493] = o_1535_;
  assign o[1494] = o_1535_;
  assign o[1495] = o_1535_;
  assign o[1496] = o_1535_;
  assign o[1497] = o_1535_;
  assign o[1498] = o_1535_;
  assign o[1499] = o_1535_;
  assign o[1500] = o_1535_;
  assign o[1501] = o_1535_;
  assign o[1502] = o_1535_;
  assign o[1503] = o_1535_;
  assign o[1504] = o_1535_;
  assign o[1505] = o_1535_;
  assign o[1506] = o_1535_;
  assign o[1507] = o_1535_;
  assign o[1508] = o_1535_;
  assign o[1509] = o_1535_;
  assign o[1510] = o_1535_;
  assign o[1511] = o_1535_;
  assign o[1512] = o_1535_;
  assign o[1513] = o_1535_;
  assign o[1514] = o_1535_;
  assign o[1515] = o_1535_;
  assign o[1516] = o_1535_;
  assign o[1517] = o_1535_;
  assign o[1518] = o_1535_;
  assign o[1519] = o_1535_;
  assign o[1520] = o_1535_;
  assign o[1521] = o_1535_;
  assign o[1522] = o_1535_;
  assign o[1523] = o_1535_;
  assign o[1524] = o_1535_;
  assign o[1525] = o_1535_;
  assign o[1526] = o_1535_;
  assign o[1527] = o_1535_;
  assign o[1528] = o_1535_;
  assign o[1529] = o_1535_;
  assign o[1530] = o_1535_;
  assign o[1531] = o_1535_;
  assign o[1532] = o_1535_;
  assign o[1533] = o_1535_;
  assign o[1534] = o_1535_;
  assign o[1535] = o_1535_;
  assign o_1471_ = i[22];
  assign o[1408] = o_1471_;
  assign o[1409] = o_1471_;
  assign o[1410] = o_1471_;
  assign o[1411] = o_1471_;
  assign o[1412] = o_1471_;
  assign o[1413] = o_1471_;
  assign o[1414] = o_1471_;
  assign o[1415] = o_1471_;
  assign o[1416] = o_1471_;
  assign o[1417] = o_1471_;
  assign o[1418] = o_1471_;
  assign o[1419] = o_1471_;
  assign o[1420] = o_1471_;
  assign o[1421] = o_1471_;
  assign o[1422] = o_1471_;
  assign o[1423] = o_1471_;
  assign o[1424] = o_1471_;
  assign o[1425] = o_1471_;
  assign o[1426] = o_1471_;
  assign o[1427] = o_1471_;
  assign o[1428] = o_1471_;
  assign o[1429] = o_1471_;
  assign o[1430] = o_1471_;
  assign o[1431] = o_1471_;
  assign o[1432] = o_1471_;
  assign o[1433] = o_1471_;
  assign o[1434] = o_1471_;
  assign o[1435] = o_1471_;
  assign o[1436] = o_1471_;
  assign o[1437] = o_1471_;
  assign o[1438] = o_1471_;
  assign o[1439] = o_1471_;
  assign o[1440] = o_1471_;
  assign o[1441] = o_1471_;
  assign o[1442] = o_1471_;
  assign o[1443] = o_1471_;
  assign o[1444] = o_1471_;
  assign o[1445] = o_1471_;
  assign o[1446] = o_1471_;
  assign o[1447] = o_1471_;
  assign o[1448] = o_1471_;
  assign o[1449] = o_1471_;
  assign o[1450] = o_1471_;
  assign o[1451] = o_1471_;
  assign o[1452] = o_1471_;
  assign o[1453] = o_1471_;
  assign o[1454] = o_1471_;
  assign o[1455] = o_1471_;
  assign o[1456] = o_1471_;
  assign o[1457] = o_1471_;
  assign o[1458] = o_1471_;
  assign o[1459] = o_1471_;
  assign o[1460] = o_1471_;
  assign o[1461] = o_1471_;
  assign o[1462] = o_1471_;
  assign o[1463] = o_1471_;
  assign o[1464] = o_1471_;
  assign o[1465] = o_1471_;
  assign o[1466] = o_1471_;
  assign o[1467] = o_1471_;
  assign o[1468] = o_1471_;
  assign o[1469] = o_1471_;
  assign o[1470] = o_1471_;
  assign o[1471] = o_1471_;
  assign o_1407_ = i[21];
  assign o[1344] = o_1407_;
  assign o[1345] = o_1407_;
  assign o[1346] = o_1407_;
  assign o[1347] = o_1407_;
  assign o[1348] = o_1407_;
  assign o[1349] = o_1407_;
  assign o[1350] = o_1407_;
  assign o[1351] = o_1407_;
  assign o[1352] = o_1407_;
  assign o[1353] = o_1407_;
  assign o[1354] = o_1407_;
  assign o[1355] = o_1407_;
  assign o[1356] = o_1407_;
  assign o[1357] = o_1407_;
  assign o[1358] = o_1407_;
  assign o[1359] = o_1407_;
  assign o[1360] = o_1407_;
  assign o[1361] = o_1407_;
  assign o[1362] = o_1407_;
  assign o[1363] = o_1407_;
  assign o[1364] = o_1407_;
  assign o[1365] = o_1407_;
  assign o[1366] = o_1407_;
  assign o[1367] = o_1407_;
  assign o[1368] = o_1407_;
  assign o[1369] = o_1407_;
  assign o[1370] = o_1407_;
  assign o[1371] = o_1407_;
  assign o[1372] = o_1407_;
  assign o[1373] = o_1407_;
  assign o[1374] = o_1407_;
  assign o[1375] = o_1407_;
  assign o[1376] = o_1407_;
  assign o[1377] = o_1407_;
  assign o[1378] = o_1407_;
  assign o[1379] = o_1407_;
  assign o[1380] = o_1407_;
  assign o[1381] = o_1407_;
  assign o[1382] = o_1407_;
  assign o[1383] = o_1407_;
  assign o[1384] = o_1407_;
  assign o[1385] = o_1407_;
  assign o[1386] = o_1407_;
  assign o[1387] = o_1407_;
  assign o[1388] = o_1407_;
  assign o[1389] = o_1407_;
  assign o[1390] = o_1407_;
  assign o[1391] = o_1407_;
  assign o[1392] = o_1407_;
  assign o[1393] = o_1407_;
  assign o[1394] = o_1407_;
  assign o[1395] = o_1407_;
  assign o[1396] = o_1407_;
  assign o[1397] = o_1407_;
  assign o[1398] = o_1407_;
  assign o[1399] = o_1407_;
  assign o[1400] = o_1407_;
  assign o[1401] = o_1407_;
  assign o[1402] = o_1407_;
  assign o[1403] = o_1407_;
  assign o[1404] = o_1407_;
  assign o[1405] = o_1407_;
  assign o[1406] = o_1407_;
  assign o[1407] = o_1407_;
  assign o_1343_ = i[20];
  assign o[1280] = o_1343_;
  assign o[1281] = o_1343_;
  assign o[1282] = o_1343_;
  assign o[1283] = o_1343_;
  assign o[1284] = o_1343_;
  assign o[1285] = o_1343_;
  assign o[1286] = o_1343_;
  assign o[1287] = o_1343_;
  assign o[1288] = o_1343_;
  assign o[1289] = o_1343_;
  assign o[1290] = o_1343_;
  assign o[1291] = o_1343_;
  assign o[1292] = o_1343_;
  assign o[1293] = o_1343_;
  assign o[1294] = o_1343_;
  assign o[1295] = o_1343_;
  assign o[1296] = o_1343_;
  assign o[1297] = o_1343_;
  assign o[1298] = o_1343_;
  assign o[1299] = o_1343_;
  assign o[1300] = o_1343_;
  assign o[1301] = o_1343_;
  assign o[1302] = o_1343_;
  assign o[1303] = o_1343_;
  assign o[1304] = o_1343_;
  assign o[1305] = o_1343_;
  assign o[1306] = o_1343_;
  assign o[1307] = o_1343_;
  assign o[1308] = o_1343_;
  assign o[1309] = o_1343_;
  assign o[1310] = o_1343_;
  assign o[1311] = o_1343_;
  assign o[1312] = o_1343_;
  assign o[1313] = o_1343_;
  assign o[1314] = o_1343_;
  assign o[1315] = o_1343_;
  assign o[1316] = o_1343_;
  assign o[1317] = o_1343_;
  assign o[1318] = o_1343_;
  assign o[1319] = o_1343_;
  assign o[1320] = o_1343_;
  assign o[1321] = o_1343_;
  assign o[1322] = o_1343_;
  assign o[1323] = o_1343_;
  assign o[1324] = o_1343_;
  assign o[1325] = o_1343_;
  assign o[1326] = o_1343_;
  assign o[1327] = o_1343_;
  assign o[1328] = o_1343_;
  assign o[1329] = o_1343_;
  assign o[1330] = o_1343_;
  assign o[1331] = o_1343_;
  assign o[1332] = o_1343_;
  assign o[1333] = o_1343_;
  assign o[1334] = o_1343_;
  assign o[1335] = o_1343_;
  assign o[1336] = o_1343_;
  assign o[1337] = o_1343_;
  assign o[1338] = o_1343_;
  assign o[1339] = o_1343_;
  assign o[1340] = o_1343_;
  assign o[1341] = o_1343_;
  assign o[1342] = o_1343_;
  assign o[1343] = o_1343_;
  assign o_1279_ = i[19];
  assign o[1216] = o_1279_;
  assign o[1217] = o_1279_;
  assign o[1218] = o_1279_;
  assign o[1219] = o_1279_;
  assign o[1220] = o_1279_;
  assign o[1221] = o_1279_;
  assign o[1222] = o_1279_;
  assign o[1223] = o_1279_;
  assign o[1224] = o_1279_;
  assign o[1225] = o_1279_;
  assign o[1226] = o_1279_;
  assign o[1227] = o_1279_;
  assign o[1228] = o_1279_;
  assign o[1229] = o_1279_;
  assign o[1230] = o_1279_;
  assign o[1231] = o_1279_;
  assign o[1232] = o_1279_;
  assign o[1233] = o_1279_;
  assign o[1234] = o_1279_;
  assign o[1235] = o_1279_;
  assign o[1236] = o_1279_;
  assign o[1237] = o_1279_;
  assign o[1238] = o_1279_;
  assign o[1239] = o_1279_;
  assign o[1240] = o_1279_;
  assign o[1241] = o_1279_;
  assign o[1242] = o_1279_;
  assign o[1243] = o_1279_;
  assign o[1244] = o_1279_;
  assign o[1245] = o_1279_;
  assign o[1246] = o_1279_;
  assign o[1247] = o_1279_;
  assign o[1248] = o_1279_;
  assign o[1249] = o_1279_;
  assign o[1250] = o_1279_;
  assign o[1251] = o_1279_;
  assign o[1252] = o_1279_;
  assign o[1253] = o_1279_;
  assign o[1254] = o_1279_;
  assign o[1255] = o_1279_;
  assign o[1256] = o_1279_;
  assign o[1257] = o_1279_;
  assign o[1258] = o_1279_;
  assign o[1259] = o_1279_;
  assign o[1260] = o_1279_;
  assign o[1261] = o_1279_;
  assign o[1262] = o_1279_;
  assign o[1263] = o_1279_;
  assign o[1264] = o_1279_;
  assign o[1265] = o_1279_;
  assign o[1266] = o_1279_;
  assign o[1267] = o_1279_;
  assign o[1268] = o_1279_;
  assign o[1269] = o_1279_;
  assign o[1270] = o_1279_;
  assign o[1271] = o_1279_;
  assign o[1272] = o_1279_;
  assign o[1273] = o_1279_;
  assign o[1274] = o_1279_;
  assign o[1275] = o_1279_;
  assign o[1276] = o_1279_;
  assign o[1277] = o_1279_;
  assign o[1278] = o_1279_;
  assign o[1279] = o_1279_;
  assign o_1215_ = i[18];
  assign o[1152] = o_1215_;
  assign o[1153] = o_1215_;
  assign o[1154] = o_1215_;
  assign o[1155] = o_1215_;
  assign o[1156] = o_1215_;
  assign o[1157] = o_1215_;
  assign o[1158] = o_1215_;
  assign o[1159] = o_1215_;
  assign o[1160] = o_1215_;
  assign o[1161] = o_1215_;
  assign o[1162] = o_1215_;
  assign o[1163] = o_1215_;
  assign o[1164] = o_1215_;
  assign o[1165] = o_1215_;
  assign o[1166] = o_1215_;
  assign o[1167] = o_1215_;
  assign o[1168] = o_1215_;
  assign o[1169] = o_1215_;
  assign o[1170] = o_1215_;
  assign o[1171] = o_1215_;
  assign o[1172] = o_1215_;
  assign o[1173] = o_1215_;
  assign o[1174] = o_1215_;
  assign o[1175] = o_1215_;
  assign o[1176] = o_1215_;
  assign o[1177] = o_1215_;
  assign o[1178] = o_1215_;
  assign o[1179] = o_1215_;
  assign o[1180] = o_1215_;
  assign o[1181] = o_1215_;
  assign o[1182] = o_1215_;
  assign o[1183] = o_1215_;
  assign o[1184] = o_1215_;
  assign o[1185] = o_1215_;
  assign o[1186] = o_1215_;
  assign o[1187] = o_1215_;
  assign o[1188] = o_1215_;
  assign o[1189] = o_1215_;
  assign o[1190] = o_1215_;
  assign o[1191] = o_1215_;
  assign o[1192] = o_1215_;
  assign o[1193] = o_1215_;
  assign o[1194] = o_1215_;
  assign o[1195] = o_1215_;
  assign o[1196] = o_1215_;
  assign o[1197] = o_1215_;
  assign o[1198] = o_1215_;
  assign o[1199] = o_1215_;
  assign o[1200] = o_1215_;
  assign o[1201] = o_1215_;
  assign o[1202] = o_1215_;
  assign o[1203] = o_1215_;
  assign o[1204] = o_1215_;
  assign o[1205] = o_1215_;
  assign o[1206] = o_1215_;
  assign o[1207] = o_1215_;
  assign o[1208] = o_1215_;
  assign o[1209] = o_1215_;
  assign o[1210] = o_1215_;
  assign o[1211] = o_1215_;
  assign o[1212] = o_1215_;
  assign o[1213] = o_1215_;
  assign o[1214] = o_1215_;
  assign o[1215] = o_1215_;
  assign o_1151_ = i[17];
  assign o[1088] = o_1151_;
  assign o[1089] = o_1151_;
  assign o[1090] = o_1151_;
  assign o[1091] = o_1151_;
  assign o[1092] = o_1151_;
  assign o[1093] = o_1151_;
  assign o[1094] = o_1151_;
  assign o[1095] = o_1151_;
  assign o[1096] = o_1151_;
  assign o[1097] = o_1151_;
  assign o[1098] = o_1151_;
  assign o[1099] = o_1151_;
  assign o[1100] = o_1151_;
  assign o[1101] = o_1151_;
  assign o[1102] = o_1151_;
  assign o[1103] = o_1151_;
  assign o[1104] = o_1151_;
  assign o[1105] = o_1151_;
  assign o[1106] = o_1151_;
  assign o[1107] = o_1151_;
  assign o[1108] = o_1151_;
  assign o[1109] = o_1151_;
  assign o[1110] = o_1151_;
  assign o[1111] = o_1151_;
  assign o[1112] = o_1151_;
  assign o[1113] = o_1151_;
  assign o[1114] = o_1151_;
  assign o[1115] = o_1151_;
  assign o[1116] = o_1151_;
  assign o[1117] = o_1151_;
  assign o[1118] = o_1151_;
  assign o[1119] = o_1151_;
  assign o[1120] = o_1151_;
  assign o[1121] = o_1151_;
  assign o[1122] = o_1151_;
  assign o[1123] = o_1151_;
  assign o[1124] = o_1151_;
  assign o[1125] = o_1151_;
  assign o[1126] = o_1151_;
  assign o[1127] = o_1151_;
  assign o[1128] = o_1151_;
  assign o[1129] = o_1151_;
  assign o[1130] = o_1151_;
  assign o[1131] = o_1151_;
  assign o[1132] = o_1151_;
  assign o[1133] = o_1151_;
  assign o[1134] = o_1151_;
  assign o[1135] = o_1151_;
  assign o[1136] = o_1151_;
  assign o[1137] = o_1151_;
  assign o[1138] = o_1151_;
  assign o[1139] = o_1151_;
  assign o[1140] = o_1151_;
  assign o[1141] = o_1151_;
  assign o[1142] = o_1151_;
  assign o[1143] = o_1151_;
  assign o[1144] = o_1151_;
  assign o[1145] = o_1151_;
  assign o[1146] = o_1151_;
  assign o[1147] = o_1151_;
  assign o[1148] = o_1151_;
  assign o[1149] = o_1151_;
  assign o[1150] = o_1151_;
  assign o[1151] = o_1151_;
  assign o_1087_ = i[16];
  assign o[1024] = o_1087_;
  assign o[1025] = o_1087_;
  assign o[1026] = o_1087_;
  assign o[1027] = o_1087_;
  assign o[1028] = o_1087_;
  assign o[1029] = o_1087_;
  assign o[1030] = o_1087_;
  assign o[1031] = o_1087_;
  assign o[1032] = o_1087_;
  assign o[1033] = o_1087_;
  assign o[1034] = o_1087_;
  assign o[1035] = o_1087_;
  assign o[1036] = o_1087_;
  assign o[1037] = o_1087_;
  assign o[1038] = o_1087_;
  assign o[1039] = o_1087_;
  assign o[1040] = o_1087_;
  assign o[1041] = o_1087_;
  assign o[1042] = o_1087_;
  assign o[1043] = o_1087_;
  assign o[1044] = o_1087_;
  assign o[1045] = o_1087_;
  assign o[1046] = o_1087_;
  assign o[1047] = o_1087_;
  assign o[1048] = o_1087_;
  assign o[1049] = o_1087_;
  assign o[1050] = o_1087_;
  assign o[1051] = o_1087_;
  assign o[1052] = o_1087_;
  assign o[1053] = o_1087_;
  assign o[1054] = o_1087_;
  assign o[1055] = o_1087_;
  assign o[1056] = o_1087_;
  assign o[1057] = o_1087_;
  assign o[1058] = o_1087_;
  assign o[1059] = o_1087_;
  assign o[1060] = o_1087_;
  assign o[1061] = o_1087_;
  assign o[1062] = o_1087_;
  assign o[1063] = o_1087_;
  assign o[1064] = o_1087_;
  assign o[1065] = o_1087_;
  assign o[1066] = o_1087_;
  assign o[1067] = o_1087_;
  assign o[1068] = o_1087_;
  assign o[1069] = o_1087_;
  assign o[1070] = o_1087_;
  assign o[1071] = o_1087_;
  assign o[1072] = o_1087_;
  assign o[1073] = o_1087_;
  assign o[1074] = o_1087_;
  assign o[1075] = o_1087_;
  assign o[1076] = o_1087_;
  assign o[1077] = o_1087_;
  assign o[1078] = o_1087_;
  assign o[1079] = o_1087_;
  assign o[1080] = o_1087_;
  assign o[1081] = o_1087_;
  assign o[1082] = o_1087_;
  assign o[1083] = o_1087_;
  assign o[1084] = o_1087_;
  assign o[1085] = o_1087_;
  assign o[1086] = o_1087_;
  assign o[1087] = o_1087_;
  assign o_1023_ = i[15];
  assign o[960] = o_1023_;
  assign o[961] = o_1023_;
  assign o[962] = o_1023_;
  assign o[963] = o_1023_;
  assign o[964] = o_1023_;
  assign o[965] = o_1023_;
  assign o[966] = o_1023_;
  assign o[967] = o_1023_;
  assign o[968] = o_1023_;
  assign o[969] = o_1023_;
  assign o[970] = o_1023_;
  assign o[971] = o_1023_;
  assign o[972] = o_1023_;
  assign o[973] = o_1023_;
  assign o[974] = o_1023_;
  assign o[975] = o_1023_;
  assign o[976] = o_1023_;
  assign o[977] = o_1023_;
  assign o[978] = o_1023_;
  assign o[979] = o_1023_;
  assign o[980] = o_1023_;
  assign o[981] = o_1023_;
  assign o[982] = o_1023_;
  assign o[983] = o_1023_;
  assign o[984] = o_1023_;
  assign o[985] = o_1023_;
  assign o[986] = o_1023_;
  assign o[987] = o_1023_;
  assign o[988] = o_1023_;
  assign o[989] = o_1023_;
  assign o[990] = o_1023_;
  assign o[991] = o_1023_;
  assign o[992] = o_1023_;
  assign o[993] = o_1023_;
  assign o[994] = o_1023_;
  assign o[995] = o_1023_;
  assign o[996] = o_1023_;
  assign o[997] = o_1023_;
  assign o[998] = o_1023_;
  assign o[999] = o_1023_;
  assign o[1000] = o_1023_;
  assign o[1001] = o_1023_;
  assign o[1002] = o_1023_;
  assign o[1003] = o_1023_;
  assign o[1004] = o_1023_;
  assign o[1005] = o_1023_;
  assign o[1006] = o_1023_;
  assign o[1007] = o_1023_;
  assign o[1008] = o_1023_;
  assign o[1009] = o_1023_;
  assign o[1010] = o_1023_;
  assign o[1011] = o_1023_;
  assign o[1012] = o_1023_;
  assign o[1013] = o_1023_;
  assign o[1014] = o_1023_;
  assign o[1015] = o_1023_;
  assign o[1016] = o_1023_;
  assign o[1017] = o_1023_;
  assign o[1018] = o_1023_;
  assign o[1019] = o_1023_;
  assign o[1020] = o_1023_;
  assign o[1021] = o_1023_;
  assign o[1022] = o_1023_;
  assign o[1023] = o_1023_;
  assign o_959_ = i[14];
  assign o[896] = o_959_;
  assign o[897] = o_959_;
  assign o[898] = o_959_;
  assign o[899] = o_959_;
  assign o[900] = o_959_;
  assign o[901] = o_959_;
  assign o[902] = o_959_;
  assign o[903] = o_959_;
  assign o[904] = o_959_;
  assign o[905] = o_959_;
  assign o[906] = o_959_;
  assign o[907] = o_959_;
  assign o[908] = o_959_;
  assign o[909] = o_959_;
  assign o[910] = o_959_;
  assign o[911] = o_959_;
  assign o[912] = o_959_;
  assign o[913] = o_959_;
  assign o[914] = o_959_;
  assign o[915] = o_959_;
  assign o[916] = o_959_;
  assign o[917] = o_959_;
  assign o[918] = o_959_;
  assign o[919] = o_959_;
  assign o[920] = o_959_;
  assign o[921] = o_959_;
  assign o[922] = o_959_;
  assign o[923] = o_959_;
  assign o[924] = o_959_;
  assign o[925] = o_959_;
  assign o[926] = o_959_;
  assign o[927] = o_959_;
  assign o[928] = o_959_;
  assign o[929] = o_959_;
  assign o[930] = o_959_;
  assign o[931] = o_959_;
  assign o[932] = o_959_;
  assign o[933] = o_959_;
  assign o[934] = o_959_;
  assign o[935] = o_959_;
  assign o[936] = o_959_;
  assign o[937] = o_959_;
  assign o[938] = o_959_;
  assign o[939] = o_959_;
  assign o[940] = o_959_;
  assign o[941] = o_959_;
  assign o[942] = o_959_;
  assign o[943] = o_959_;
  assign o[944] = o_959_;
  assign o[945] = o_959_;
  assign o[946] = o_959_;
  assign o[947] = o_959_;
  assign o[948] = o_959_;
  assign o[949] = o_959_;
  assign o[950] = o_959_;
  assign o[951] = o_959_;
  assign o[952] = o_959_;
  assign o[953] = o_959_;
  assign o[954] = o_959_;
  assign o[955] = o_959_;
  assign o[956] = o_959_;
  assign o[957] = o_959_;
  assign o[958] = o_959_;
  assign o[959] = o_959_;
  assign o_895_ = i[13];
  assign o[832] = o_895_;
  assign o[833] = o_895_;
  assign o[834] = o_895_;
  assign o[835] = o_895_;
  assign o[836] = o_895_;
  assign o[837] = o_895_;
  assign o[838] = o_895_;
  assign o[839] = o_895_;
  assign o[840] = o_895_;
  assign o[841] = o_895_;
  assign o[842] = o_895_;
  assign o[843] = o_895_;
  assign o[844] = o_895_;
  assign o[845] = o_895_;
  assign o[846] = o_895_;
  assign o[847] = o_895_;
  assign o[848] = o_895_;
  assign o[849] = o_895_;
  assign o[850] = o_895_;
  assign o[851] = o_895_;
  assign o[852] = o_895_;
  assign o[853] = o_895_;
  assign o[854] = o_895_;
  assign o[855] = o_895_;
  assign o[856] = o_895_;
  assign o[857] = o_895_;
  assign o[858] = o_895_;
  assign o[859] = o_895_;
  assign o[860] = o_895_;
  assign o[861] = o_895_;
  assign o[862] = o_895_;
  assign o[863] = o_895_;
  assign o[864] = o_895_;
  assign o[865] = o_895_;
  assign o[866] = o_895_;
  assign o[867] = o_895_;
  assign o[868] = o_895_;
  assign o[869] = o_895_;
  assign o[870] = o_895_;
  assign o[871] = o_895_;
  assign o[872] = o_895_;
  assign o[873] = o_895_;
  assign o[874] = o_895_;
  assign o[875] = o_895_;
  assign o[876] = o_895_;
  assign o[877] = o_895_;
  assign o[878] = o_895_;
  assign o[879] = o_895_;
  assign o[880] = o_895_;
  assign o[881] = o_895_;
  assign o[882] = o_895_;
  assign o[883] = o_895_;
  assign o[884] = o_895_;
  assign o[885] = o_895_;
  assign o[886] = o_895_;
  assign o[887] = o_895_;
  assign o[888] = o_895_;
  assign o[889] = o_895_;
  assign o[890] = o_895_;
  assign o[891] = o_895_;
  assign o[892] = o_895_;
  assign o[893] = o_895_;
  assign o[894] = o_895_;
  assign o[895] = o_895_;
  assign o_831_ = i[12];
  assign o[768] = o_831_;
  assign o[769] = o_831_;
  assign o[770] = o_831_;
  assign o[771] = o_831_;
  assign o[772] = o_831_;
  assign o[773] = o_831_;
  assign o[774] = o_831_;
  assign o[775] = o_831_;
  assign o[776] = o_831_;
  assign o[777] = o_831_;
  assign o[778] = o_831_;
  assign o[779] = o_831_;
  assign o[780] = o_831_;
  assign o[781] = o_831_;
  assign o[782] = o_831_;
  assign o[783] = o_831_;
  assign o[784] = o_831_;
  assign o[785] = o_831_;
  assign o[786] = o_831_;
  assign o[787] = o_831_;
  assign o[788] = o_831_;
  assign o[789] = o_831_;
  assign o[790] = o_831_;
  assign o[791] = o_831_;
  assign o[792] = o_831_;
  assign o[793] = o_831_;
  assign o[794] = o_831_;
  assign o[795] = o_831_;
  assign o[796] = o_831_;
  assign o[797] = o_831_;
  assign o[798] = o_831_;
  assign o[799] = o_831_;
  assign o[800] = o_831_;
  assign o[801] = o_831_;
  assign o[802] = o_831_;
  assign o[803] = o_831_;
  assign o[804] = o_831_;
  assign o[805] = o_831_;
  assign o[806] = o_831_;
  assign o[807] = o_831_;
  assign o[808] = o_831_;
  assign o[809] = o_831_;
  assign o[810] = o_831_;
  assign o[811] = o_831_;
  assign o[812] = o_831_;
  assign o[813] = o_831_;
  assign o[814] = o_831_;
  assign o[815] = o_831_;
  assign o[816] = o_831_;
  assign o[817] = o_831_;
  assign o[818] = o_831_;
  assign o[819] = o_831_;
  assign o[820] = o_831_;
  assign o[821] = o_831_;
  assign o[822] = o_831_;
  assign o[823] = o_831_;
  assign o[824] = o_831_;
  assign o[825] = o_831_;
  assign o[826] = o_831_;
  assign o[827] = o_831_;
  assign o[828] = o_831_;
  assign o[829] = o_831_;
  assign o[830] = o_831_;
  assign o[831] = o_831_;
  assign o_767_ = i[11];
  assign o[704] = o_767_;
  assign o[705] = o_767_;
  assign o[706] = o_767_;
  assign o[707] = o_767_;
  assign o[708] = o_767_;
  assign o[709] = o_767_;
  assign o[710] = o_767_;
  assign o[711] = o_767_;
  assign o[712] = o_767_;
  assign o[713] = o_767_;
  assign o[714] = o_767_;
  assign o[715] = o_767_;
  assign o[716] = o_767_;
  assign o[717] = o_767_;
  assign o[718] = o_767_;
  assign o[719] = o_767_;
  assign o[720] = o_767_;
  assign o[721] = o_767_;
  assign o[722] = o_767_;
  assign o[723] = o_767_;
  assign o[724] = o_767_;
  assign o[725] = o_767_;
  assign o[726] = o_767_;
  assign o[727] = o_767_;
  assign o[728] = o_767_;
  assign o[729] = o_767_;
  assign o[730] = o_767_;
  assign o[731] = o_767_;
  assign o[732] = o_767_;
  assign o[733] = o_767_;
  assign o[734] = o_767_;
  assign o[735] = o_767_;
  assign o[736] = o_767_;
  assign o[737] = o_767_;
  assign o[738] = o_767_;
  assign o[739] = o_767_;
  assign o[740] = o_767_;
  assign o[741] = o_767_;
  assign o[742] = o_767_;
  assign o[743] = o_767_;
  assign o[744] = o_767_;
  assign o[745] = o_767_;
  assign o[746] = o_767_;
  assign o[747] = o_767_;
  assign o[748] = o_767_;
  assign o[749] = o_767_;
  assign o[750] = o_767_;
  assign o[751] = o_767_;
  assign o[752] = o_767_;
  assign o[753] = o_767_;
  assign o[754] = o_767_;
  assign o[755] = o_767_;
  assign o[756] = o_767_;
  assign o[757] = o_767_;
  assign o[758] = o_767_;
  assign o[759] = o_767_;
  assign o[760] = o_767_;
  assign o[761] = o_767_;
  assign o[762] = o_767_;
  assign o[763] = o_767_;
  assign o[764] = o_767_;
  assign o[765] = o_767_;
  assign o[766] = o_767_;
  assign o[767] = o_767_;
  assign o_703_ = i[10];
  assign o[640] = o_703_;
  assign o[641] = o_703_;
  assign o[642] = o_703_;
  assign o[643] = o_703_;
  assign o[644] = o_703_;
  assign o[645] = o_703_;
  assign o[646] = o_703_;
  assign o[647] = o_703_;
  assign o[648] = o_703_;
  assign o[649] = o_703_;
  assign o[650] = o_703_;
  assign o[651] = o_703_;
  assign o[652] = o_703_;
  assign o[653] = o_703_;
  assign o[654] = o_703_;
  assign o[655] = o_703_;
  assign o[656] = o_703_;
  assign o[657] = o_703_;
  assign o[658] = o_703_;
  assign o[659] = o_703_;
  assign o[660] = o_703_;
  assign o[661] = o_703_;
  assign o[662] = o_703_;
  assign o[663] = o_703_;
  assign o[664] = o_703_;
  assign o[665] = o_703_;
  assign o[666] = o_703_;
  assign o[667] = o_703_;
  assign o[668] = o_703_;
  assign o[669] = o_703_;
  assign o[670] = o_703_;
  assign o[671] = o_703_;
  assign o[672] = o_703_;
  assign o[673] = o_703_;
  assign o[674] = o_703_;
  assign o[675] = o_703_;
  assign o[676] = o_703_;
  assign o[677] = o_703_;
  assign o[678] = o_703_;
  assign o[679] = o_703_;
  assign o[680] = o_703_;
  assign o[681] = o_703_;
  assign o[682] = o_703_;
  assign o[683] = o_703_;
  assign o[684] = o_703_;
  assign o[685] = o_703_;
  assign o[686] = o_703_;
  assign o[687] = o_703_;
  assign o[688] = o_703_;
  assign o[689] = o_703_;
  assign o[690] = o_703_;
  assign o[691] = o_703_;
  assign o[692] = o_703_;
  assign o[693] = o_703_;
  assign o[694] = o_703_;
  assign o[695] = o_703_;
  assign o[696] = o_703_;
  assign o[697] = o_703_;
  assign o[698] = o_703_;
  assign o[699] = o_703_;
  assign o[700] = o_703_;
  assign o[701] = o_703_;
  assign o[702] = o_703_;
  assign o[703] = o_703_;
  assign o_639_ = i[9];
  assign o[576] = o_639_;
  assign o[577] = o_639_;
  assign o[578] = o_639_;
  assign o[579] = o_639_;
  assign o[580] = o_639_;
  assign o[581] = o_639_;
  assign o[582] = o_639_;
  assign o[583] = o_639_;
  assign o[584] = o_639_;
  assign o[585] = o_639_;
  assign o[586] = o_639_;
  assign o[587] = o_639_;
  assign o[588] = o_639_;
  assign o[589] = o_639_;
  assign o[590] = o_639_;
  assign o[591] = o_639_;
  assign o[592] = o_639_;
  assign o[593] = o_639_;
  assign o[594] = o_639_;
  assign o[595] = o_639_;
  assign o[596] = o_639_;
  assign o[597] = o_639_;
  assign o[598] = o_639_;
  assign o[599] = o_639_;
  assign o[600] = o_639_;
  assign o[601] = o_639_;
  assign o[602] = o_639_;
  assign o[603] = o_639_;
  assign o[604] = o_639_;
  assign o[605] = o_639_;
  assign o[606] = o_639_;
  assign o[607] = o_639_;
  assign o[608] = o_639_;
  assign o[609] = o_639_;
  assign o[610] = o_639_;
  assign o[611] = o_639_;
  assign o[612] = o_639_;
  assign o[613] = o_639_;
  assign o[614] = o_639_;
  assign o[615] = o_639_;
  assign o[616] = o_639_;
  assign o[617] = o_639_;
  assign o[618] = o_639_;
  assign o[619] = o_639_;
  assign o[620] = o_639_;
  assign o[621] = o_639_;
  assign o[622] = o_639_;
  assign o[623] = o_639_;
  assign o[624] = o_639_;
  assign o[625] = o_639_;
  assign o[626] = o_639_;
  assign o[627] = o_639_;
  assign o[628] = o_639_;
  assign o[629] = o_639_;
  assign o[630] = o_639_;
  assign o[631] = o_639_;
  assign o[632] = o_639_;
  assign o[633] = o_639_;
  assign o[634] = o_639_;
  assign o[635] = o_639_;
  assign o[636] = o_639_;
  assign o[637] = o_639_;
  assign o[638] = o_639_;
  assign o[639] = o_639_;
  assign o_575_ = i[8];
  assign o[512] = o_575_;
  assign o[513] = o_575_;
  assign o[514] = o_575_;
  assign o[515] = o_575_;
  assign o[516] = o_575_;
  assign o[517] = o_575_;
  assign o[518] = o_575_;
  assign o[519] = o_575_;
  assign o[520] = o_575_;
  assign o[521] = o_575_;
  assign o[522] = o_575_;
  assign o[523] = o_575_;
  assign o[524] = o_575_;
  assign o[525] = o_575_;
  assign o[526] = o_575_;
  assign o[527] = o_575_;
  assign o[528] = o_575_;
  assign o[529] = o_575_;
  assign o[530] = o_575_;
  assign o[531] = o_575_;
  assign o[532] = o_575_;
  assign o[533] = o_575_;
  assign o[534] = o_575_;
  assign o[535] = o_575_;
  assign o[536] = o_575_;
  assign o[537] = o_575_;
  assign o[538] = o_575_;
  assign o[539] = o_575_;
  assign o[540] = o_575_;
  assign o[541] = o_575_;
  assign o[542] = o_575_;
  assign o[543] = o_575_;
  assign o[544] = o_575_;
  assign o[545] = o_575_;
  assign o[546] = o_575_;
  assign o[547] = o_575_;
  assign o[548] = o_575_;
  assign o[549] = o_575_;
  assign o[550] = o_575_;
  assign o[551] = o_575_;
  assign o[552] = o_575_;
  assign o[553] = o_575_;
  assign o[554] = o_575_;
  assign o[555] = o_575_;
  assign o[556] = o_575_;
  assign o[557] = o_575_;
  assign o[558] = o_575_;
  assign o[559] = o_575_;
  assign o[560] = o_575_;
  assign o[561] = o_575_;
  assign o[562] = o_575_;
  assign o[563] = o_575_;
  assign o[564] = o_575_;
  assign o[565] = o_575_;
  assign o[566] = o_575_;
  assign o[567] = o_575_;
  assign o[568] = o_575_;
  assign o[569] = o_575_;
  assign o[570] = o_575_;
  assign o[571] = o_575_;
  assign o[572] = o_575_;
  assign o[573] = o_575_;
  assign o[574] = o_575_;
  assign o[575] = o_575_;
  assign o_511_ = i[7];
  assign o[448] = o_511_;
  assign o[449] = o_511_;
  assign o[450] = o_511_;
  assign o[451] = o_511_;
  assign o[452] = o_511_;
  assign o[453] = o_511_;
  assign o[454] = o_511_;
  assign o[455] = o_511_;
  assign o[456] = o_511_;
  assign o[457] = o_511_;
  assign o[458] = o_511_;
  assign o[459] = o_511_;
  assign o[460] = o_511_;
  assign o[461] = o_511_;
  assign o[462] = o_511_;
  assign o[463] = o_511_;
  assign o[464] = o_511_;
  assign o[465] = o_511_;
  assign o[466] = o_511_;
  assign o[467] = o_511_;
  assign o[468] = o_511_;
  assign o[469] = o_511_;
  assign o[470] = o_511_;
  assign o[471] = o_511_;
  assign o[472] = o_511_;
  assign o[473] = o_511_;
  assign o[474] = o_511_;
  assign o[475] = o_511_;
  assign o[476] = o_511_;
  assign o[477] = o_511_;
  assign o[478] = o_511_;
  assign o[479] = o_511_;
  assign o[480] = o_511_;
  assign o[481] = o_511_;
  assign o[482] = o_511_;
  assign o[483] = o_511_;
  assign o[484] = o_511_;
  assign o[485] = o_511_;
  assign o[486] = o_511_;
  assign o[487] = o_511_;
  assign o[488] = o_511_;
  assign o[489] = o_511_;
  assign o[490] = o_511_;
  assign o[491] = o_511_;
  assign o[492] = o_511_;
  assign o[493] = o_511_;
  assign o[494] = o_511_;
  assign o[495] = o_511_;
  assign o[496] = o_511_;
  assign o[497] = o_511_;
  assign o[498] = o_511_;
  assign o[499] = o_511_;
  assign o[500] = o_511_;
  assign o[501] = o_511_;
  assign o[502] = o_511_;
  assign o[503] = o_511_;
  assign o[504] = o_511_;
  assign o[505] = o_511_;
  assign o[506] = o_511_;
  assign o[507] = o_511_;
  assign o[508] = o_511_;
  assign o[509] = o_511_;
  assign o[510] = o_511_;
  assign o[511] = o_511_;
  assign o_447_ = i[6];
  assign o[384] = o_447_;
  assign o[385] = o_447_;
  assign o[386] = o_447_;
  assign o[387] = o_447_;
  assign o[388] = o_447_;
  assign o[389] = o_447_;
  assign o[390] = o_447_;
  assign o[391] = o_447_;
  assign o[392] = o_447_;
  assign o[393] = o_447_;
  assign o[394] = o_447_;
  assign o[395] = o_447_;
  assign o[396] = o_447_;
  assign o[397] = o_447_;
  assign o[398] = o_447_;
  assign o[399] = o_447_;
  assign o[400] = o_447_;
  assign o[401] = o_447_;
  assign o[402] = o_447_;
  assign o[403] = o_447_;
  assign o[404] = o_447_;
  assign o[405] = o_447_;
  assign o[406] = o_447_;
  assign o[407] = o_447_;
  assign o[408] = o_447_;
  assign o[409] = o_447_;
  assign o[410] = o_447_;
  assign o[411] = o_447_;
  assign o[412] = o_447_;
  assign o[413] = o_447_;
  assign o[414] = o_447_;
  assign o[415] = o_447_;
  assign o[416] = o_447_;
  assign o[417] = o_447_;
  assign o[418] = o_447_;
  assign o[419] = o_447_;
  assign o[420] = o_447_;
  assign o[421] = o_447_;
  assign o[422] = o_447_;
  assign o[423] = o_447_;
  assign o[424] = o_447_;
  assign o[425] = o_447_;
  assign o[426] = o_447_;
  assign o[427] = o_447_;
  assign o[428] = o_447_;
  assign o[429] = o_447_;
  assign o[430] = o_447_;
  assign o[431] = o_447_;
  assign o[432] = o_447_;
  assign o[433] = o_447_;
  assign o[434] = o_447_;
  assign o[435] = o_447_;
  assign o[436] = o_447_;
  assign o[437] = o_447_;
  assign o[438] = o_447_;
  assign o[439] = o_447_;
  assign o[440] = o_447_;
  assign o[441] = o_447_;
  assign o[442] = o_447_;
  assign o[443] = o_447_;
  assign o[444] = o_447_;
  assign o[445] = o_447_;
  assign o[446] = o_447_;
  assign o[447] = o_447_;
  assign o_383_ = i[5];
  assign o[320] = o_383_;
  assign o[321] = o_383_;
  assign o[322] = o_383_;
  assign o[323] = o_383_;
  assign o[324] = o_383_;
  assign o[325] = o_383_;
  assign o[326] = o_383_;
  assign o[327] = o_383_;
  assign o[328] = o_383_;
  assign o[329] = o_383_;
  assign o[330] = o_383_;
  assign o[331] = o_383_;
  assign o[332] = o_383_;
  assign o[333] = o_383_;
  assign o[334] = o_383_;
  assign o[335] = o_383_;
  assign o[336] = o_383_;
  assign o[337] = o_383_;
  assign o[338] = o_383_;
  assign o[339] = o_383_;
  assign o[340] = o_383_;
  assign o[341] = o_383_;
  assign o[342] = o_383_;
  assign o[343] = o_383_;
  assign o[344] = o_383_;
  assign o[345] = o_383_;
  assign o[346] = o_383_;
  assign o[347] = o_383_;
  assign o[348] = o_383_;
  assign o[349] = o_383_;
  assign o[350] = o_383_;
  assign o[351] = o_383_;
  assign o[352] = o_383_;
  assign o[353] = o_383_;
  assign o[354] = o_383_;
  assign o[355] = o_383_;
  assign o[356] = o_383_;
  assign o[357] = o_383_;
  assign o[358] = o_383_;
  assign o[359] = o_383_;
  assign o[360] = o_383_;
  assign o[361] = o_383_;
  assign o[362] = o_383_;
  assign o[363] = o_383_;
  assign o[364] = o_383_;
  assign o[365] = o_383_;
  assign o[366] = o_383_;
  assign o[367] = o_383_;
  assign o[368] = o_383_;
  assign o[369] = o_383_;
  assign o[370] = o_383_;
  assign o[371] = o_383_;
  assign o[372] = o_383_;
  assign o[373] = o_383_;
  assign o[374] = o_383_;
  assign o[375] = o_383_;
  assign o[376] = o_383_;
  assign o[377] = o_383_;
  assign o[378] = o_383_;
  assign o[379] = o_383_;
  assign o[380] = o_383_;
  assign o[381] = o_383_;
  assign o[382] = o_383_;
  assign o[383] = o_383_;
  assign o_319_ = i[4];
  assign o[256] = o_319_;
  assign o[257] = o_319_;
  assign o[258] = o_319_;
  assign o[259] = o_319_;
  assign o[260] = o_319_;
  assign o[261] = o_319_;
  assign o[262] = o_319_;
  assign o[263] = o_319_;
  assign o[264] = o_319_;
  assign o[265] = o_319_;
  assign o[266] = o_319_;
  assign o[267] = o_319_;
  assign o[268] = o_319_;
  assign o[269] = o_319_;
  assign o[270] = o_319_;
  assign o[271] = o_319_;
  assign o[272] = o_319_;
  assign o[273] = o_319_;
  assign o[274] = o_319_;
  assign o[275] = o_319_;
  assign o[276] = o_319_;
  assign o[277] = o_319_;
  assign o[278] = o_319_;
  assign o[279] = o_319_;
  assign o[280] = o_319_;
  assign o[281] = o_319_;
  assign o[282] = o_319_;
  assign o[283] = o_319_;
  assign o[284] = o_319_;
  assign o[285] = o_319_;
  assign o[286] = o_319_;
  assign o[287] = o_319_;
  assign o[288] = o_319_;
  assign o[289] = o_319_;
  assign o[290] = o_319_;
  assign o[291] = o_319_;
  assign o[292] = o_319_;
  assign o[293] = o_319_;
  assign o[294] = o_319_;
  assign o[295] = o_319_;
  assign o[296] = o_319_;
  assign o[297] = o_319_;
  assign o[298] = o_319_;
  assign o[299] = o_319_;
  assign o[300] = o_319_;
  assign o[301] = o_319_;
  assign o[302] = o_319_;
  assign o[303] = o_319_;
  assign o[304] = o_319_;
  assign o[305] = o_319_;
  assign o[306] = o_319_;
  assign o[307] = o_319_;
  assign o[308] = o_319_;
  assign o[309] = o_319_;
  assign o[310] = o_319_;
  assign o[311] = o_319_;
  assign o[312] = o_319_;
  assign o[313] = o_319_;
  assign o[314] = o_319_;
  assign o[315] = o_319_;
  assign o[316] = o_319_;
  assign o[317] = o_319_;
  assign o[318] = o_319_;
  assign o[319] = o_319_;
  assign o_255_ = i[3];
  assign o[192] = o_255_;
  assign o[193] = o_255_;
  assign o[194] = o_255_;
  assign o[195] = o_255_;
  assign o[196] = o_255_;
  assign o[197] = o_255_;
  assign o[198] = o_255_;
  assign o[199] = o_255_;
  assign o[200] = o_255_;
  assign o[201] = o_255_;
  assign o[202] = o_255_;
  assign o[203] = o_255_;
  assign o[204] = o_255_;
  assign o[205] = o_255_;
  assign o[206] = o_255_;
  assign o[207] = o_255_;
  assign o[208] = o_255_;
  assign o[209] = o_255_;
  assign o[210] = o_255_;
  assign o[211] = o_255_;
  assign o[212] = o_255_;
  assign o[213] = o_255_;
  assign o[214] = o_255_;
  assign o[215] = o_255_;
  assign o[216] = o_255_;
  assign o[217] = o_255_;
  assign o[218] = o_255_;
  assign o[219] = o_255_;
  assign o[220] = o_255_;
  assign o[221] = o_255_;
  assign o[222] = o_255_;
  assign o[223] = o_255_;
  assign o[224] = o_255_;
  assign o[225] = o_255_;
  assign o[226] = o_255_;
  assign o[227] = o_255_;
  assign o[228] = o_255_;
  assign o[229] = o_255_;
  assign o[230] = o_255_;
  assign o[231] = o_255_;
  assign o[232] = o_255_;
  assign o[233] = o_255_;
  assign o[234] = o_255_;
  assign o[235] = o_255_;
  assign o[236] = o_255_;
  assign o[237] = o_255_;
  assign o[238] = o_255_;
  assign o[239] = o_255_;
  assign o[240] = o_255_;
  assign o[241] = o_255_;
  assign o[242] = o_255_;
  assign o[243] = o_255_;
  assign o[244] = o_255_;
  assign o[245] = o_255_;
  assign o[246] = o_255_;
  assign o[247] = o_255_;
  assign o[248] = o_255_;
  assign o[249] = o_255_;
  assign o[250] = o_255_;
  assign o[251] = o_255_;
  assign o[252] = o_255_;
  assign o[253] = o_255_;
  assign o[254] = o_255_;
  assign o[255] = o_255_;
  assign o_191_ = i[2];
  assign o[128] = o_191_;
  assign o[129] = o_191_;
  assign o[130] = o_191_;
  assign o[131] = o_191_;
  assign o[132] = o_191_;
  assign o[133] = o_191_;
  assign o[134] = o_191_;
  assign o[135] = o_191_;
  assign o[136] = o_191_;
  assign o[137] = o_191_;
  assign o[138] = o_191_;
  assign o[139] = o_191_;
  assign o[140] = o_191_;
  assign o[141] = o_191_;
  assign o[142] = o_191_;
  assign o[143] = o_191_;
  assign o[144] = o_191_;
  assign o[145] = o_191_;
  assign o[146] = o_191_;
  assign o[147] = o_191_;
  assign o[148] = o_191_;
  assign o[149] = o_191_;
  assign o[150] = o_191_;
  assign o[151] = o_191_;
  assign o[152] = o_191_;
  assign o[153] = o_191_;
  assign o[154] = o_191_;
  assign o[155] = o_191_;
  assign o[156] = o_191_;
  assign o[157] = o_191_;
  assign o[158] = o_191_;
  assign o[159] = o_191_;
  assign o[160] = o_191_;
  assign o[161] = o_191_;
  assign o[162] = o_191_;
  assign o[163] = o_191_;
  assign o[164] = o_191_;
  assign o[165] = o_191_;
  assign o[166] = o_191_;
  assign o[167] = o_191_;
  assign o[168] = o_191_;
  assign o[169] = o_191_;
  assign o[170] = o_191_;
  assign o[171] = o_191_;
  assign o[172] = o_191_;
  assign o[173] = o_191_;
  assign o[174] = o_191_;
  assign o[175] = o_191_;
  assign o[176] = o_191_;
  assign o[177] = o_191_;
  assign o[178] = o_191_;
  assign o[179] = o_191_;
  assign o[180] = o_191_;
  assign o[181] = o_191_;
  assign o[182] = o_191_;
  assign o[183] = o_191_;
  assign o[184] = o_191_;
  assign o[185] = o_191_;
  assign o[186] = o_191_;
  assign o[187] = o_191_;
  assign o[188] = o_191_;
  assign o[189] = o_191_;
  assign o[190] = o_191_;
  assign o[191] = o_191_;
  assign o_127_ = i[1];
  assign o[64] = o_127_;
  assign o[65] = o_127_;
  assign o[66] = o_127_;
  assign o[67] = o_127_;
  assign o[68] = o_127_;
  assign o[69] = o_127_;
  assign o[70] = o_127_;
  assign o[71] = o_127_;
  assign o[72] = o_127_;
  assign o[73] = o_127_;
  assign o[74] = o_127_;
  assign o[75] = o_127_;
  assign o[76] = o_127_;
  assign o[77] = o_127_;
  assign o[78] = o_127_;
  assign o[79] = o_127_;
  assign o[80] = o_127_;
  assign o[81] = o_127_;
  assign o[82] = o_127_;
  assign o[83] = o_127_;
  assign o[84] = o_127_;
  assign o[85] = o_127_;
  assign o[86] = o_127_;
  assign o[87] = o_127_;
  assign o[88] = o_127_;
  assign o[89] = o_127_;
  assign o[90] = o_127_;
  assign o[91] = o_127_;
  assign o[92] = o_127_;
  assign o[93] = o_127_;
  assign o[94] = o_127_;
  assign o[95] = o_127_;
  assign o[96] = o_127_;
  assign o[97] = o_127_;
  assign o[98] = o_127_;
  assign o[99] = o_127_;
  assign o[100] = o_127_;
  assign o[101] = o_127_;
  assign o[102] = o_127_;
  assign o[103] = o_127_;
  assign o[104] = o_127_;
  assign o[105] = o_127_;
  assign o[106] = o_127_;
  assign o[107] = o_127_;
  assign o[108] = o_127_;
  assign o[109] = o_127_;
  assign o[110] = o_127_;
  assign o[111] = o_127_;
  assign o[112] = o_127_;
  assign o[113] = o_127_;
  assign o[114] = o_127_;
  assign o[115] = o_127_;
  assign o[116] = o_127_;
  assign o[117] = o_127_;
  assign o[118] = o_127_;
  assign o[119] = o_127_;
  assign o[120] = o_127_;
  assign o[121] = o_127_;
  assign o[122] = o_127_;
  assign o[123] = o_127_;
  assign o[124] = o_127_;
  assign o[125] = o_127_;
  assign o[126] = o_127_;
  assign o[127] = o_127_;
  assign o_63_ = i[0];
  assign o[0] = o_63_;
  assign o[1] = o_63_;
  assign o[2] = o_63_;
  assign o[3] = o_63_;
  assign o[4] = o_63_;
  assign o[5] = o_63_;
  assign o[6] = o_63_;
  assign o[7] = o_63_;
  assign o[8] = o_63_;
  assign o[9] = o_63_;
  assign o[10] = o_63_;
  assign o[11] = o_63_;
  assign o[12] = o_63_;
  assign o[13] = o_63_;
  assign o[14] = o_63_;
  assign o[15] = o_63_;
  assign o[16] = o_63_;
  assign o[17] = o_63_;
  assign o[18] = o_63_;
  assign o[19] = o_63_;
  assign o[20] = o_63_;
  assign o[21] = o_63_;
  assign o[22] = o_63_;
  assign o[23] = o_63_;
  assign o[24] = o_63_;
  assign o[25] = o_63_;
  assign o[26] = o_63_;
  assign o[27] = o_63_;
  assign o[28] = o_63_;
  assign o[29] = o_63_;
  assign o[30] = o_63_;
  assign o[31] = o_63_;
  assign o[32] = o_63_;
  assign o[33] = o_63_;
  assign o[34] = o_63_;
  assign o[35] = o_63_;
  assign o[36] = o_63_;
  assign o[37] = o_63_;
  assign o[38] = o_63_;
  assign o[39] = o_63_;
  assign o[40] = o_63_;
  assign o[41] = o_63_;
  assign o[42] = o_63_;
  assign o[43] = o_63_;
  assign o[44] = o_63_;
  assign o[45] = o_63_;
  assign o[46] = o_63_;
  assign o[47] = o_63_;
  assign o[48] = o_63_;
  assign o[49] = o_63_;
  assign o[50] = o_63_;
  assign o[51] = o_63_;
  assign o[52] = o_63_;
  assign o[53] = o_63_;
  assign o[54] = o_63_;
  assign o[55] = o_63_;
  assign o[56] = o_63_;
  assign o[57] = o_63_;
  assign o[58] = o_63_;
  assign o[59] = o_63_;
  assign o[60] = o_63_;
  assign o[61] = o_63_;
  assign o[62] = o_63_;
  assign o[63] = o_63_;

endmodule

