

module top
(
  clk_i,
  reset_i,
  valid_i,
  data_i,
  ready_and_o,
  valid_o,
  data_o,
  yumi_i
);

  input [2047:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input valid_i;
  input yumi_i;
  output ready_and_o;
  output valid_o;

  bsg_parallel_in_serial_out
  wrapper
  (
    .data_i(data_i),
    .data_o(data_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .valid_i(valid_i),
    .yumi_i(yumi_i),
    .ready_and_o(ready_and_o),
    .valid_o(valid_o)
  );


endmodule



module bsg_array_reverse_width_p32_els_p64
(
  i,
  o
);

  input [2047:0] i;
  output [2047:0] o;
  wire [2047:0] o;
  assign o[2047] = i[31];
  assign o[2046] = i[30];
  assign o[2045] = i[29];
  assign o[2044] = i[28];
  assign o[2043] = i[27];
  assign o[2042] = i[26];
  assign o[2041] = i[25];
  assign o[2040] = i[24];
  assign o[2039] = i[23];
  assign o[2038] = i[22];
  assign o[2037] = i[21];
  assign o[2036] = i[20];
  assign o[2035] = i[19];
  assign o[2034] = i[18];
  assign o[2033] = i[17];
  assign o[2032] = i[16];
  assign o[2031] = i[15];
  assign o[2030] = i[14];
  assign o[2029] = i[13];
  assign o[2028] = i[12];
  assign o[2027] = i[11];
  assign o[2026] = i[10];
  assign o[2025] = i[9];
  assign o[2024] = i[8];
  assign o[2023] = i[7];
  assign o[2022] = i[6];
  assign o[2021] = i[5];
  assign o[2020] = i[4];
  assign o[2019] = i[3];
  assign o[2018] = i[2];
  assign o[2017] = i[1];
  assign o[2016] = i[0];
  assign o[2015] = i[63];
  assign o[2014] = i[62];
  assign o[2013] = i[61];
  assign o[2012] = i[60];
  assign o[2011] = i[59];
  assign o[2010] = i[58];
  assign o[2009] = i[57];
  assign o[2008] = i[56];
  assign o[2007] = i[55];
  assign o[2006] = i[54];
  assign o[2005] = i[53];
  assign o[2004] = i[52];
  assign o[2003] = i[51];
  assign o[2002] = i[50];
  assign o[2001] = i[49];
  assign o[2000] = i[48];
  assign o[1999] = i[47];
  assign o[1998] = i[46];
  assign o[1997] = i[45];
  assign o[1996] = i[44];
  assign o[1995] = i[43];
  assign o[1994] = i[42];
  assign o[1993] = i[41];
  assign o[1992] = i[40];
  assign o[1991] = i[39];
  assign o[1990] = i[38];
  assign o[1989] = i[37];
  assign o[1988] = i[36];
  assign o[1987] = i[35];
  assign o[1986] = i[34];
  assign o[1985] = i[33];
  assign o[1984] = i[32];
  assign o[1983] = i[95];
  assign o[1982] = i[94];
  assign o[1981] = i[93];
  assign o[1980] = i[92];
  assign o[1979] = i[91];
  assign o[1978] = i[90];
  assign o[1977] = i[89];
  assign o[1976] = i[88];
  assign o[1975] = i[87];
  assign o[1974] = i[86];
  assign o[1973] = i[85];
  assign o[1972] = i[84];
  assign o[1971] = i[83];
  assign o[1970] = i[82];
  assign o[1969] = i[81];
  assign o[1968] = i[80];
  assign o[1967] = i[79];
  assign o[1966] = i[78];
  assign o[1965] = i[77];
  assign o[1964] = i[76];
  assign o[1963] = i[75];
  assign o[1962] = i[74];
  assign o[1961] = i[73];
  assign o[1960] = i[72];
  assign o[1959] = i[71];
  assign o[1958] = i[70];
  assign o[1957] = i[69];
  assign o[1956] = i[68];
  assign o[1955] = i[67];
  assign o[1954] = i[66];
  assign o[1953] = i[65];
  assign o[1952] = i[64];
  assign o[1951] = i[127];
  assign o[1950] = i[126];
  assign o[1949] = i[125];
  assign o[1948] = i[124];
  assign o[1947] = i[123];
  assign o[1946] = i[122];
  assign o[1945] = i[121];
  assign o[1944] = i[120];
  assign o[1943] = i[119];
  assign o[1942] = i[118];
  assign o[1941] = i[117];
  assign o[1940] = i[116];
  assign o[1939] = i[115];
  assign o[1938] = i[114];
  assign o[1937] = i[113];
  assign o[1936] = i[112];
  assign o[1935] = i[111];
  assign o[1934] = i[110];
  assign o[1933] = i[109];
  assign o[1932] = i[108];
  assign o[1931] = i[107];
  assign o[1930] = i[106];
  assign o[1929] = i[105];
  assign o[1928] = i[104];
  assign o[1927] = i[103];
  assign o[1926] = i[102];
  assign o[1925] = i[101];
  assign o[1924] = i[100];
  assign o[1923] = i[99];
  assign o[1922] = i[98];
  assign o[1921] = i[97];
  assign o[1920] = i[96];
  assign o[1919] = i[159];
  assign o[1918] = i[158];
  assign o[1917] = i[157];
  assign o[1916] = i[156];
  assign o[1915] = i[155];
  assign o[1914] = i[154];
  assign o[1913] = i[153];
  assign o[1912] = i[152];
  assign o[1911] = i[151];
  assign o[1910] = i[150];
  assign o[1909] = i[149];
  assign o[1908] = i[148];
  assign o[1907] = i[147];
  assign o[1906] = i[146];
  assign o[1905] = i[145];
  assign o[1904] = i[144];
  assign o[1903] = i[143];
  assign o[1902] = i[142];
  assign o[1901] = i[141];
  assign o[1900] = i[140];
  assign o[1899] = i[139];
  assign o[1898] = i[138];
  assign o[1897] = i[137];
  assign o[1896] = i[136];
  assign o[1895] = i[135];
  assign o[1894] = i[134];
  assign o[1893] = i[133];
  assign o[1892] = i[132];
  assign o[1891] = i[131];
  assign o[1890] = i[130];
  assign o[1889] = i[129];
  assign o[1888] = i[128];
  assign o[1887] = i[191];
  assign o[1886] = i[190];
  assign o[1885] = i[189];
  assign o[1884] = i[188];
  assign o[1883] = i[187];
  assign o[1882] = i[186];
  assign o[1881] = i[185];
  assign o[1880] = i[184];
  assign o[1879] = i[183];
  assign o[1878] = i[182];
  assign o[1877] = i[181];
  assign o[1876] = i[180];
  assign o[1875] = i[179];
  assign o[1874] = i[178];
  assign o[1873] = i[177];
  assign o[1872] = i[176];
  assign o[1871] = i[175];
  assign o[1870] = i[174];
  assign o[1869] = i[173];
  assign o[1868] = i[172];
  assign o[1867] = i[171];
  assign o[1866] = i[170];
  assign o[1865] = i[169];
  assign o[1864] = i[168];
  assign o[1863] = i[167];
  assign o[1862] = i[166];
  assign o[1861] = i[165];
  assign o[1860] = i[164];
  assign o[1859] = i[163];
  assign o[1858] = i[162];
  assign o[1857] = i[161];
  assign o[1856] = i[160];
  assign o[1855] = i[223];
  assign o[1854] = i[222];
  assign o[1853] = i[221];
  assign o[1852] = i[220];
  assign o[1851] = i[219];
  assign o[1850] = i[218];
  assign o[1849] = i[217];
  assign o[1848] = i[216];
  assign o[1847] = i[215];
  assign o[1846] = i[214];
  assign o[1845] = i[213];
  assign o[1844] = i[212];
  assign o[1843] = i[211];
  assign o[1842] = i[210];
  assign o[1841] = i[209];
  assign o[1840] = i[208];
  assign o[1839] = i[207];
  assign o[1838] = i[206];
  assign o[1837] = i[205];
  assign o[1836] = i[204];
  assign o[1835] = i[203];
  assign o[1834] = i[202];
  assign o[1833] = i[201];
  assign o[1832] = i[200];
  assign o[1831] = i[199];
  assign o[1830] = i[198];
  assign o[1829] = i[197];
  assign o[1828] = i[196];
  assign o[1827] = i[195];
  assign o[1826] = i[194];
  assign o[1825] = i[193];
  assign o[1824] = i[192];
  assign o[1823] = i[255];
  assign o[1822] = i[254];
  assign o[1821] = i[253];
  assign o[1820] = i[252];
  assign o[1819] = i[251];
  assign o[1818] = i[250];
  assign o[1817] = i[249];
  assign o[1816] = i[248];
  assign o[1815] = i[247];
  assign o[1814] = i[246];
  assign o[1813] = i[245];
  assign o[1812] = i[244];
  assign o[1811] = i[243];
  assign o[1810] = i[242];
  assign o[1809] = i[241];
  assign o[1808] = i[240];
  assign o[1807] = i[239];
  assign o[1806] = i[238];
  assign o[1805] = i[237];
  assign o[1804] = i[236];
  assign o[1803] = i[235];
  assign o[1802] = i[234];
  assign o[1801] = i[233];
  assign o[1800] = i[232];
  assign o[1799] = i[231];
  assign o[1798] = i[230];
  assign o[1797] = i[229];
  assign o[1796] = i[228];
  assign o[1795] = i[227];
  assign o[1794] = i[226];
  assign o[1793] = i[225];
  assign o[1792] = i[224];
  assign o[1791] = i[287];
  assign o[1790] = i[286];
  assign o[1789] = i[285];
  assign o[1788] = i[284];
  assign o[1787] = i[283];
  assign o[1786] = i[282];
  assign o[1785] = i[281];
  assign o[1784] = i[280];
  assign o[1783] = i[279];
  assign o[1782] = i[278];
  assign o[1781] = i[277];
  assign o[1780] = i[276];
  assign o[1779] = i[275];
  assign o[1778] = i[274];
  assign o[1777] = i[273];
  assign o[1776] = i[272];
  assign o[1775] = i[271];
  assign o[1774] = i[270];
  assign o[1773] = i[269];
  assign o[1772] = i[268];
  assign o[1771] = i[267];
  assign o[1770] = i[266];
  assign o[1769] = i[265];
  assign o[1768] = i[264];
  assign o[1767] = i[263];
  assign o[1766] = i[262];
  assign o[1765] = i[261];
  assign o[1764] = i[260];
  assign o[1763] = i[259];
  assign o[1762] = i[258];
  assign o[1761] = i[257];
  assign o[1760] = i[256];
  assign o[1759] = i[319];
  assign o[1758] = i[318];
  assign o[1757] = i[317];
  assign o[1756] = i[316];
  assign o[1755] = i[315];
  assign o[1754] = i[314];
  assign o[1753] = i[313];
  assign o[1752] = i[312];
  assign o[1751] = i[311];
  assign o[1750] = i[310];
  assign o[1749] = i[309];
  assign o[1748] = i[308];
  assign o[1747] = i[307];
  assign o[1746] = i[306];
  assign o[1745] = i[305];
  assign o[1744] = i[304];
  assign o[1743] = i[303];
  assign o[1742] = i[302];
  assign o[1741] = i[301];
  assign o[1740] = i[300];
  assign o[1739] = i[299];
  assign o[1738] = i[298];
  assign o[1737] = i[297];
  assign o[1736] = i[296];
  assign o[1735] = i[295];
  assign o[1734] = i[294];
  assign o[1733] = i[293];
  assign o[1732] = i[292];
  assign o[1731] = i[291];
  assign o[1730] = i[290];
  assign o[1729] = i[289];
  assign o[1728] = i[288];
  assign o[1727] = i[351];
  assign o[1726] = i[350];
  assign o[1725] = i[349];
  assign o[1724] = i[348];
  assign o[1723] = i[347];
  assign o[1722] = i[346];
  assign o[1721] = i[345];
  assign o[1720] = i[344];
  assign o[1719] = i[343];
  assign o[1718] = i[342];
  assign o[1717] = i[341];
  assign o[1716] = i[340];
  assign o[1715] = i[339];
  assign o[1714] = i[338];
  assign o[1713] = i[337];
  assign o[1712] = i[336];
  assign o[1711] = i[335];
  assign o[1710] = i[334];
  assign o[1709] = i[333];
  assign o[1708] = i[332];
  assign o[1707] = i[331];
  assign o[1706] = i[330];
  assign o[1705] = i[329];
  assign o[1704] = i[328];
  assign o[1703] = i[327];
  assign o[1702] = i[326];
  assign o[1701] = i[325];
  assign o[1700] = i[324];
  assign o[1699] = i[323];
  assign o[1698] = i[322];
  assign o[1697] = i[321];
  assign o[1696] = i[320];
  assign o[1695] = i[383];
  assign o[1694] = i[382];
  assign o[1693] = i[381];
  assign o[1692] = i[380];
  assign o[1691] = i[379];
  assign o[1690] = i[378];
  assign o[1689] = i[377];
  assign o[1688] = i[376];
  assign o[1687] = i[375];
  assign o[1686] = i[374];
  assign o[1685] = i[373];
  assign o[1684] = i[372];
  assign o[1683] = i[371];
  assign o[1682] = i[370];
  assign o[1681] = i[369];
  assign o[1680] = i[368];
  assign o[1679] = i[367];
  assign o[1678] = i[366];
  assign o[1677] = i[365];
  assign o[1676] = i[364];
  assign o[1675] = i[363];
  assign o[1674] = i[362];
  assign o[1673] = i[361];
  assign o[1672] = i[360];
  assign o[1671] = i[359];
  assign o[1670] = i[358];
  assign o[1669] = i[357];
  assign o[1668] = i[356];
  assign o[1667] = i[355];
  assign o[1666] = i[354];
  assign o[1665] = i[353];
  assign o[1664] = i[352];
  assign o[1663] = i[415];
  assign o[1662] = i[414];
  assign o[1661] = i[413];
  assign o[1660] = i[412];
  assign o[1659] = i[411];
  assign o[1658] = i[410];
  assign o[1657] = i[409];
  assign o[1656] = i[408];
  assign o[1655] = i[407];
  assign o[1654] = i[406];
  assign o[1653] = i[405];
  assign o[1652] = i[404];
  assign o[1651] = i[403];
  assign o[1650] = i[402];
  assign o[1649] = i[401];
  assign o[1648] = i[400];
  assign o[1647] = i[399];
  assign o[1646] = i[398];
  assign o[1645] = i[397];
  assign o[1644] = i[396];
  assign o[1643] = i[395];
  assign o[1642] = i[394];
  assign o[1641] = i[393];
  assign o[1640] = i[392];
  assign o[1639] = i[391];
  assign o[1638] = i[390];
  assign o[1637] = i[389];
  assign o[1636] = i[388];
  assign o[1635] = i[387];
  assign o[1634] = i[386];
  assign o[1633] = i[385];
  assign o[1632] = i[384];
  assign o[1631] = i[447];
  assign o[1630] = i[446];
  assign o[1629] = i[445];
  assign o[1628] = i[444];
  assign o[1627] = i[443];
  assign o[1626] = i[442];
  assign o[1625] = i[441];
  assign o[1624] = i[440];
  assign o[1623] = i[439];
  assign o[1622] = i[438];
  assign o[1621] = i[437];
  assign o[1620] = i[436];
  assign o[1619] = i[435];
  assign o[1618] = i[434];
  assign o[1617] = i[433];
  assign o[1616] = i[432];
  assign o[1615] = i[431];
  assign o[1614] = i[430];
  assign o[1613] = i[429];
  assign o[1612] = i[428];
  assign o[1611] = i[427];
  assign o[1610] = i[426];
  assign o[1609] = i[425];
  assign o[1608] = i[424];
  assign o[1607] = i[423];
  assign o[1606] = i[422];
  assign o[1605] = i[421];
  assign o[1604] = i[420];
  assign o[1603] = i[419];
  assign o[1602] = i[418];
  assign o[1601] = i[417];
  assign o[1600] = i[416];
  assign o[1599] = i[479];
  assign o[1598] = i[478];
  assign o[1597] = i[477];
  assign o[1596] = i[476];
  assign o[1595] = i[475];
  assign o[1594] = i[474];
  assign o[1593] = i[473];
  assign o[1592] = i[472];
  assign o[1591] = i[471];
  assign o[1590] = i[470];
  assign o[1589] = i[469];
  assign o[1588] = i[468];
  assign o[1587] = i[467];
  assign o[1586] = i[466];
  assign o[1585] = i[465];
  assign o[1584] = i[464];
  assign o[1583] = i[463];
  assign o[1582] = i[462];
  assign o[1581] = i[461];
  assign o[1580] = i[460];
  assign o[1579] = i[459];
  assign o[1578] = i[458];
  assign o[1577] = i[457];
  assign o[1576] = i[456];
  assign o[1575] = i[455];
  assign o[1574] = i[454];
  assign o[1573] = i[453];
  assign o[1572] = i[452];
  assign o[1571] = i[451];
  assign o[1570] = i[450];
  assign o[1569] = i[449];
  assign o[1568] = i[448];
  assign o[1567] = i[511];
  assign o[1566] = i[510];
  assign o[1565] = i[509];
  assign o[1564] = i[508];
  assign o[1563] = i[507];
  assign o[1562] = i[506];
  assign o[1561] = i[505];
  assign o[1560] = i[504];
  assign o[1559] = i[503];
  assign o[1558] = i[502];
  assign o[1557] = i[501];
  assign o[1556] = i[500];
  assign o[1555] = i[499];
  assign o[1554] = i[498];
  assign o[1553] = i[497];
  assign o[1552] = i[496];
  assign o[1551] = i[495];
  assign o[1550] = i[494];
  assign o[1549] = i[493];
  assign o[1548] = i[492];
  assign o[1547] = i[491];
  assign o[1546] = i[490];
  assign o[1545] = i[489];
  assign o[1544] = i[488];
  assign o[1543] = i[487];
  assign o[1542] = i[486];
  assign o[1541] = i[485];
  assign o[1540] = i[484];
  assign o[1539] = i[483];
  assign o[1538] = i[482];
  assign o[1537] = i[481];
  assign o[1536] = i[480];
  assign o[1535] = i[543];
  assign o[1534] = i[542];
  assign o[1533] = i[541];
  assign o[1532] = i[540];
  assign o[1531] = i[539];
  assign o[1530] = i[538];
  assign o[1529] = i[537];
  assign o[1528] = i[536];
  assign o[1527] = i[535];
  assign o[1526] = i[534];
  assign o[1525] = i[533];
  assign o[1524] = i[532];
  assign o[1523] = i[531];
  assign o[1522] = i[530];
  assign o[1521] = i[529];
  assign o[1520] = i[528];
  assign o[1519] = i[527];
  assign o[1518] = i[526];
  assign o[1517] = i[525];
  assign o[1516] = i[524];
  assign o[1515] = i[523];
  assign o[1514] = i[522];
  assign o[1513] = i[521];
  assign o[1512] = i[520];
  assign o[1511] = i[519];
  assign o[1510] = i[518];
  assign o[1509] = i[517];
  assign o[1508] = i[516];
  assign o[1507] = i[515];
  assign o[1506] = i[514];
  assign o[1505] = i[513];
  assign o[1504] = i[512];
  assign o[1503] = i[575];
  assign o[1502] = i[574];
  assign o[1501] = i[573];
  assign o[1500] = i[572];
  assign o[1499] = i[571];
  assign o[1498] = i[570];
  assign o[1497] = i[569];
  assign o[1496] = i[568];
  assign o[1495] = i[567];
  assign o[1494] = i[566];
  assign o[1493] = i[565];
  assign o[1492] = i[564];
  assign o[1491] = i[563];
  assign o[1490] = i[562];
  assign o[1489] = i[561];
  assign o[1488] = i[560];
  assign o[1487] = i[559];
  assign o[1486] = i[558];
  assign o[1485] = i[557];
  assign o[1484] = i[556];
  assign o[1483] = i[555];
  assign o[1482] = i[554];
  assign o[1481] = i[553];
  assign o[1480] = i[552];
  assign o[1479] = i[551];
  assign o[1478] = i[550];
  assign o[1477] = i[549];
  assign o[1476] = i[548];
  assign o[1475] = i[547];
  assign o[1474] = i[546];
  assign o[1473] = i[545];
  assign o[1472] = i[544];
  assign o[1471] = i[607];
  assign o[1470] = i[606];
  assign o[1469] = i[605];
  assign o[1468] = i[604];
  assign o[1467] = i[603];
  assign o[1466] = i[602];
  assign o[1465] = i[601];
  assign o[1464] = i[600];
  assign o[1463] = i[599];
  assign o[1462] = i[598];
  assign o[1461] = i[597];
  assign o[1460] = i[596];
  assign o[1459] = i[595];
  assign o[1458] = i[594];
  assign o[1457] = i[593];
  assign o[1456] = i[592];
  assign o[1455] = i[591];
  assign o[1454] = i[590];
  assign o[1453] = i[589];
  assign o[1452] = i[588];
  assign o[1451] = i[587];
  assign o[1450] = i[586];
  assign o[1449] = i[585];
  assign o[1448] = i[584];
  assign o[1447] = i[583];
  assign o[1446] = i[582];
  assign o[1445] = i[581];
  assign o[1444] = i[580];
  assign o[1443] = i[579];
  assign o[1442] = i[578];
  assign o[1441] = i[577];
  assign o[1440] = i[576];
  assign o[1439] = i[639];
  assign o[1438] = i[638];
  assign o[1437] = i[637];
  assign o[1436] = i[636];
  assign o[1435] = i[635];
  assign o[1434] = i[634];
  assign o[1433] = i[633];
  assign o[1432] = i[632];
  assign o[1431] = i[631];
  assign o[1430] = i[630];
  assign o[1429] = i[629];
  assign o[1428] = i[628];
  assign o[1427] = i[627];
  assign o[1426] = i[626];
  assign o[1425] = i[625];
  assign o[1424] = i[624];
  assign o[1423] = i[623];
  assign o[1422] = i[622];
  assign o[1421] = i[621];
  assign o[1420] = i[620];
  assign o[1419] = i[619];
  assign o[1418] = i[618];
  assign o[1417] = i[617];
  assign o[1416] = i[616];
  assign o[1415] = i[615];
  assign o[1414] = i[614];
  assign o[1413] = i[613];
  assign o[1412] = i[612];
  assign o[1411] = i[611];
  assign o[1410] = i[610];
  assign o[1409] = i[609];
  assign o[1408] = i[608];
  assign o[1407] = i[671];
  assign o[1406] = i[670];
  assign o[1405] = i[669];
  assign o[1404] = i[668];
  assign o[1403] = i[667];
  assign o[1402] = i[666];
  assign o[1401] = i[665];
  assign o[1400] = i[664];
  assign o[1399] = i[663];
  assign o[1398] = i[662];
  assign o[1397] = i[661];
  assign o[1396] = i[660];
  assign o[1395] = i[659];
  assign o[1394] = i[658];
  assign o[1393] = i[657];
  assign o[1392] = i[656];
  assign o[1391] = i[655];
  assign o[1390] = i[654];
  assign o[1389] = i[653];
  assign o[1388] = i[652];
  assign o[1387] = i[651];
  assign o[1386] = i[650];
  assign o[1385] = i[649];
  assign o[1384] = i[648];
  assign o[1383] = i[647];
  assign o[1382] = i[646];
  assign o[1381] = i[645];
  assign o[1380] = i[644];
  assign o[1379] = i[643];
  assign o[1378] = i[642];
  assign o[1377] = i[641];
  assign o[1376] = i[640];
  assign o[1375] = i[703];
  assign o[1374] = i[702];
  assign o[1373] = i[701];
  assign o[1372] = i[700];
  assign o[1371] = i[699];
  assign o[1370] = i[698];
  assign o[1369] = i[697];
  assign o[1368] = i[696];
  assign o[1367] = i[695];
  assign o[1366] = i[694];
  assign o[1365] = i[693];
  assign o[1364] = i[692];
  assign o[1363] = i[691];
  assign o[1362] = i[690];
  assign o[1361] = i[689];
  assign o[1360] = i[688];
  assign o[1359] = i[687];
  assign o[1358] = i[686];
  assign o[1357] = i[685];
  assign o[1356] = i[684];
  assign o[1355] = i[683];
  assign o[1354] = i[682];
  assign o[1353] = i[681];
  assign o[1352] = i[680];
  assign o[1351] = i[679];
  assign o[1350] = i[678];
  assign o[1349] = i[677];
  assign o[1348] = i[676];
  assign o[1347] = i[675];
  assign o[1346] = i[674];
  assign o[1345] = i[673];
  assign o[1344] = i[672];
  assign o[1343] = i[735];
  assign o[1342] = i[734];
  assign o[1341] = i[733];
  assign o[1340] = i[732];
  assign o[1339] = i[731];
  assign o[1338] = i[730];
  assign o[1337] = i[729];
  assign o[1336] = i[728];
  assign o[1335] = i[727];
  assign o[1334] = i[726];
  assign o[1333] = i[725];
  assign o[1332] = i[724];
  assign o[1331] = i[723];
  assign o[1330] = i[722];
  assign o[1329] = i[721];
  assign o[1328] = i[720];
  assign o[1327] = i[719];
  assign o[1326] = i[718];
  assign o[1325] = i[717];
  assign o[1324] = i[716];
  assign o[1323] = i[715];
  assign o[1322] = i[714];
  assign o[1321] = i[713];
  assign o[1320] = i[712];
  assign o[1319] = i[711];
  assign o[1318] = i[710];
  assign o[1317] = i[709];
  assign o[1316] = i[708];
  assign o[1315] = i[707];
  assign o[1314] = i[706];
  assign o[1313] = i[705];
  assign o[1312] = i[704];
  assign o[1311] = i[767];
  assign o[1310] = i[766];
  assign o[1309] = i[765];
  assign o[1308] = i[764];
  assign o[1307] = i[763];
  assign o[1306] = i[762];
  assign o[1305] = i[761];
  assign o[1304] = i[760];
  assign o[1303] = i[759];
  assign o[1302] = i[758];
  assign o[1301] = i[757];
  assign o[1300] = i[756];
  assign o[1299] = i[755];
  assign o[1298] = i[754];
  assign o[1297] = i[753];
  assign o[1296] = i[752];
  assign o[1295] = i[751];
  assign o[1294] = i[750];
  assign o[1293] = i[749];
  assign o[1292] = i[748];
  assign o[1291] = i[747];
  assign o[1290] = i[746];
  assign o[1289] = i[745];
  assign o[1288] = i[744];
  assign o[1287] = i[743];
  assign o[1286] = i[742];
  assign o[1285] = i[741];
  assign o[1284] = i[740];
  assign o[1283] = i[739];
  assign o[1282] = i[738];
  assign o[1281] = i[737];
  assign o[1280] = i[736];
  assign o[1279] = i[799];
  assign o[1278] = i[798];
  assign o[1277] = i[797];
  assign o[1276] = i[796];
  assign o[1275] = i[795];
  assign o[1274] = i[794];
  assign o[1273] = i[793];
  assign o[1272] = i[792];
  assign o[1271] = i[791];
  assign o[1270] = i[790];
  assign o[1269] = i[789];
  assign o[1268] = i[788];
  assign o[1267] = i[787];
  assign o[1266] = i[786];
  assign o[1265] = i[785];
  assign o[1264] = i[784];
  assign o[1263] = i[783];
  assign o[1262] = i[782];
  assign o[1261] = i[781];
  assign o[1260] = i[780];
  assign o[1259] = i[779];
  assign o[1258] = i[778];
  assign o[1257] = i[777];
  assign o[1256] = i[776];
  assign o[1255] = i[775];
  assign o[1254] = i[774];
  assign o[1253] = i[773];
  assign o[1252] = i[772];
  assign o[1251] = i[771];
  assign o[1250] = i[770];
  assign o[1249] = i[769];
  assign o[1248] = i[768];
  assign o[1247] = i[831];
  assign o[1246] = i[830];
  assign o[1245] = i[829];
  assign o[1244] = i[828];
  assign o[1243] = i[827];
  assign o[1242] = i[826];
  assign o[1241] = i[825];
  assign o[1240] = i[824];
  assign o[1239] = i[823];
  assign o[1238] = i[822];
  assign o[1237] = i[821];
  assign o[1236] = i[820];
  assign o[1235] = i[819];
  assign o[1234] = i[818];
  assign o[1233] = i[817];
  assign o[1232] = i[816];
  assign o[1231] = i[815];
  assign o[1230] = i[814];
  assign o[1229] = i[813];
  assign o[1228] = i[812];
  assign o[1227] = i[811];
  assign o[1226] = i[810];
  assign o[1225] = i[809];
  assign o[1224] = i[808];
  assign o[1223] = i[807];
  assign o[1222] = i[806];
  assign o[1221] = i[805];
  assign o[1220] = i[804];
  assign o[1219] = i[803];
  assign o[1218] = i[802];
  assign o[1217] = i[801];
  assign o[1216] = i[800];
  assign o[1215] = i[863];
  assign o[1214] = i[862];
  assign o[1213] = i[861];
  assign o[1212] = i[860];
  assign o[1211] = i[859];
  assign o[1210] = i[858];
  assign o[1209] = i[857];
  assign o[1208] = i[856];
  assign o[1207] = i[855];
  assign o[1206] = i[854];
  assign o[1205] = i[853];
  assign o[1204] = i[852];
  assign o[1203] = i[851];
  assign o[1202] = i[850];
  assign o[1201] = i[849];
  assign o[1200] = i[848];
  assign o[1199] = i[847];
  assign o[1198] = i[846];
  assign o[1197] = i[845];
  assign o[1196] = i[844];
  assign o[1195] = i[843];
  assign o[1194] = i[842];
  assign o[1193] = i[841];
  assign o[1192] = i[840];
  assign o[1191] = i[839];
  assign o[1190] = i[838];
  assign o[1189] = i[837];
  assign o[1188] = i[836];
  assign o[1187] = i[835];
  assign o[1186] = i[834];
  assign o[1185] = i[833];
  assign o[1184] = i[832];
  assign o[1183] = i[895];
  assign o[1182] = i[894];
  assign o[1181] = i[893];
  assign o[1180] = i[892];
  assign o[1179] = i[891];
  assign o[1178] = i[890];
  assign o[1177] = i[889];
  assign o[1176] = i[888];
  assign o[1175] = i[887];
  assign o[1174] = i[886];
  assign o[1173] = i[885];
  assign o[1172] = i[884];
  assign o[1171] = i[883];
  assign o[1170] = i[882];
  assign o[1169] = i[881];
  assign o[1168] = i[880];
  assign o[1167] = i[879];
  assign o[1166] = i[878];
  assign o[1165] = i[877];
  assign o[1164] = i[876];
  assign o[1163] = i[875];
  assign o[1162] = i[874];
  assign o[1161] = i[873];
  assign o[1160] = i[872];
  assign o[1159] = i[871];
  assign o[1158] = i[870];
  assign o[1157] = i[869];
  assign o[1156] = i[868];
  assign o[1155] = i[867];
  assign o[1154] = i[866];
  assign o[1153] = i[865];
  assign o[1152] = i[864];
  assign o[1151] = i[927];
  assign o[1150] = i[926];
  assign o[1149] = i[925];
  assign o[1148] = i[924];
  assign o[1147] = i[923];
  assign o[1146] = i[922];
  assign o[1145] = i[921];
  assign o[1144] = i[920];
  assign o[1143] = i[919];
  assign o[1142] = i[918];
  assign o[1141] = i[917];
  assign o[1140] = i[916];
  assign o[1139] = i[915];
  assign o[1138] = i[914];
  assign o[1137] = i[913];
  assign o[1136] = i[912];
  assign o[1135] = i[911];
  assign o[1134] = i[910];
  assign o[1133] = i[909];
  assign o[1132] = i[908];
  assign o[1131] = i[907];
  assign o[1130] = i[906];
  assign o[1129] = i[905];
  assign o[1128] = i[904];
  assign o[1127] = i[903];
  assign o[1126] = i[902];
  assign o[1125] = i[901];
  assign o[1124] = i[900];
  assign o[1123] = i[899];
  assign o[1122] = i[898];
  assign o[1121] = i[897];
  assign o[1120] = i[896];
  assign o[1119] = i[959];
  assign o[1118] = i[958];
  assign o[1117] = i[957];
  assign o[1116] = i[956];
  assign o[1115] = i[955];
  assign o[1114] = i[954];
  assign o[1113] = i[953];
  assign o[1112] = i[952];
  assign o[1111] = i[951];
  assign o[1110] = i[950];
  assign o[1109] = i[949];
  assign o[1108] = i[948];
  assign o[1107] = i[947];
  assign o[1106] = i[946];
  assign o[1105] = i[945];
  assign o[1104] = i[944];
  assign o[1103] = i[943];
  assign o[1102] = i[942];
  assign o[1101] = i[941];
  assign o[1100] = i[940];
  assign o[1099] = i[939];
  assign o[1098] = i[938];
  assign o[1097] = i[937];
  assign o[1096] = i[936];
  assign o[1095] = i[935];
  assign o[1094] = i[934];
  assign o[1093] = i[933];
  assign o[1092] = i[932];
  assign o[1091] = i[931];
  assign o[1090] = i[930];
  assign o[1089] = i[929];
  assign o[1088] = i[928];
  assign o[1087] = i[991];
  assign o[1086] = i[990];
  assign o[1085] = i[989];
  assign o[1084] = i[988];
  assign o[1083] = i[987];
  assign o[1082] = i[986];
  assign o[1081] = i[985];
  assign o[1080] = i[984];
  assign o[1079] = i[983];
  assign o[1078] = i[982];
  assign o[1077] = i[981];
  assign o[1076] = i[980];
  assign o[1075] = i[979];
  assign o[1074] = i[978];
  assign o[1073] = i[977];
  assign o[1072] = i[976];
  assign o[1071] = i[975];
  assign o[1070] = i[974];
  assign o[1069] = i[973];
  assign o[1068] = i[972];
  assign o[1067] = i[971];
  assign o[1066] = i[970];
  assign o[1065] = i[969];
  assign o[1064] = i[968];
  assign o[1063] = i[967];
  assign o[1062] = i[966];
  assign o[1061] = i[965];
  assign o[1060] = i[964];
  assign o[1059] = i[963];
  assign o[1058] = i[962];
  assign o[1057] = i[961];
  assign o[1056] = i[960];
  assign o[1055] = i[1023];
  assign o[1054] = i[1022];
  assign o[1053] = i[1021];
  assign o[1052] = i[1020];
  assign o[1051] = i[1019];
  assign o[1050] = i[1018];
  assign o[1049] = i[1017];
  assign o[1048] = i[1016];
  assign o[1047] = i[1015];
  assign o[1046] = i[1014];
  assign o[1045] = i[1013];
  assign o[1044] = i[1012];
  assign o[1043] = i[1011];
  assign o[1042] = i[1010];
  assign o[1041] = i[1009];
  assign o[1040] = i[1008];
  assign o[1039] = i[1007];
  assign o[1038] = i[1006];
  assign o[1037] = i[1005];
  assign o[1036] = i[1004];
  assign o[1035] = i[1003];
  assign o[1034] = i[1002];
  assign o[1033] = i[1001];
  assign o[1032] = i[1000];
  assign o[1031] = i[999];
  assign o[1030] = i[998];
  assign o[1029] = i[997];
  assign o[1028] = i[996];
  assign o[1027] = i[995];
  assign o[1026] = i[994];
  assign o[1025] = i[993];
  assign o[1024] = i[992];
  assign o[1023] = i[1055];
  assign o[1022] = i[1054];
  assign o[1021] = i[1053];
  assign o[1020] = i[1052];
  assign o[1019] = i[1051];
  assign o[1018] = i[1050];
  assign o[1017] = i[1049];
  assign o[1016] = i[1048];
  assign o[1015] = i[1047];
  assign o[1014] = i[1046];
  assign o[1013] = i[1045];
  assign o[1012] = i[1044];
  assign o[1011] = i[1043];
  assign o[1010] = i[1042];
  assign o[1009] = i[1041];
  assign o[1008] = i[1040];
  assign o[1007] = i[1039];
  assign o[1006] = i[1038];
  assign o[1005] = i[1037];
  assign o[1004] = i[1036];
  assign o[1003] = i[1035];
  assign o[1002] = i[1034];
  assign o[1001] = i[1033];
  assign o[1000] = i[1032];
  assign o[999] = i[1031];
  assign o[998] = i[1030];
  assign o[997] = i[1029];
  assign o[996] = i[1028];
  assign o[995] = i[1027];
  assign o[994] = i[1026];
  assign o[993] = i[1025];
  assign o[992] = i[1024];
  assign o[991] = i[1087];
  assign o[990] = i[1086];
  assign o[989] = i[1085];
  assign o[988] = i[1084];
  assign o[987] = i[1083];
  assign o[986] = i[1082];
  assign o[985] = i[1081];
  assign o[984] = i[1080];
  assign o[983] = i[1079];
  assign o[982] = i[1078];
  assign o[981] = i[1077];
  assign o[980] = i[1076];
  assign o[979] = i[1075];
  assign o[978] = i[1074];
  assign o[977] = i[1073];
  assign o[976] = i[1072];
  assign o[975] = i[1071];
  assign o[974] = i[1070];
  assign o[973] = i[1069];
  assign o[972] = i[1068];
  assign o[971] = i[1067];
  assign o[970] = i[1066];
  assign o[969] = i[1065];
  assign o[968] = i[1064];
  assign o[967] = i[1063];
  assign o[966] = i[1062];
  assign o[965] = i[1061];
  assign o[964] = i[1060];
  assign o[963] = i[1059];
  assign o[962] = i[1058];
  assign o[961] = i[1057];
  assign o[960] = i[1056];
  assign o[959] = i[1119];
  assign o[958] = i[1118];
  assign o[957] = i[1117];
  assign o[956] = i[1116];
  assign o[955] = i[1115];
  assign o[954] = i[1114];
  assign o[953] = i[1113];
  assign o[952] = i[1112];
  assign o[951] = i[1111];
  assign o[950] = i[1110];
  assign o[949] = i[1109];
  assign o[948] = i[1108];
  assign o[947] = i[1107];
  assign o[946] = i[1106];
  assign o[945] = i[1105];
  assign o[944] = i[1104];
  assign o[943] = i[1103];
  assign o[942] = i[1102];
  assign o[941] = i[1101];
  assign o[940] = i[1100];
  assign o[939] = i[1099];
  assign o[938] = i[1098];
  assign o[937] = i[1097];
  assign o[936] = i[1096];
  assign o[935] = i[1095];
  assign o[934] = i[1094];
  assign o[933] = i[1093];
  assign o[932] = i[1092];
  assign o[931] = i[1091];
  assign o[930] = i[1090];
  assign o[929] = i[1089];
  assign o[928] = i[1088];
  assign o[927] = i[1151];
  assign o[926] = i[1150];
  assign o[925] = i[1149];
  assign o[924] = i[1148];
  assign o[923] = i[1147];
  assign o[922] = i[1146];
  assign o[921] = i[1145];
  assign o[920] = i[1144];
  assign o[919] = i[1143];
  assign o[918] = i[1142];
  assign o[917] = i[1141];
  assign o[916] = i[1140];
  assign o[915] = i[1139];
  assign o[914] = i[1138];
  assign o[913] = i[1137];
  assign o[912] = i[1136];
  assign o[911] = i[1135];
  assign o[910] = i[1134];
  assign o[909] = i[1133];
  assign o[908] = i[1132];
  assign o[907] = i[1131];
  assign o[906] = i[1130];
  assign o[905] = i[1129];
  assign o[904] = i[1128];
  assign o[903] = i[1127];
  assign o[902] = i[1126];
  assign o[901] = i[1125];
  assign o[900] = i[1124];
  assign o[899] = i[1123];
  assign o[898] = i[1122];
  assign o[897] = i[1121];
  assign o[896] = i[1120];
  assign o[895] = i[1183];
  assign o[894] = i[1182];
  assign o[893] = i[1181];
  assign o[892] = i[1180];
  assign o[891] = i[1179];
  assign o[890] = i[1178];
  assign o[889] = i[1177];
  assign o[888] = i[1176];
  assign o[887] = i[1175];
  assign o[886] = i[1174];
  assign o[885] = i[1173];
  assign o[884] = i[1172];
  assign o[883] = i[1171];
  assign o[882] = i[1170];
  assign o[881] = i[1169];
  assign o[880] = i[1168];
  assign o[879] = i[1167];
  assign o[878] = i[1166];
  assign o[877] = i[1165];
  assign o[876] = i[1164];
  assign o[875] = i[1163];
  assign o[874] = i[1162];
  assign o[873] = i[1161];
  assign o[872] = i[1160];
  assign o[871] = i[1159];
  assign o[870] = i[1158];
  assign o[869] = i[1157];
  assign o[868] = i[1156];
  assign o[867] = i[1155];
  assign o[866] = i[1154];
  assign o[865] = i[1153];
  assign o[864] = i[1152];
  assign o[863] = i[1215];
  assign o[862] = i[1214];
  assign o[861] = i[1213];
  assign o[860] = i[1212];
  assign o[859] = i[1211];
  assign o[858] = i[1210];
  assign o[857] = i[1209];
  assign o[856] = i[1208];
  assign o[855] = i[1207];
  assign o[854] = i[1206];
  assign o[853] = i[1205];
  assign o[852] = i[1204];
  assign o[851] = i[1203];
  assign o[850] = i[1202];
  assign o[849] = i[1201];
  assign o[848] = i[1200];
  assign o[847] = i[1199];
  assign o[846] = i[1198];
  assign o[845] = i[1197];
  assign o[844] = i[1196];
  assign o[843] = i[1195];
  assign o[842] = i[1194];
  assign o[841] = i[1193];
  assign o[840] = i[1192];
  assign o[839] = i[1191];
  assign o[838] = i[1190];
  assign o[837] = i[1189];
  assign o[836] = i[1188];
  assign o[835] = i[1187];
  assign o[834] = i[1186];
  assign o[833] = i[1185];
  assign o[832] = i[1184];
  assign o[831] = i[1247];
  assign o[830] = i[1246];
  assign o[829] = i[1245];
  assign o[828] = i[1244];
  assign o[827] = i[1243];
  assign o[826] = i[1242];
  assign o[825] = i[1241];
  assign o[824] = i[1240];
  assign o[823] = i[1239];
  assign o[822] = i[1238];
  assign o[821] = i[1237];
  assign o[820] = i[1236];
  assign o[819] = i[1235];
  assign o[818] = i[1234];
  assign o[817] = i[1233];
  assign o[816] = i[1232];
  assign o[815] = i[1231];
  assign o[814] = i[1230];
  assign o[813] = i[1229];
  assign o[812] = i[1228];
  assign o[811] = i[1227];
  assign o[810] = i[1226];
  assign o[809] = i[1225];
  assign o[808] = i[1224];
  assign o[807] = i[1223];
  assign o[806] = i[1222];
  assign o[805] = i[1221];
  assign o[804] = i[1220];
  assign o[803] = i[1219];
  assign o[802] = i[1218];
  assign o[801] = i[1217];
  assign o[800] = i[1216];
  assign o[799] = i[1279];
  assign o[798] = i[1278];
  assign o[797] = i[1277];
  assign o[796] = i[1276];
  assign o[795] = i[1275];
  assign o[794] = i[1274];
  assign o[793] = i[1273];
  assign o[792] = i[1272];
  assign o[791] = i[1271];
  assign o[790] = i[1270];
  assign o[789] = i[1269];
  assign o[788] = i[1268];
  assign o[787] = i[1267];
  assign o[786] = i[1266];
  assign o[785] = i[1265];
  assign o[784] = i[1264];
  assign o[783] = i[1263];
  assign o[782] = i[1262];
  assign o[781] = i[1261];
  assign o[780] = i[1260];
  assign o[779] = i[1259];
  assign o[778] = i[1258];
  assign o[777] = i[1257];
  assign o[776] = i[1256];
  assign o[775] = i[1255];
  assign o[774] = i[1254];
  assign o[773] = i[1253];
  assign o[772] = i[1252];
  assign o[771] = i[1251];
  assign o[770] = i[1250];
  assign o[769] = i[1249];
  assign o[768] = i[1248];
  assign o[767] = i[1311];
  assign o[766] = i[1310];
  assign o[765] = i[1309];
  assign o[764] = i[1308];
  assign o[763] = i[1307];
  assign o[762] = i[1306];
  assign o[761] = i[1305];
  assign o[760] = i[1304];
  assign o[759] = i[1303];
  assign o[758] = i[1302];
  assign o[757] = i[1301];
  assign o[756] = i[1300];
  assign o[755] = i[1299];
  assign o[754] = i[1298];
  assign o[753] = i[1297];
  assign o[752] = i[1296];
  assign o[751] = i[1295];
  assign o[750] = i[1294];
  assign o[749] = i[1293];
  assign o[748] = i[1292];
  assign o[747] = i[1291];
  assign o[746] = i[1290];
  assign o[745] = i[1289];
  assign o[744] = i[1288];
  assign o[743] = i[1287];
  assign o[742] = i[1286];
  assign o[741] = i[1285];
  assign o[740] = i[1284];
  assign o[739] = i[1283];
  assign o[738] = i[1282];
  assign o[737] = i[1281];
  assign o[736] = i[1280];
  assign o[735] = i[1343];
  assign o[734] = i[1342];
  assign o[733] = i[1341];
  assign o[732] = i[1340];
  assign o[731] = i[1339];
  assign o[730] = i[1338];
  assign o[729] = i[1337];
  assign o[728] = i[1336];
  assign o[727] = i[1335];
  assign o[726] = i[1334];
  assign o[725] = i[1333];
  assign o[724] = i[1332];
  assign o[723] = i[1331];
  assign o[722] = i[1330];
  assign o[721] = i[1329];
  assign o[720] = i[1328];
  assign o[719] = i[1327];
  assign o[718] = i[1326];
  assign o[717] = i[1325];
  assign o[716] = i[1324];
  assign o[715] = i[1323];
  assign o[714] = i[1322];
  assign o[713] = i[1321];
  assign o[712] = i[1320];
  assign o[711] = i[1319];
  assign o[710] = i[1318];
  assign o[709] = i[1317];
  assign o[708] = i[1316];
  assign o[707] = i[1315];
  assign o[706] = i[1314];
  assign o[705] = i[1313];
  assign o[704] = i[1312];
  assign o[703] = i[1375];
  assign o[702] = i[1374];
  assign o[701] = i[1373];
  assign o[700] = i[1372];
  assign o[699] = i[1371];
  assign o[698] = i[1370];
  assign o[697] = i[1369];
  assign o[696] = i[1368];
  assign o[695] = i[1367];
  assign o[694] = i[1366];
  assign o[693] = i[1365];
  assign o[692] = i[1364];
  assign o[691] = i[1363];
  assign o[690] = i[1362];
  assign o[689] = i[1361];
  assign o[688] = i[1360];
  assign o[687] = i[1359];
  assign o[686] = i[1358];
  assign o[685] = i[1357];
  assign o[684] = i[1356];
  assign o[683] = i[1355];
  assign o[682] = i[1354];
  assign o[681] = i[1353];
  assign o[680] = i[1352];
  assign o[679] = i[1351];
  assign o[678] = i[1350];
  assign o[677] = i[1349];
  assign o[676] = i[1348];
  assign o[675] = i[1347];
  assign o[674] = i[1346];
  assign o[673] = i[1345];
  assign o[672] = i[1344];
  assign o[671] = i[1407];
  assign o[670] = i[1406];
  assign o[669] = i[1405];
  assign o[668] = i[1404];
  assign o[667] = i[1403];
  assign o[666] = i[1402];
  assign o[665] = i[1401];
  assign o[664] = i[1400];
  assign o[663] = i[1399];
  assign o[662] = i[1398];
  assign o[661] = i[1397];
  assign o[660] = i[1396];
  assign o[659] = i[1395];
  assign o[658] = i[1394];
  assign o[657] = i[1393];
  assign o[656] = i[1392];
  assign o[655] = i[1391];
  assign o[654] = i[1390];
  assign o[653] = i[1389];
  assign o[652] = i[1388];
  assign o[651] = i[1387];
  assign o[650] = i[1386];
  assign o[649] = i[1385];
  assign o[648] = i[1384];
  assign o[647] = i[1383];
  assign o[646] = i[1382];
  assign o[645] = i[1381];
  assign o[644] = i[1380];
  assign o[643] = i[1379];
  assign o[642] = i[1378];
  assign o[641] = i[1377];
  assign o[640] = i[1376];
  assign o[639] = i[1439];
  assign o[638] = i[1438];
  assign o[637] = i[1437];
  assign o[636] = i[1436];
  assign o[635] = i[1435];
  assign o[634] = i[1434];
  assign o[633] = i[1433];
  assign o[632] = i[1432];
  assign o[631] = i[1431];
  assign o[630] = i[1430];
  assign o[629] = i[1429];
  assign o[628] = i[1428];
  assign o[627] = i[1427];
  assign o[626] = i[1426];
  assign o[625] = i[1425];
  assign o[624] = i[1424];
  assign o[623] = i[1423];
  assign o[622] = i[1422];
  assign o[621] = i[1421];
  assign o[620] = i[1420];
  assign o[619] = i[1419];
  assign o[618] = i[1418];
  assign o[617] = i[1417];
  assign o[616] = i[1416];
  assign o[615] = i[1415];
  assign o[614] = i[1414];
  assign o[613] = i[1413];
  assign o[612] = i[1412];
  assign o[611] = i[1411];
  assign o[610] = i[1410];
  assign o[609] = i[1409];
  assign o[608] = i[1408];
  assign o[607] = i[1471];
  assign o[606] = i[1470];
  assign o[605] = i[1469];
  assign o[604] = i[1468];
  assign o[603] = i[1467];
  assign o[602] = i[1466];
  assign o[601] = i[1465];
  assign o[600] = i[1464];
  assign o[599] = i[1463];
  assign o[598] = i[1462];
  assign o[597] = i[1461];
  assign o[596] = i[1460];
  assign o[595] = i[1459];
  assign o[594] = i[1458];
  assign o[593] = i[1457];
  assign o[592] = i[1456];
  assign o[591] = i[1455];
  assign o[590] = i[1454];
  assign o[589] = i[1453];
  assign o[588] = i[1452];
  assign o[587] = i[1451];
  assign o[586] = i[1450];
  assign o[585] = i[1449];
  assign o[584] = i[1448];
  assign o[583] = i[1447];
  assign o[582] = i[1446];
  assign o[581] = i[1445];
  assign o[580] = i[1444];
  assign o[579] = i[1443];
  assign o[578] = i[1442];
  assign o[577] = i[1441];
  assign o[576] = i[1440];
  assign o[575] = i[1503];
  assign o[574] = i[1502];
  assign o[573] = i[1501];
  assign o[572] = i[1500];
  assign o[571] = i[1499];
  assign o[570] = i[1498];
  assign o[569] = i[1497];
  assign o[568] = i[1496];
  assign o[567] = i[1495];
  assign o[566] = i[1494];
  assign o[565] = i[1493];
  assign o[564] = i[1492];
  assign o[563] = i[1491];
  assign o[562] = i[1490];
  assign o[561] = i[1489];
  assign o[560] = i[1488];
  assign o[559] = i[1487];
  assign o[558] = i[1486];
  assign o[557] = i[1485];
  assign o[556] = i[1484];
  assign o[555] = i[1483];
  assign o[554] = i[1482];
  assign o[553] = i[1481];
  assign o[552] = i[1480];
  assign o[551] = i[1479];
  assign o[550] = i[1478];
  assign o[549] = i[1477];
  assign o[548] = i[1476];
  assign o[547] = i[1475];
  assign o[546] = i[1474];
  assign o[545] = i[1473];
  assign o[544] = i[1472];
  assign o[543] = i[1535];
  assign o[542] = i[1534];
  assign o[541] = i[1533];
  assign o[540] = i[1532];
  assign o[539] = i[1531];
  assign o[538] = i[1530];
  assign o[537] = i[1529];
  assign o[536] = i[1528];
  assign o[535] = i[1527];
  assign o[534] = i[1526];
  assign o[533] = i[1525];
  assign o[532] = i[1524];
  assign o[531] = i[1523];
  assign o[530] = i[1522];
  assign o[529] = i[1521];
  assign o[528] = i[1520];
  assign o[527] = i[1519];
  assign o[526] = i[1518];
  assign o[525] = i[1517];
  assign o[524] = i[1516];
  assign o[523] = i[1515];
  assign o[522] = i[1514];
  assign o[521] = i[1513];
  assign o[520] = i[1512];
  assign o[519] = i[1511];
  assign o[518] = i[1510];
  assign o[517] = i[1509];
  assign o[516] = i[1508];
  assign o[515] = i[1507];
  assign o[514] = i[1506];
  assign o[513] = i[1505];
  assign o[512] = i[1504];
  assign o[511] = i[1567];
  assign o[510] = i[1566];
  assign o[509] = i[1565];
  assign o[508] = i[1564];
  assign o[507] = i[1563];
  assign o[506] = i[1562];
  assign o[505] = i[1561];
  assign o[504] = i[1560];
  assign o[503] = i[1559];
  assign o[502] = i[1558];
  assign o[501] = i[1557];
  assign o[500] = i[1556];
  assign o[499] = i[1555];
  assign o[498] = i[1554];
  assign o[497] = i[1553];
  assign o[496] = i[1552];
  assign o[495] = i[1551];
  assign o[494] = i[1550];
  assign o[493] = i[1549];
  assign o[492] = i[1548];
  assign o[491] = i[1547];
  assign o[490] = i[1546];
  assign o[489] = i[1545];
  assign o[488] = i[1544];
  assign o[487] = i[1543];
  assign o[486] = i[1542];
  assign o[485] = i[1541];
  assign o[484] = i[1540];
  assign o[483] = i[1539];
  assign o[482] = i[1538];
  assign o[481] = i[1537];
  assign o[480] = i[1536];
  assign o[479] = i[1599];
  assign o[478] = i[1598];
  assign o[477] = i[1597];
  assign o[476] = i[1596];
  assign o[475] = i[1595];
  assign o[474] = i[1594];
  assign o[473] = i[1593];
  assign o[472] = i[1592];
  assign o[471] = i[1591];
  assign o[470] = i[1590];
  assign o[469] = i[1589];
  assign o[468] = i[1588];
  assign o[467] = i[1587];
  assign o[466] = i[1586];
  assign o[465] = i[1585];
  assign o[464] = i[1584];
  assign o[463] = i[1583];
  assign o[462] = i[1582];
  assign o[461] = i[1581];
  assign o[460] = i[1580];
  assign o[459] = i[1579];
  assign o[458] = i[1578];
  assign o[457] = i[1577];
  assign o[456] = i[1576];
  assign o[455] = i[1575];
  assign o[454] = i[1574];
  assign o[453] = i[1573];
  assign o[452] = i[1572];
  assign o[451] = i[1571];
  assign o[450] = i[1570];
  assign o[449] = i[1569];
  assign o[448] = i[1568];
  assign o[447] = i[1631];
  assign o[446] = i[1630];
  assign o[445] = i[1629];
  assign o[444] = i[1628];
  assign o[443] = i[1627];
  assign o[442] = i[1626];
  assign o[441] = i[1625];
  assign o[440] = i[1624];
  assign o[439] = i[1623];
  assign o[438] = i[1622];
  assign o[437] = i[1621];
  assign o[436] = i[1620];
  assign o[435] = i[1619];
  assign o[434] = i[1618];
  assign o[433] = i[1617];
  assign o[432] = i[1616];
  assign o[431] = i[1615];
  assign o[430] = i[1614];
  assign o[429] = i[1613];
  assign o[428] = i[1612];
  assign o[427] = i[1611];
  assign o[426] = i[1610];
  assign o[425] = i[1609];
  assign o[424] = i[1608];
  assign o[423] = i[1607];
  assign o[422] = i[1606];
  assign o[421] = i[1605];
  assign o[420] = i[1604];
  assign o[419] = i[1603];
  assign o[418] = i[1602];
  assign o[417] = i[1601];
  assign o[416] = i[1600];
  assign o[415] = i[1663];
  assign o[414] = i[1662];
  assign o[413] = i[1661];
  assign o[412] = i[1660];
  assign o[411] = i[1659];
  assign o[410] = i[1658];
  assign o[409] = i[1657];
  assign o[408] = i[1656];
  assign o[407] = i[1655];
  assign o[406] = i[1654];
  assign o[405] = i[1653];
  assign o[404] = i[1652];
  assign o[403] = i[1651];
  assign o[402] = i[1650];
  assign o[401] = i[1649];
  assign o[400] = i[1648];
  assign o[399] = i[1647];
  assign o[398] = i[1646];
  assign o[397] = i[1645];
  assign o[396] = i[1644];
  assign o[395] = i[1643];
  assign o[394] = i[1642];
  assign o[393] = i[1641];
  assign o[392] = i[1640];
  assign o[391] = i[1639];
  assign o[390] = i[1638];
  assign o[389] = i[1637];
  assign o[388] = i[1636];
  assign o[387] = i[1635];
  assign o[386] = i[1634];
  assign o[385] = i[1633];
  assign o[384] = i[1632];
  assign o[383] = i[1695];
  assign o[382] = i[1694];
  assign o[381] = i[1693];
  assign o[380] = i[1692];
  assign o[379] = i[1691];
  assign o[378] = i[1690];
  assign o[377] = i[1689];
  assign o[376] = i[1688];
  assign o[375] = i[1687];
  assign o[374] = i[1686];
  assign o[373] = i[1685];
  assign o[372] = i[1684];
  assign o[371] = i[1683];
  assign o[370] = i[1682];
  assign o[369] = i[1681];
  assign o[368] = i[1680];
  assign o[367] = i[1679];
  assign o[366] = i[1678];
  assign o[365] = i[1677];
  assign o[364] = i[1676];
  assign o[363] = i[1675];
  assign o[362] = i[1674];
  assign o[361] = i[1673];
  assign o[360] = i[1672];
  assign o[359] = i[1671];
  assign o[358] = i[1670];
  assign o[357] = i[1669];
  assign o[356] = i[1668];
  assign o[355] = i[1667];
  assign o[354] = i[1666];
  assign o[353] = i[1665];
  assign o[352] = i[1664];
  assign o[351] = i[1727];
  assign o[350] = i[1726];
  assign o[349] = i[1725];
  assign o[348] = i[1724];
  assign o[347] = i[1723];
  assign o[346] = i[1722];
  assign o[345] = i[1721];
  assign o[344] = i[1720];
  assign o[343] = i[1719];
  assign o[342] = i[1718];
  assign o[341] = i[1717];
  assign o[340] = i[1716];
  assign o[339] = i[1715];
  assign o[338] = i[1714];
  assign o[337] = i[1713];
  assign o[336] = i[1712];
  assign o[335] = i[1711];
  assign o[334] = i[1710];
  assign o[333] = i[1709];
  assign o[332] = i[1708];
  assign o[331] = i[1707];
  assign o[330] = i[1706];
  assign o[329] = i[1705];
  assign o[328] = i[1704];
  assign o[327] = i[1703];
  assign o[326] = i[1702];
  assign o[325] = i[1701];
  assign o[324] = i[1700];
  assign o[323] = i[1699];
  assign o[322] = i[1698];
  assign o[321] = i[1697];
  assign o[320] = i[1696];
  assign o[319] = i[1759];
  assign o[318] = i[1758];
  assign o[317] = i[1757];
  assign o[316] = i[1756];
  assign o[315] = i[1755];
  assign o[314] = i[1754];
  assign o[313] = i[1753];
  assign o[312] = i[1752];
  assign o[311] = i[1751];
  assign o[310] = i[1750];
  assign o[309] = i[1749];
  assign o[308] = i[1748];
  assign o[307] = i[1747];
  assign o[306] = i[1746];
  assign o[305] = i[1745];
  assign o[304] = i[1744];
  assign o[303] = i[1743];
  assign o[302] = i[1742];
  assign o[301] = i[1741];
  assign o[300] = i[1740];
  assign o[299] = i[1739];
  assign o[298] = i[1738];
  assign o[297] = i[1737];
  assign o[296] = i[1736];
  assign o[295] = i[1735];
  assign o[294] = i[1734];
  assign o[293] = i[1733];
  assign o[292] = i[1732];
  assign o[291] = i[1731];
  assign o[290] = i[1730];
  assign o[289] = i[1729];
  assign o[288] = i[1728];
  assign o[287] = i[1791];
  assign o[286] = i[1790];
  assign o[285] = i[1789];
  assign o[284] = i[1788];
  assign o[283] = i[1787];
  assign o[282] = i[1786];
  assign o[281] = i[1785];
  assign o[280] = i[1784];
  assign o[279] = i[1783];
  assign o[278] = i[1782];
  assign o[277] = i[1781];
  assign o[276] = i[1780];
  assign o[275] = i[1779];
  assign o[274] = i[1778];
  assign o[273] = i[1777];
  assign o[272] = i[1776];
  assign o[271] = i[1775];
  assign o[270] = i[1774];
  assign o[269] = i[1773];
  assign o[268] = i[1772];
  assign o[267] = i[1771];
  assign o[266] = i[1770];
  assign o[265] = i[1769];
  assign o[264] = i[1768];
  assign o[263] = i[1767];
  assign o[262] = i[1766];
  assign o[261] = i[1765];
  assign o[260] = i[1764];
  assign o[259] = i[1763];
  assign o[258] = i[1762];
  assign o[257] = i[1761];
  assign o[256] = i[1760];
  assign o[255] = i[1823];
  assign o[254] = i[1822];
  assign o[253] = i[1821];
  assign o[252] = i[1820];
  assign o[251] = i[1819];
  assign o[250] = i[1818];
  assign o[249] = i[1817];
  assign o[248] = i[1816];
  assign o[247] = i[1815];
  assign o[246] = i[1814];
  assign o[245] = i[1813];
  assign o[244] = i[1812];
  assign o[243] = i[1811];
  assign o[242] = i[1810];
  assign o[241] = i[1809];
  assign o[240] = i[1808];
  assign o[239] = i[1807];
  assign o[238] = i[1806];
  assign o[237] = i[1805];
  assign o[236] = i[1804];
  assign o[235] = i[1803];
  assign o[234] = i[1802];
  assign o[233] = i[1801];
  assign o[232] = i[1800];
  assign o[231] = i[1799];
  assign o[230] = i[1798];
  assign o[229] = i[1797];
  assign o[228] = i[1796];
  assign o[227] = i[1795];
  assign o[226] = i[1794];
  assign o[225] = i[1793];
  assign o[224] = i[1792];
  assign o[223] = i[1855];
  assign o[222] = i[1854];
  assign o[221] = i[1853];
  assign o[220] = i[1852];
  assign o[219] = i[1851];
  assign o[218] = i[1850];
  assign o[217] = i[1849];
  assign o[216] = i[1848];
  assign o[215] = i[1847];
  assign o[214] = i[1846];
  assign o[213] = i[1845];
  assign o[212] = i[1844];
  assign o[211] = i[1843];
  assign o[210] = i[1842];
  assign o[209] = i[1841];
  assign o[208] = i[1840];
  assign o[207] = i[1839];
  assign o[206] = i[1838];
  assign o[205] = i[1837];
  assign o[204] = i[1836];
  assign o[203] = i[1835];
  assign o[202] = i[1834];
  assign o[201] = i[1833];
  assign o[200] = i[1832];
  assign o[199] = i[1831];
  assign o[198] = i[1830];
  assign o[197] = i[1829];
  assign o[196] = i[1828];
  assign o[195] = i[1827];
  assign o[194] = i[1826];
  assign o[193] = i[1825];
  assign o[192] = i[1824];
  assign o[191] = i[1887];
  assign o[190] = i[1886];
  assign o[189] = i[1885];
  assign o[188] = i[1884];
  assign o[187] = i[1883];
  assign o[186] = i[1882];
  assign o[185] = i[1881];
  assign o[184] = i[1880];
  assign o[183] = i[1879];
  assign o[182] = i[1878];
  assign o[181] = i[1877];
  assign o[180] = i[1876];
  assign o[179] = i[1875];
  assign o[178] = i[1874];
  assign o[177] = i[1873];
  assign o[176] = i[1872];
  assign o[175] = i[1871];
  assign o[174] = i[1870];
  assign o[173] = i[1869];
  assign o[172] = i[1868];
  assign o[171] = i[1867];
  assign o[170] = i[1866];
  assign o[169] = i[1865];
  assign o[168] = i[1864];
  assign o[167] = i[1863];
  assign o[166] = i[1862];
  assign o[165] = i[1861];
  assign o[164] = i[1860];
  assign o[163] = i[1859];
  assign o[162] = i[1858];
  assign o[161] = i[1857];
  assign o[160] = i[1856];
  assign o[159] = i[1919];
  assign o[158] = i[1918];
  assign o[157] = i[1917];
  assign o[156] = i[1916];
  assign o[155] = i[1915];
  assign o[154] = i[1914];
  assign o[153] = i[1913];
  assign o[152] = i[1912];
  assign o[151] = i[1911];
  assign o[150] = i[1910];
  assign o[149] = i[1909];
  assign o[148] = i[1908];
  assign o[147] = i[1907];
  assign o[146] = i[1906];
  assign o[145] = i[1905];
  assign o[144] = i[1904];
  assign o[143] = i[1903];
  assign o[142] = i[1902];
  assign o[141] = i[1901];
  assign o[140] = i[1900];
  assign o[139] = i[1899];
  assign o[138] = i[1898];
  assign o[137] = i[1897];
  assign o[136] = i[1896];
  assign o[135] = i[1895];
  assign o[134] = i[1894];
  assign o[133] = i[1893];
  assign o[132] = i[1892];
  assign o[131] = i[1891];
  assign o[130] = i[1890];
  assign o[129] = i[1889];
  assign o[128] = i[1888];
  assign o[127] = i[1951];
  assign o[126] = i[1950];
  assign o[125] = i[1949];
  assign o[124] = i[1948];
  assign o[123] = i[1947];
  assign o[122] = i[1946];
  assign o[121] = i[1945];
  assign o[120] = i[1944];
  assign o[119] = i[1943];
  assign o[118] = i[1942];
  assign o[117] = i[1941];
  assign o[116] = i[1940];
  assign o[115] = i[1939];
  assign o[114] = i[1938];
  assign o[113] = i[1937];
  assign o[112] = i[1936];
  assign o[111] = i[1935];
  assign o[110] = i[1934];
  assign o[109] = i[1933];
  assign o[108] = i[1932];
  assign o[107] = i[1931];
  assign o[106] = i[1930];
  assign o[105] = i[1929];
  assign o[104] = i[1928];
  assign o[103] = i[1927];
  assign o[102] = i[1926];
  assign o[101] = i[1925];
  assign o[100] = i[1924];
  assign o[99] = i[1923];
  assign o[98] = i[1922];
  assign o[97] = i[1921];
  assign o[96] = i[1920];
  assign o[95] = i[1983];
  assign o[94] = i[1982];
  assign o[93] = i[1981];
  assign o[92] = i[1980];
  assign o[91] = i[1979];
  assign o[90] = i[1978];
  assign o[89] = i[1977];
  assign o[88] = i[1976];
  assign o[87] = i[1975];
  assign o[86] = i[1974];
  assign o[85] = i[1973];
  assign o[84] = i[1972];
  assign o[83] = i[1971];
  assign o[82] = i[1970];
  assign o[81] = i[1969];
  assign o[80] = i[1968];
  assign o[79] = i[1967];
  assign o[78] = i[1966];
  assign o[77] = i[1965];
  assign o[76] = i[1964];
  assign o[75] = i[1963];
  assign o[74] = i[1962];
  assign o[73] = i[1961];
  assign o[72] = i[1960];
  assign o[71] = i[1959];
  assign o[70] = i[1958];
  assign o[69] = i[1957];
  assign o[68] = i[1956];
  assign o[67] = i[1955];
  assign o[66] = i[1954];
  assign o[65] = i[1953];
  assign o[64] = i[1952];
  assign o[63] = i[2015];
  assign o[62] = i[2014];
  assign o[61] = i[2013];
  assign o[60] = i[2012];
  assign o[59] = i[2011];
  assign o[58] = i[2010];
  assign o[57] = i[2009];
  assign o[56] = i[2008];
  assign o[55] = i[2007];
  assign o[54] = i[2006];
  assign o[53] = i[2005];
  assign o[52] = i[2004];
  assign o[51] = i[2003];
  assign o[50] = i[2002];
  assign o[49] = i[2001];
  assign o[48] = i[2000];
  assign o[47] = i[1999];
  assign o[46] = i[1998];
  assign o[45] = i[1997];
  assign o[44] = i[1996];
  assign o[43] = i[1995];
  assign o[42] = i[1994];
  assign o[41] = i[1993];
  assign o[40] = i[1992];
  assign o[39] = i[1991];
  assign o[38] = i[1990];
  assign o[37] = i[1989];
  assign o[36] = i[1988];
  assign o[35] = i[1987];
  assign o[34] = i[1986];
  assign o[33] = i[1985];
  assign o[32] = i[1984];
  assign o[31] = i[2047];
  assign o[30] = i[2046];
  assign o[29] = i[2045];
  assign o[28] = i[2044];
  assign o[27] = i[2043];
  assign o[26] = i[2042];
  assign o[25] = i[2041];
  assign o[24] = i[2040];
  assign o[23] = i[2039];
  assign o[22] = i[2038];
  assign o[21] = i[2037];
  assign o[20] = i[2036];
  assign o[19] = i[2035];
  assign o[18] = i[2034];
  assign o[17] = i[2033];
  assign o[16] = i[2032];
  assign o[15] = i[2031];
  assign o[14] = i[2030];
  assign o[13] = i[2029];
  assign o[12] = i[2028];
  assign o[11] = i[2027];
  assign o[10] = i[2026];
  assign o[9] = i[2025];
  assign o[8] = i[2024];
  assign o[7] = i[2023];
  assign o[6] = i[2022];
  assign o[5] = i[2021];
  assign o[4] = i[2020];
  assign o[3] = i[2019];
  assign o[2] = i[2018];
  assign o[1] = i[2017];
  assign o[0] = i[2016];

endmodule



module bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  wire [63:0] \nz.mem ;
  reg \nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,
  \nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,\nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,
  \nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,
  \nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,
  \nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,
  \nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,
  \nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,\nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,
  \nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,\nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,
  \nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,
  \nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,
  \nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,
  \nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,
  \nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,\nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,
  \nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,
  \nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,
  \nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,
  \nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[31] = (N3)? \nz.mem [31] : 
                        (N0)? \nz.mem [63] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[30] = (N3)? \nz.mem [30] : 
                        (N0)? \nz.mem [62] : 1'b0;
  assign r_data_o[29] = (N3)? \nz.mem [29] : 
                        (N0)? \nz.mem [61] : 1'b0;
  assign r_data_o[28] = (N3)? \nz.mem [28] : 
                        (N0)? \nz.mem [60] : 1'b0;
  assign r_data_o[27] = (N3)? \nz.mem [27] : 
                        (N0)? \nz.mem [59] : 1'b0;
  assign r_data_o[26] = (N3)? \nz.mem [26] : 
                        (N0)? \nz.mem [58] : 1'b0;
  assign r_data_o[25] = (N3)? \nz.mem [25] : 
                        (N0)? \nz.mem [57] : 1'b0;
  assign r_data_o[24] = (N3)? \nz.mem [24] : 
                        (N0)? \nz.mem [56] : 1'b0;
  assign r_data_o[23] = (N3)? \nz.mem [23] : 
                        (N0)? \nz.mem [55] : 1'b0;
  assign r_data_o[22] = (N3)? \nz.mem [22] : 
                        (N0)? \nz.mem [54] : 1'b0;
  assign r_data_o[21] = (N3)? \nz.mem [21] : 
                        (N0)? \nz.mem [53] : 1'b0;
  assign r_data_o[20] = (N3)? \nz.mem [20] : 
                        (N0)? \nz.mem [52] : 1'b0;
  assign r_data_o[19] = (N3)? \nz.mem [19] : 
                        (N0)? \nz.mem [51] : 1'b0;
  assign r_data_o[18] = (N3)? \nz.mem [18] : 
                        (N0)? \nz.mem [50] : 1'b0;
  assign r_data_o[17] = (N3)? \nz.mem [17] : 
                        (N0)? \nz.mem [49] : 1'b0;
  assign r_data_o[16] = (N3)? \nz.mem [16] : 
                        (N0)? \nz.mem [48] : 1'b0;
  assign r_data_o[15] = (N3)? \nz.mem [15] : 
                        (N0)? \nz.mem [47] : 1'b0;
  assign r_data_o[14] = (N3)? \nz.mem [14] : 
                        (N0)? \nz.mem [46] : 1'b0;
  assign r_data_o[13] = (N3)? \nz.mem [13] : 
                        (N0)? \nz.mem [45] : 1'b0;
  assign r_data_o[12] = (N3)? \nz.mem [12] : 
                        (N0)? \nz.mem [44] : 1'b0;
  assign r_data_o[11] = (N3)? \nz.mem [11] : 
                        (N0)? \nz.mem [43] : 1'b0;
  assign r_data_o[10] = (N3)? \nz.mem [10] : 
                        (N0)? \nz.mem [42] : 1'b0;
  assign r_data_o[9] = (N3)? \nz.mem [9] : 
                       (N0)? \nz.mem [41] : 1'b0;
  assign r_data_o[8] = (N3)? \nz.mem [8] : 
                       (N0)? \nz.mem [40] : 1'b0;
  assign r_data_o[7] = (N3)? \nz.mem [7] : 
                       (N0)? \nz.mem [39] : 1'b0;
  assign r_data_o[6] = (N3)? \nz.mem [6] : 
                       (N0)? \nz.mem [38] : 1'b0;
  assign r_data_o[5] = (N3)? \nz.mem [5] : 
                       (N0)? \nz.mem [37] : 1'b0;
  assign r_data_o[4] = (N3)? \nz.mem [4] : 
                       (N0)? \nz.mem [36] : 1'b0;
  assign r_data_o[3] = (N3)? \nz.mem [3] : 
                       (N0)? \nz.mem [35] : 1'b0;
  assign r_data_o[2] = (N3)? \nz.mem [2] : 
                       (N0)? \nz.mem [34] : 1'b0;
  assign r_data_o[1] = (N3)? \nz.mem [1] : 
                       (N0)? \nz.mem [33] : 1'b0;
  assign r_data_o[0] = (N3)? \nz.mem [0] : 
                       (N0)? \nz.mem [32] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      \nz.mem_63_sv2v_reg  <= w_data_i[31];
      \nz.mem_62_sv2v_reg  <= w_data_i[30];
      \nz.mem_61_sv2v_reg  <= w_data_i[29];
      \nz.mem_60_sv2v_reg  <= w_data_i[28];
      \nz.mem_59_sv2v_reg  <= w_data_i[27];
      \nz.mem_58_sv2v_reg  <= w_data_i[26];
      \nz.mem_57_sv2v_reg  <= w_data_i[25];
      \nz.mem_56_sv2v_reg  <= w_data_i[24];
      \nz.mem_55_sv2v_reg  <= w_data_i[23];
      \nz.mem_54_sv2v_reg  <= w_data_i[22];
      \nz.mem_53_sv2v_reg  <= w_data_i[21];
      \nz.mem_52_sv2v_reg  <= w_data_i[20];
      \nz.mem_51_sv2v_reg  <= w_data_i[19];
      \nz.mem_50_sv2v_reg  <= w_data_i[18];
      \nz.mem_49_sv2v_reg  <= w_data_i[17];
      \nz.mem_48_sv2v_reg  <= w_data_i[16];
      \nz.mem_47_sv2v_reg  <= w_data_i[15];
      \nz.mem_46_sv2v_reg  <= w_data_i[14];
      \nz.mem_45_sv2v_reg  <= w_data_i[13];
      \nz.mem_44_sv2v_reg  <= w_data_i[12];
      \nz.mem_43_sv2v_reg  <= w_data_i[11];
      \nz.mem_42_sv2v_reg  <= w_data_i[10];
      \nz.mem_41_sv2v_reg  <= w_data_i[9];
      \nz.mem_40_sv2v_reg  <= w_data_i[8];
      \nz.mem_39_sv2v_reg  <= w_data_i[7];
      \nz.mem_38_sv2v_reg  <= w_data_i[6];
      \nz.mem_37_sv2v_reg  <= w_data_i[5];
      \nz.mem_36_sv2v_reg  <= w_data_i[4];
      \nz.mem_35_sv2v_reg  <= w_data_i[3];
      \nz.mem_34_sv2v_reg  <= w_data_i[2];
      \nz.mem_33_sv2v_reg  <= w_data_i[1];
      \nz.mem_32_sv2v_reg  <= w_data_i[0];
    end 
    if(N7) begin
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;

  bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p32
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,enq_i,tail_r,_0_net_,head_r,empty_r,full_r,N0,N1,N2,N3,N4,N5,N6,N7,
  N8,N9,N10,N11,N12,N13,N14;
  reg full_r_sv2v_reg,tail_r_sv2v_reg,head_r_sv2v_reg,empty_r_sv2v_reg;
  assign full_r = full_r_sv2v_reg;
  assign tail_r = tail_r_sv2v_reg;
  assign head_r = head_r_sv2v_reg;
  assign empty_r = empty_r_sv2v_reg;

  bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign _0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N5;
  assign N5 = ~full_r;
  assign N1 = enq_i;
  assign N0 = ~tail_r;
  assign N2 = ~head_r;
  assign N3 = N7 | N9;
  assign N7 = empty_r & N6;
  assign N6 = ~enq_i;
  assign N9 = N8 & N6;
  assign N8 = N5 & yumi_i;
  assign N4 = N13 | N14;
  assign N13 = N11 & N12;
  assign N11 = N10 & enq_i;
  assign N10 = ~empty_r;
  assign N12 = ~yumi_i;
  assign N14 = full_r & N12;

  always @(posedge clk_i) begin
    if(reset_i) begin
      full_r_sv2v_reg <= 1'b0;
      empty_r_sv2v_reg <= 1'b1;
    end else if(1'b1) begin
      full_r_sv2v_reg <= N4;
      empty_r_sv2v_reg <= N3;
    end 
    if(reset_i) begin
      tail_r_sv2v_reg <= 1'b0;
    end else if(N1) begin
      tail_r_sv2v_reg <= N0;
    end 
    if(reset_i) begin
      head_r_sv2v_reg <= 1'b0;
    end else if(yumi_i) begin
      head_r_sv2v_reg <= N2;
    end 
  end


endmodule



module bsg_parallel_in_serial_out
(
  clk_i,
  reset_i,
  valid_i,
  data_i,
  ready_and_o,
  valid_o,
  data_o,
  yumi_i
);

  input [2047:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input valid_i;
  input yumi_i;
  output ready_and_o;
  output valid_o;
  wire [31:0] data_o;
  wire ready_and_o,valid_o,fifo0_ready_lo,fifo_v_li,fifo0_yumi_li,
  \piso.fifo1_ready_lo ,\piso.fifo1_yumi_li ,_0_net_,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16;
  wire [2047:0] data_li,fifo_data_lo;
  wire [5:0] \piso.shift_ctr_r ;

  bsg_array_reverse_width_p32_els_p64
  \hi2lo.bar 
  (
    .i(data_i),
    .o(data_li)
  );


  bsg_two_fifo_width_p32
  \two_fifo.fifo0 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(fifo0_ready_lo),
    .data_i(data_li[2047:2016]),
    .v_i(fifo_v_li),
    .v_o(valid_o),
    .data_o(fifo_data_lo[2047:2016]),
    .yumi_i(fifo0_yumi_li)
  );


  bsg_one_fifo
  \piso.fifo1 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(\piso.fifo1_ready_lo ),
    .data_i(data_li[2015:0]),
    .v_i(fifo_v_li),
    .data_o(fifo_data_lo[2015:0]),
    .yumi_i(\piso.fifo1_yumi_li )
  );


  bsg_counter_clear_up
  \piso.shift_ctr 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(fifo0_yumi_li),
    .up_i(_0_net_),
    .count_o(\piso.shift_ctr_r )
  );


  bsg_mux
  \piso.data_o_mux 
  (
    .data_i(fifo_data_lo),
    .sel_i(\piso.shift_ctr_r ),
    .data_o(data_o)
  );

  assign N0 = ~\piso.shift_ctr_r [5];
  assign N1 = ~\piso.shift_ctr_r [4];
  assign N2 = ~\piso.shift_ctr_r [3];
  assign N3 = ~\piso.shift_ctr_r [2];
  assign N4 = ~\piso.shift_ctr_r [1];
  assign N5 = N1 | N0;
  assign N6 = N2 | N5;
  assign N7 = N3 | N6;
  assign N8 = N4 | N7;
  assign N9 = \piso.shift_ctr_r [0] | N8;
  assign N10 = ~N9;
  assign N11 = \piso.shift_ctr_r [4] & \piso.shift_ctr_r [5];
  assign N12 = \piso.shift_ctr_r [3] & N11;
  assign N13 = \piso.shift_ctr_r [2] & N12;
  assign N14 = \piso.shift_ctr_r [1] & N13;
  assign N15 = \piso.shift_ctr_r [0] & N14;
  assign ready_and_o = fifo0_ready_lo & \piso.fifo1_ready_lo ;
  assign fifo_v_li = valid_i & ready_and_o;
  assign fifo0_yumi_li = N15 & yumi_i;
  assign \piso.fifo1_yumi_li  = N10 & yumi_i;
  assign _0_net_ = N16 & yumi_i;
  assign N16 = ~fifo0_yumi_li;

endmodule

