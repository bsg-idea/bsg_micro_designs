

module top
(
  en_ls_i,
  clk_i,
  reset_i,
  clk_o,
  reset_o,
  fsb_v_i_o,
  fsb_data_i_o,
  fsb_yumi_o_i,
  fsb_v_o_i,
  fsb_data_o_i,
  fsb_ready_i_o,
  node_v_i_o,
  node_data_i_o,
  node_ready_o_i,
  node_v_o_i,
  node_data_o_i,
  node_yumi_i_o
);

  output [49:0] fsb_data_i_o;
  input [49:0] fsb_data_o_i;
  output [49:0] node_data_i_o;
  input [49:0] node_data_o_i;
  input en_ls_i;
  input clk_i;
  input reset_i;
  input fsb_yumi_o_i;
  input fsb_v_o_i;
  input node_ready_o_i;
  input node_v_o_i;
  output clk_o;
  output reset_o;
  output fsb_v_i_o;
  output fsb_ready_i_o;
  output node_v_i_o;
  output node_yumi_i_o;

  bsg_fsb_node_level_shift_node_domain
  wrapper
  (
    .fsb_data_i_o(fsb_data_i_o),
    .fsb_data_o_i(fsb_data_o_i),
    .node_data_i_o(node_data_i_o),
    .node_data_o_i(node_data_o_i),
    .en_ls_i(en_ls_i),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .fsb_yumi_o_i(fsb_yumi_o_i),
    .fsb_v_o_i(fsb_v_o_i),
    .node_ready_o_i(node_ready_o_i),
    .node_v_o_i(node_v_o_i),
    .clk_o(clk_o),
    .reset_o(reset_o),
    .fsb_v_i_o(fsb_v_i_o),
    .fsb_ready_i_o(fsb_ready_i_o),
    .node_v_i_o(node_v_i_o),
    .node_yumi_i_o(node_yumi_i_o)
  );


endmodule



module bsg_level_shift_up_down_sink_width_p1
(
  v0_data_i,
  v1_en_i,
  v1_data_o
);

  input [0:0] v0_data_i;
  output [0:0] v1_data_o;
  input v1_en_i;
  wire [0:0] v1_data_o;
  assign v1_data_o[0] = v0_data_i[0] & v1_en_i;

endmodule



module bsg_level_shift_up_down_source_width_p1
(
  v0_en_i,
  v0_data_i,
  v1_data_o
);

  input [0:0] v0_data_i;
  output [0:0] v1_data_o;
  input v0_en_i;
  wire [0:0] v1_data_o;
  assign v1_data_o[0] = v0_data_i[0] & v0_en_i;

endmodule



module bsg_level_shift_up_down_source_width_p50
(
  v0_en_i,
  v0_data_i,
  v1_data_o
);

  input [49:0] v0_data_i;
  output [49:0] v1_data_o;
  input v0_en_i;
  wire [49:0] v1_data_o;
  assign v1_data_o[49] = v0_data_i[49] & v0_en_i;
  assign v1_data_o[48] = v0_data_i[48] & v0_en_i;
  assign v1_data_o[47] = v0_data_i[47] & v0_en_i;
  assign v1_data_o[46] = v0_data_i[46] & v0_en_i;
  assign v1_data_o[45] = v0_data_i[45] & v0_en_i;
  assign v1_data_o[44] = v0_data_i[44] & v0_en_i;
  assign v1_data_o[43] = v0_data_i[43] & v0_en_i;
  assign v1_data_o[42] = v0_data_i[42] & v0_en_i;
  assign v1_data_o[41] = v0_data_i[41] & v0_en_i;
  assign v1_data_o[40] = v0_data_i[40] & v0_en_i;
  assign v1_data_o[39] = v0_data_i[39] & v0_en_i;
  assign v1_data_o[38] = v0_data_i[38] & v0_en_i;
  assign v1_data_o[37] = v0_data_i[37] & v0_en_i;
  assign v1_data_o[36] = v0_data_i[36] & v0_en_i;
  assign v1_data_o[35] = v0_data_i[35] & v0_en_i;
  assign v1_data_o[34] = v0_data_i[34] & v0_en_i;
  assign v1_data_o[33] = v0_data_i[33] & v0_en_i;
  assign v1_data_o[32] = v0_data_i[32] & v0_en_i;
  assign v1_data_o[31] = v0_data_i[31] & v0_en_i;
  assign v1_data_o[30] = v0_data_i[30] & v0_en_i;
  assign v1_data_o[29] = v0_data_i[29] & v0_en_i;
  assign v1_data_o[28] = v0_data_i[28] & v0_en_i;
  assign v1_data_o[27] = v0_data_i[27] & v0_en_i;
  assign v1_data_o[26] = v0_data_i[26] & v0_en_i;
  assign v1_data_o[25] = v0_data_i[25] & v0_en_i;
  assign v1_data_o[24] = v0_data_i[24] & v0_en_i;
  assign v1_data_o[23] = v0_data_i[23] & v0_en_i;
  assign v1_data_o[22] = v0_data_i[22] & v0_en_i;
  assign v1_data_o[21] = v0_data_i[21] & v0_en_i;
  assign v1_data_o[20] = v0_data_i[20] & v0_en_i;
  assign v1_data_o[19] = v0_data_i[19] & v0_en_i;
  assign v1_data_o[18] = v0_data_i[18] & v0_en_i;
  assign v1_data_o[17] = v0_data_i[17] & v0_en_i;
  assign v1_data_o[16] = v0_data_i[16] & v0_en_i;
  assign v1_data_o[15] = v0_data_i[15] & v0_en_i;
  assign v1_data_o[14] = v0_data_i[14] & v0_en_i;
  assign v1_data_o[13] = v0_data_i[13] & v0_en_i;
  assign v1_data_o[12] = v0_data_i[12] & v0_en_i;
  assign v1_data_o[11] = v0_data_i[11] & v0_en_i;
  assign v1_data_o[10] = v0_data_i[10] & v0_en_i;
  assign v1_data_o[9] = v0_data_i[9] & v0_en_i;
  assign v1_data_o[8] = v0_data_i[8] & v0_en_i;
  assign v1_data_o[7] = v0_data_i[7] & v0_en_i;
  assign v1_data_o[6] = v0_data_i[6] & v0_en_i;
  assign v1_data_o[5] = v0_data_i[5] & v0_en_i;
  assign v1_data_o[4] = v0_data_i[4] & v0_en_i;
  assign v1_data_o[3] = v0_data_i[3] & v0_en_i;
  assign v1_data_o[2] = v0_data_i[2] & v0_en_i;
  assign v1_data_o[1] = v0_data_i[1] & v0_en_i;
  assign v1_data_o[0] = v0_data_i[0] & v0_en_i;

endmodule



module bsg_level_shift_up_down_sink_width_p50
(
  v0_data_i,
  v1_en_i,
  v1_data_o
);

  input [49:0] v0_data_i;
  output [49:0] v1_data_o;
  input v1_en_i;
  wire [49:0] v1_data_o;
  assign v1_data_o[49] = v0_data_i[49] & v1_en_i;
  assign v1_data_o[48] = v0_data_i[48] & v1_en_i;
  assign v1_data_o[47] = v0_data_i[47] & v1_en_i;
  assign v1_data_o[46] = v0_data_i[46] & v1_en_i;
  assign v1_data_o[45] = v0_data_i[45] & v1_en_i;
  assign v1_data_o[44] = v0_data_i[44] & v1_en_i;
  assign v1_data_o[43] = v0_data_i[43] & v1_en_i;
  assign v1_data_o[42] = v0_data_i[42] & v1_en_i;
  assign v1_data_o[41] = v0_data_i[41] & v1_en_i;
  assign v1_data_o[40] = v0_data_i[40] & v1_en_i;
  assign v1_data_o[39] = v0_data_i[39] & v1_en_i;
  assign v1_data_o[38] = v0_data_i[38] & v1_en_i;
  assign v1_data_o[37] = v0_data_i[37] & v1_en_i;
  assign v1_data_o[36] = v0_data_i[36] & v1_en_i;
  assign v1_data_o[35] = v0_data_i[35] & v1_en_i;
  assign v1_data_o[34] = v0_data_i[34] & v1_en_i;
  assign v1_data_o[33] = v0_data_i[33] & v1_en_i;
  assign v1_data_o[32] = v0_data_i[32] & v1_en_i;
  assign v1_data_o[31] = v0_data_i[31] & v1_en_i;
  assign v1_data_o[30] = v0_data_i[30] & v1_en_i;
  assign v1_data_o[29] = v0_data_i[29] & v1_en_i;
  assign v1_data_o[28] = v0_data_i[28] & v1_en_i;
  assign v1_data_o[27] = v0_data_i[27] & v1_en_i;
  assign v1_data_o[26] = v0_data_i[26] & v1_en_i;
  assign v1_data_o[25] = v0_data_i[25] & v1_en_i;
  assign v1_data_o[24] = v0_data_i[24] & v1_en_i;
  assign v1_data_o[23] = v0_data_i[23] & v1_en_i;
  assign v1_data_o[22] = v0_data_i[22] & v1_en_i;
  assign v1_data_o[21] = v0_data_i[21] & v1_en_i;
  assign v1_data_o[20] = v0_data_i[20] & v1_en_i;
  assign v1_data_o[19] = v0_data_i[19] & v1_en_i;
  assign v1_data_o[18] = v0_data_i[18] & v1_en_i;
  assign v1_data_o[17] = v0_data_i[17] & v1_en_i;
  assign v1_data_o[16] = v0_data_i[16] & v1_en_i;
  assign v1_data_o[15] = v0_data_i[15] & v1_en_i;
  assign v1_data_o[14] = v0_data_i[14] & v1_en_i;
  assign v1_data_o[13] = v0_data_i[13] & v1_en_i;
  assign v1_data_o[12] = v0_data_i[12] & v1_en_i;
  assign v1_data_o[11] = v0_data_i[11] & v1_en_i;
  assign v1_data_o[10] = v0_data_i[10] & v1_en_i;
  assign v1_data_o[9] = v0_data_i[9] & v1_en_i;
  assign v1_data_o[8] = v0_data_i[8] & v1_en_i;
  assign v1_data_o[7] = v0_data_i[7] & v1_en_i;
  assign v1_data_o[6] = v0_data_i[6] & v1_en_i;
  assign v1_data_o[5] = v0_data_i[5] & v1_en_i;
  assign v1_data_o[4] = v0_data_i[4] & v1_en_i;
  assign v1_data_o[3] = v0_data_i[3] & v1_en_i;
  assign v1_data_o[2] = v0_data_i[2] & v1_en_i;
  assign v1_data_o[1] = v0_data_i[1] & v1_en_i;
  assign v1_data_o[0] = v0_data_i[0] & v1_en_i;

endmodule



module bsg_fsb_node_level_shift_node_domain
(
  en_ls_i,
  clk_i,
  reset_i,
  clk_o,
  reset_o,
  fsb_v_i_o,
  fsb_data_i_o,
  fsb_yumi_o_i,
  fsb_v_o_i,
  fsb_data_o_i,
  fsb_ready_i_o,
  node_v_i_o,
  node_data_i_o,
  node_ready_o_i,
  node_v_o_i,
  node_data_o_i,
  node_yumi_i_o
);

  output [49:0] fsb_data_i_o;
  input [49:0] fsb_data_o_i;
  output [49:0] node_data_i_o;
  input [49:0] node_data_o_i;
  input en_ls_i;
  input clk_i;
  input reset_i;
  input fsb_yumi_o_i;
  input fsb_v_o_i;
  input node_ready_o_i;
  input node_v_o_i;
  output clk_o;
  output reset_o;
  output fsb_v_i_o;
  output fsb_ready_i_o;
  output node_v_i_o;
  output node_yumi_i_o;
  wire [49:0] fsb_data_i_o,node_data_i_o;
  wire clk_o,reset_o,fsb_v_i_o,fsb_ready_i_o,node_v_i_o,node_yumi_i_o;

  bsg_level_shift_up_down_sink_width_p1
  clk_ls_inst
  (
    .v0_data_i(clk_i),
    .v1_en_i(1'b1),
    .v1_data_o(clk_o)
  );


  bsg_level_shift_up_down_sink_width_p1
  reset_ls_inst
  (
    .v0_data_i(reset_i),
    .v1_en_i(1'b1),
    .v1_data_o(reset_o)
  );


  bsg_level_shift_up_down_source_width_p1
  n2f_v_ls_inst
  (
    .v0_en_i(en_ls_i),
    .v0_data_i(node_v_o_i),
    .v1_data_o(fsb_v_i_o)
  );


  bsg_level_shift_up_down_source_width_p50
  n2f_data_ls_inst
  (
    .v0_en_i(en_ls_i),
    .v0_data_i(node_data_o_i),
    .v1_data_o(fsb_data_i_o)
  );


  bsg_level_shift_up_down_sink_width_p1
  f2n_yumi_ls_inst
  (
    .v0_data_i(fsb_yumi_o_i),
    .v1_en_i(en_ls_i),
    .v1_data_o(node_yumi_i_o)
  );


  bsg_level_shift_up_down_sink_width_p1
  f2n_v_ls_inst
  (
    .v0_data_i(fsb_v_o_i),
    .v1_en_i(en_ls_i),
    .v1_data_o(node_v_i_o)
  );


  bsg_level_shift_up_down_sink_width_p50
  f2n_data_ls_inst
  (
    .v0_data_i(fsb_data_o_i),
    .v1_en_i(en_ls_i),
    .v1_data_o(node_data_i_o)
  );


  bsg_level_shift_up_down_source_width_p1
  n2f_ready_ls_inst
  (
    .v0_en_i(en_ls_i),
    .v0_data_i(node_ready_o_i),
    .v1_data_o(fsb_ready_i_o)
  );


endmodule

